magic
tech sky130A
timestamp 1483428465
<< checkpaint >>
rect -785 -785 785 785
<< metal4 >>
rect -155 139 155 155
rect -155 -139 -139 139
rect 139 -139 155 139
rect -155 -155 155 -139
<< via4 >>
rect -139 -139 139 139
<< metal5 >>
rect -155 139 155 155
rect -155 -139 -139 139
rect 139 -139 155 139
rect -155 -155 155 -139
<< end >>
