magic
tech sky130A
timestamp 1483428465
<< checkpaint >>
rect -739 -654 739 654
<< metal3 >>
rect -109 16 109 24
rect -109 -16 -96 16
rect -64 -16 -56 16
rect -24 -16 -16 16
rect 16 -16 24 16
rect 56 -16 64 16
rect 96 -16 109 16
rect -109 -24 109 -16
<< via3 >>
rect -96 -16 -64 16
rect -56 -16 -24 16
rect -16 -16 16 16
rect 24 -16 56 16
rect 64 -16 96 16
<< metal4 >>
rect -109 16 109 24
rect -109 -16 -96 16
rect -64 -16 -56 16
rect -24 -16 -16 16
rect 16 -16 24 16
rect 56 -16 64 16
rect 96 -16 109 16
rect -109 -24 109 -16
<< end >>
