magic
tech sky130A
timestamp 1483428465
<< checkpaint >>
rect -1130 -1085 1130 1085
<< metal4 >>
rect -500 379 500 455
rect -500 -379 -459 379
rect 459 -379 500 379
rect -500 -455 500 -379
<< via4 >>
rect -459 -379 459 379
<< metal5 >>
rect -500 379 500 455
rect -500 -379 -459 379
rect 459 -379 500 379
rect -500 -455 500 -379
<< end >>
