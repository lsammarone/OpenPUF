magic
tech sky130A
magscale 1 2
timestamp 1654736712
<< metal4 >>
rect -1000 278 1000 443
rect -1000 -278 -918 278
rect 918 -278 1000 278
rect -1000 -443 1000 -278
<< via4 >>
rect -918 -278 918 278
<< metal5 >>
rect -1000 278 1000 443
rect -1000 -278 -918 278
rect 918 -278 1000 278
rect -1000 -443 1000 -278
<< end >>
