magic
tech sky130A
magscale 1 2
timestamp 1654736712
<< metal4 >>
rect -1000 278 1000 443
rect -1000 42 -918 278
rect -682 42 -598 278
rect -362 42 -278 278
rect -42 42 42 278
rect -1000 -42 42 42
rect -1000 -278 -918 -42
rect -682 -278 42 -42
rect 918 -278 1000 278
rect -1000 -443 1000 -278
<< via4 >>
rect -918 42 -682 278
rect -598 42 -362 278
rect -278 42 -42 278
rect -918 -278 -682 -42
rect 42 -278 918 278
<< metal5 >>
rect -1000 278 1000 443
rect -1000 42 -918 278
rect -682 42 -598 278
rect -362 42 -278 278
rect -42 42 42 278
rect -1000 -42 42 42
rect -1000 -278 -918 -42
rect -682 -278 42 -42
rect 918 -278 1000 278
rect -1000 -443 1000 -278
<< end >>
