magic
tech sky130A
timestamp 1654736712
<< metal1 >>
rect -86 13 86 24
rect -86 -13 -77 13
rect -51 -13 -45 13
rect -19 -13 -13 13
rect 13 -13 19 13
rect 45 -13 51 13
rect 77 -13 86 13
rect -86 -24 86 -13
<< via1 >>
rect -77 -13 -51 13
rect -45 -13 -19 13
rect -13 -13 13 13
rect 19 -13 45 13
rect 51 -13 77 13
<< metal2 >>
rect -86 13 86 24
rect -86 -13 -77 13
rect -51 -13 -45 13
rect -19 -13 -13 13
rect 13 -13 19 13
rect 45 -13 51 13
rect 77 -13 86 13
rect -86 -24 86 -13
<< end >>
