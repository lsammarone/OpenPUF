magic
tech sky130A
magscale 1 2
timestamp 1656715967
<< nwell >>
rect 2282 4746 3458 4824
rect 4170 4746 5346 4824
rect 17380 4746 18556 4824
rect 19268 4746 20444 4824
<< locali >>
rect 4626 5009 4668 5012
rect 2742 5005 2784 5008
rect 2742 4971 2746 5005
rect 2780 4971 2784 5005
rect 2742 4968 2784 4971
rect 4626 4975 4630 5009
rect 4664 4975 4668 5009
rect 19724 5009 19766 5012
rect 4626 4972 4668 4975
rect 17840 5005 17882 5008
rect 17840 4971 17844 5005
rect 17878 4971 17882 5005
rect 17840 4968 17882 4971
rect 19724 4975 19728 5009
rect 19762 4975 19766 5009
rect 19724 4972 19766 4975
<< viali >>
rect 2368 5146 2402 5180
rect 2560 5146 2594 5180
rect 2752 5146 2786 5180
rect 2944 5146 2978 5180
rect 3136 5146 3170 5180
rect 4142 5140 4176 5174
rect 4292 5140 4326 5174
rect 4442 5140 4476 5174
rect 4592 5140 4626 5174
rect 4742 5140 4776 5174
rect 17585 5143 17619 5177
rect 17713 5143 17747 5177
rect 17841 5143 17875 5177
rect 17969 5143 18003 5177
rect 18097 5143 18131 5177
rect 19320 5140 19354 5174
rect 19448 5140 19482 5174
rect 19576 5140 19610 5174
rect 19704 5140 19738 5174
rect 19832 5140 19866 5174
rect 2245 4973 2279 5007
rect 2411 4971 2445 5005
rect 2575 4969 2609 5003
rect 2746 4971 2780 5005
rect 2915 4967 2949 5001
rect 3084 4966 3118 5000
rect 3250 4972 3284 5006
rect 3420 4974 3454 5008
rect 4134 4971 4168 5005
rect 4294 4971 4328 5005
rect 4461 4965 4495 4999
rect 4630 4975 4664 5009
rect 4794 4962 4828 4996
rect 4964 4968 4998 5002
rect 5134 4970 5168 5004
rect 5293 4972 5327 5006
rect 17343 4967 17377 5001
rect 17506 4962 17540 4996
rect 17679 4966 17713 5000
rect 17844 4971 17878 5005
rect 18011 4958 18045 4992
rect 18179 4956 18213 4990
rect 18349 4965 18383 4999
rect 19222 4966 19256 5000
rect 19395 4967 19429 5001
rect 19557 4972 19591 5006
rect 19728 4975 19762 5009
rect 19897 4961 19931 4995
rect 20062 4961 20096 4995
rect 20232 4959 20266 4993
rect 20395 4963 20429 4997
<< metal1 >>
rect 3656 5194 3912 5246
rect 2304 5180 4916 5194
rect 18772 5192 18996 5254
rect 2304 5146 2368 5180
rect 2402 5146 2560 5180
rect 2594 5146 2752 5180
rect 2786 5146 2944 5180
rect 2978 5146 3136 5180
rect 3170 5174 4916 5180
rect 3170 5146 4142 5174
rect 2304 5140 4142 5146
rect 4176 5140 4292 5174
rect 4326 5140 4442 5174
rect 4476 5140 4592 5174
rect 4626 5140 4742 5174
rect 4776 5140 4916 5174
rect 2304 5128 4916 5140
rect 17570 5177 19902 5192
rect 17570 5143 17585 5177
rect 17619 5143 17713 5177
rect 17747 5143 17841 5177
rect 17875 5143 17969 5177
rect 18003 5143 18097 5177
rect 18131 5174 19902 5177
rect 18131 5143 19320 5174
rect 17570 5140 19320 5143
rect 19354 5140 19448 5174
rect 19482 5140 19576 5174
rect 19610 5140 19704 5174
rect 19738 5140 19832 5174
rect 19866 5140 19902 5174
rect 17570 5124 19902 5140
rect 2230 5008 3467 5020
rect 2230 5007 3420 5008
rect 2230 4973 2245 5007
rect 2279 5006 3420 5007
rect 2279 5005 3250 5006
rect 2279 5002 2411 5005
rect 2445 5004 2746 5005
rect 2780 5004 3250 5005
rect 2445 5003 2740 5004
rect 2445 5002 2575 5003
rect 2279 4973 2282 5002
rect 2230 4950 2282 4973
rect 2334 4950 2389 5002
rect 2445 4971 2495 5002
rect 2441 4950 2495 4971
rect 2547 4969 2575 5002
rect 2609 5002 2740 5003
rect 2609 4969 2611 5002
rect 2547 4950 2611 4969
rect 2663 4952 2740 5002
rect 2792 5003 3250 5004
rect 3284 5003 3420 5006
rect 2792 4952 2874 5003
rect 2926 5001 2991 5003
rect 2949 4967 2991 5001
rect 2663 4951 2874 4952
rect 2926 4951 2991 4967
rect 3043 5000 3096 5003
rect 3043 4966 3084 5000
rect 3043 4951 3096 4966
rect 3148 4951 3202 5003
rect 3284 4972 3299 5003
rect 3254 4951 3299 4972
rect 3351 4951 3396 5003
rect 3454 4974 3467 5008
rect 3448 4951 3467 4974
rect 2663 4950 3467 4951
rect 2230 4936 3467 4950
rect 4120 5009 5346 5018
rect 4120 5005 4630 5009
rect 4120 4971 4134 5005
rect 4168 4999 4294 5005
rect 4328 4999 4630 5005
rect 4168 4971 4171 4999
rect 4120 4947 4171 4971
rect 4223 4947 4278 4999
rect 4330 4947 4384 4999
rect 4436 4965 4461 4999
rect 4495 4965 4500 4999
rect 4436 4947 4500 4965
rect 4552 4975 4630 4999
rect 4664 5006 5346 5009
rect 4664 5004 5293 5006
rect 4664 5002 5134 5004
rect 4664 5000 4964 5002
rect 4998 5000 5134 5002
rect 5168 5000 5293 5004
rect 5327 5000 5346 5006
rect 4664 4975 4763 5000
rect 4815 4996 4880 5000
rect 4552 4948 4763 4975
rect 4828 4962 4880 4996
rect 4815 4948 4880 4962
rect 4932 4968 4964 5000
rect 4932 4948 4985 4968
rect 5037 4948 5091 5000
rect 5168 4970 5188 5000
rect 5143 4948 5188 4970
rect 5240 4948 5285 5000
rect 5337 4948 5346 5000
rect 4552 4947 5346 4948
rect 4120 4934 5346 4947
rect 17321 5008 18588 5020
rect 17321 5001 17391 5008
rect 17321 4967 17343 5001
rect 17377 4967 17391 5001
rect 17321 4956 17391 4967
rect 17443 5006 18588 5008
rect 17443 4956 17503 5006
rect 17321 4954 17503 4956
rect 17555 4954 17610 5006
rect 17662 5000 17712 5006
rect 17764 5005 18588 5006
rect 17764 5004 17844 5005
rect 17878 5004 18588 5005
rect 17662 4966 17679 5000
rect 17662 4954 17712 4966
rect 17764 4954 17838 5004
rect 17321 4952 17838 4954
rect 17890 4952 17992 5004
rect 18044 4992 18129 5004
rect 18045 4958 18129 4992
rect 18181 4990 18226 5004
rect 18044 4952 18129 4958
rect 18213 4956 18226 4990
rect 18181 4952 18226 4956
rect 18278 4952 18326 5004
rect 18378 5003 18588 5004
rect 18378 4999 18415 5003
rect 18383 4965 18415 4999
rect 18378 4952 18415 4965
rect 17321 4951 18415 4952
rect 18467 4951 18511 5003
rect 18563 4951 18588 5003
rect 17321 4936 18588 4951
rect 19207 5009 20463 5018
rect 19207 5006 19728 5009
rect 19207 5002 19557 5006
rect 19591 5002 19728 5006
rect 19762 5002 20463 5009
rect 19207 5000 19225 5002
rect 19207 4966 19222 5000
rect 19207 4950 19225 4966
rect 19277 4950 19319 5002
rect 19371 5001 19418 5002
rect 19371 4967 19395 5001
rect 19371 4950 19418 4967
rect 19470 4950 19526 5002
rect 19591 4972 19622 5002
rect 19578 4950 19622 4972
rect 19674 4950 19720 5002
rect 19772 5001 20463 5002
rect 19772 4950 19839 5001
rect 19207 4949 19839 4950
rect 19891 4995 19953 5001
rect 19891 4961 19897 4995
rect 19931 4961 19953 4995
rect 19891 4949 19953 4961
rect 20005 4995 20070 5001
rect 20005 4961 20062 4995
rect 20005 4949 20070 4961
rect 20122 4949 20197 5001
rect 20249 4993 20312 5001
rect 20266 4959 20312 4993
rect 20249 4949 20312 4959
rect 20364 4997 20463 5001
rect 20364 4963 20395 4997
rect 20429 4963 20463 4997
rect 20364 4949 20463 4963
rect 19207 4934 20463 4949
<< via1 >>
rect 2282 4950 2334 5002
rect 2389 4971 2411 5002
rect 2411 4971 2441 5002
rect 2389 4950 2441 4971
rect 2495 4950 2547 5002
rect 2611 4950 2663 5002
rect 2740 4971 2746 5004
rect 2746 4971 2780 5004
rect 2780 4971 2792 5004
rect 2740 4952 2792 4971
rect 2874 5001 2926 5003
rect 2874 4967 2915 5001
rect 2915 4967 2926 5001
rect 2874 4951 2926 4967
rect 2991 4951 3043 5003
rect 3096 5000 3148 5003
rect 3096 4966 3118 5000
rect 3118 4966 3148 5000
rect 3096 4951 3148 4966
rect 3202 4972 3250 5003
rect 3250 4972 3254 5003
rect 3202 4951 3254 4972
rect 3299 4951 3351 5003
rect 3396 4974 3420 5003
rect 3420 4974 3448 5003
rect 3396 4951 3448 4974
rect 4171 4947 4223 4999
rect 4278 4971 4294 4999
rect 4294 4971 4328 4999
rect 4328 4971 4330 4999
rect 4278 4947 4330 4971
rect 4384 4947 4436 4999
rect 4500 4947 4552 4999
rect 4763 4996 4815 5000
rect 4763 4962 4794 4996
rect 4794 4962 4815 4996
rect 4763 4948 4815 4962
rect 4880 4948 4932 5000
rect 4985 4968 4998 5000
rect 4998 4968 5037 5000
rect 4985 4948 5037 4968
rect 5091 4970 5134 5000
rect 5134 4970 5143 5000
rect 5091 4948 5143 4970
rect 5188 4948 5240 5000
rect 5285 4972 5293 5000
rect 5293 4972 5327 5000
rect 5327 4972 5337 5000
rect 5285 4948 5337 4972
rect 17391 4956 17443 5008
rect 17503 4996 17555 5006
rect 17503 4962 17506 4996
rect 17506 4962 17540 4996
rect 17540 4962 17555 4996
rect 17503 4954 17555 4962
rect 17610 4954 17662 5006
rect 17712 5000 17764 5006
rect 17712 4966 17713 5000
rect 17713 4966 17764 5000
rect 17712 4954 17764 4966
rect 17838 4971 17844 5004
rect 17844 4971 17878 5004
rect 17878 4971 17890 5004
rect 17838 4952 17890 4971
rect 17992 4992 18044 5004
rect 17992 4958 18011 4992
rect 18011 4958 18044 4992
rect 18129 4990 18181 5004
rect 17992 4952 18044 4958
rect 18129 4956 18179 4990
rect 18179 4956 18181 4990
rect 18129 4952 18181 4956
rect 18226 4952 18278 5004
rect 18326 4999 18378 5004
rect 18326 4965 18349 4999
rect 18349 4965 18378 4999
rect 18326 4952 18378 4965
rect 18415 4951 18467 5003
rect 18511 4951 18563 5003
rect 19225 5000 19277 5002
rect 19225 4966 19256 5000
rect 19256 4966 19277 5000
rect 19225 4950 19277 4966
rect 19319 4950 19371 5002
rect 19418 5001 19470 5002
rect 19418 4967 19429 5001
rect 19429 4967 19470 5001
rect 19418 4950 19470 4967
rect 19526 4972 19557 5002
rect 19557 4972 19578 5002
rect 19526 4950 19578 4972
rect 19622 4950 19674 5002
rect 19720 4975 19728 5002
rect 19728 4975 19762 5002
rect 19762 4975 19772 5002
rect 19720 4950 19772 4975
rect 19839 4949 19891 5001
rect 19953 4949 20005 5001
rect 20070 4995 20122 5001
rect 20070 4961 20096 4995
rect 20096 4961 20122 4995
rect 20070 4949 20122 4961
rect 20197 4993 20249 5001
rect 20197 4959 20232 4993
rect 20232 4959 20249 4993
rect 20197 4949 20249 4959
rect 20312 4949 20364 5001
<< metal2 >>
rect -1439 5082 -413 5083
rect 446 5082 1472 5084
rect 13643 5082 14669 5084
rect 15544 5082 16570 5083
rect 21211 5082 22237 5086
rect 23115 5082 24141 5083
rect -3546 5020 11208 5082
rect 11562 5020 26308 5082
rect -3544 5004 11208 5020
rect -3544 5002 2740 5004
rect -3544 4950 2282 5002
rect 2334 4950 2389 5002
rect 2441 4950 2495 5002
rect 2547 4950 2611 5002
rect 2663 4952 2740 5002
rect 2792 5003 11208 5004
rect 2792 4952 2874 5003
rect 2663 4951 2874 4952
rect 2926 4951 2991 5003
rect 3043 4951 3096 5003
rect 3148 4951 3202 5003
rect 3254 4951 3299 5003
rect 3351 4951 3396 5003
rect 3448 5000 11208 5003
rect 3448 4999 4763 5000
rect 3448 4951 4171 4999
rect 2663 4950 4171 4951
rect -3544 4947 4171 4950
rect 4223 4947 4278 4999
rect 4330 4947 4384 4999
rect 4436 4947 4500 4999
rect 4552 4948 4763 4999
rect 4815 4948 4880 5000
rect 4932 4948 4985 5000
rect 5037 4948 5091 5000
rect 5143 4948 5188 5000
rect 5240 4948 5285 5000
rect 5337 4948 11208 5000
rect 11563 5008 26308 5020
rect 11563 4956 17391 5008
rect 17443 5006 26308 5008
rect 17443 4956 17503 5006
rect 4552 4947 11208 4948
rect -3544 4894 11208 4947
rect 11562 4954 17503 4956
rect 17555 4954 17610 5006
rect 17662 4954 17712 5006
rect 17764 5004 26308 5006
rect 17764 4954 17838 5004
rect 11562 4952 17838 4954
rect 17890 4952 17992 5004
rect 18044 4952 18129 5004
rect 18181 4952 18226 5004
rect 18278 4952 18326 5004
rect 18378 5003 26308 5004
rect 18378 4952 18415 5003
rect 11562 4951 18415 4952
rect 18467 4951 18511 5003
rect 18563 5002 26308 5003
rect 18563 4951 19225 5002
rect 11562 4950 19225 4951
rect 19277 4950 19319 5002
rect 19371 4950 19418 5002
rect 19470 4950 19526 5002
rect 19578 4950 19622 5002
rect 19674 4950 19720 5002
rect 19772 5001 26308 5002
rect 19772 4950 19839 5001
rect 11562 4949 19839 4950
rect 19891 4949 19953 5001
rect 20005 4949 20070 5001
rect 20122 4949 20197 5001
rect 20249 4949 20312 5001
rect 20364 4949 26308 5001
rect 11562 4894 26308 4949
rect -3326 4637 -2300 4894
rect -1439 4637 -413 4894
rect 446 4637 1472 4894
rect 2150 4886 5358 4894
rect 2150 4637 3470 4886
rect -3544 4590 3470 4637
rect 4034 4633 5358 4886
rect 6115 4633 7141 4894
rect 8010 4633 9036 4894
rect 9879 4633 10905 4894
rect 11756 4637 12782 4894
rect 13643 4637 14669 4894
rect 15544 4637 16570 4894
rect 17248 4886 20456 4894
rect 17248 4637 18568 4886
rect 19132 4637 20456 4886
rect 21211 4637 22237 4894
rect 23115 4637 24141 4894
rect 24991 4637 26017 4894
rect 4034 4590 11208 4633
rect -3544 4528 11208 4590
rect 11562 4590 26307 4637
rect 11562 4528 26306 4590
rect 2150 4524 3470 4528
rect 4034 4524 11208 4528
rect 17248 4524 18568 4528
rect 19132 4524 20456 4528
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0
timestamp 1656715967
transform 1 0 19092 0 -1 5396
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1656715967
transform 1 0 17210 0 -1 5398
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_2
timestamp 1656715967
transform 1 0 3994 0 -1 5396
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_3
timestamp 1656715967
transform 1 0 2112 0 -1 5398
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_4
timestamp 1656715967
transform 1 0 19092 0 -1 5396
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_5
timestamp 1656715967
transform 1 0 17210 0 -1 5398
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_6
timestamp 1656715967
transform 1 0 3994 0 -1 5396
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_7
timestamp 1656715967
transform 1 0 2112 0 -1 5398
box -38 -48 1510 592
use unitcell2buf  unitcell2buf_0
timestamp 1656715967
transform 1 0 23448 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_1
timestamp 1656715967
transform 1 0 21560 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_2
timestamp 1656715967
transform 1 0 19672 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_3
timestamp 1656715967
transform 1 0 17784 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_4
timestamp 1656715967
transform 1 0 15896 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_5
timestamp 1656715967
transform 1 0 14008 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_6
timestamp 1656715967
transform 1 0 12120 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_7
timestamp 1656715967
transform 1 0 8350 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_8
timestamp 1656715967
transform 1 0 6462 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_9
timestamp 1656715967
transform 1 0 4574 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_10
timestamp 1656715967
transform 1 0 2686 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_11
timestamp 1656715967
transform 1 0 798 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_12
timestamp 1656715967
transform 1 0 -2978 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_13
timestamp 1656715967
transform 1 0 -1090 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_14
timestamp 1656715967
transform 1 0 23448 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_15
timestamp 1656715967
transform 1 0 21560 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_16
timestamp 1656715967
transform 1 0 19672 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_17
timestamp 1656715967
transform 1 0 17784 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_18
timestamp 1656715967
transform 1 0 15896 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_19
timestamp 1656715967
transform 1 0 14008 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_20
timestamp 1656715967
transform 1 0 12120 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_21
timestamp 1656715967
transform 1 0 8350 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_22
timestamp 1656715967
transform 1 0 6462 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_23
timestamp 1656715967
transform 1 0 4574 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_24
timestamp 1656715967
transform 1 0 2686 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_25
timestamp 1656715967
transform 1 0 798 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_26
timestamp 1656715967
transform 1 0 -2978 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_27
timestamp 1656715967
transform 1 0 -1090 0 1 3712
box -574 -1185 1322 1192
use unitcell2bufcut  unitcell2bufcut_0
timestamp 1656715967
transform 1 0 25336 0 1 3712
box -574 -1184 1322 1192
use unitcell2bufcut  unitcell2bufcut_1
timestamp 1656715967
transform 1 0 10238 0 1 3712
box -574 -1184 1322 1192
use unitcell2bufcut  unitcell2bufcut_2
timestamp 1656715967
transform 1 0 25336 0 1 3712
box -574 -1184 1322 1192
use unitcell2bufcut  unitcell2bufcut_3
timestamp 1656715967
transform 1 0 10238 0 1 3712
box -574 -1184 1322 1192
<< properties >>
string GDS_END 9427070
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/design_merged.gds
string GDS_START 9400314
<< end >>
