magic
tech sky130A
magscale 1 2
timestamp 1656715967
<< metal4 >>
rect -309 918 309 1000
rect -309 -918 -278 918
rect 278 -918 309 918
rect -309 -1000 309 -918
<< via4 >>
rect -278 -918 278 918
<< metal5 >>
rect -309 918 309 1000
rect -309 -918 -278 918
rect 278 -918 309 918
rect -309 -1000 309 -918
<< properties >>
string GDS_END 9321222
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/design_merged.gds
string GDS_START 9320322
<< end >>
