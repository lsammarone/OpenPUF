magic
tech sky130A
timestamp 1656729169
<< error_p >>
rect -71 71 71 89
rect -71 59 89 71
rect -71 -59 -59 59
rect 71 -59 89 59
rect -71 -71 89 -59
<< via4 >>
rect -59 -59 59 59
<< metal5 >>
rect -71 59 71 71
rect -71 -59 -59 59
rect 59 -59 71 59
rect -71 -71 71 -59
<< properties >>
string GDS_END 9297588
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/merge/design_merged.gds
string GDS_START 9297392
<< end >>
