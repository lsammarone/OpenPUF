magic
tech sky130A
timestamp 1483428465
<< checkpaint >>
rect -720 -675 720 675
<< metal3 >>
rect -90 36 90 45
rect -90 -36 -76 36
rect 76 -36 90 36
rect -90 -45 90 -36
<< via3 >>
rect -76 -36 76 36
<< metal4 >>
rect -90 36 90 45
rect -90 -36 -76 36
rect 76 -36 90 36
rect -90 -45 90 -36
<< end >>
