magic
tech sky130A
magscale 1 2
timestamp 1483428465
<< checkpaint >>
rect -1569 -2260 1569 2260
<< metal4 >>
rect -309 918 309 1000
rect -309 -918 -278 918
rect 278 -918 309 918
rect -309 -1000 309 -918
<< via4 >>
rect -278 -918 278 918
<< metal5 >>
rect -309 918 309 1000
rect -309 -918 -278 918
rect 278 -918 309 918
rect -309 -1000 309 -918
<< end >>
