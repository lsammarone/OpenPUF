magic
tech sky130A
magscale 1 2
timestamp 1656715967
<< metal4 >>
rect -392 918 392 963
rect -392 -918 -278 918
rect 278 -918 392 918
rect -392 -963 392 -918
<< via4 >>
rect -278 -918 278 918
<< metal5 >>
rect -392 918 392 963
rect -392 -918 -278 918
rect 278 -918 392 918
rect -392 -963 392 -918
<< properties >>
string GDS_END 9318454
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/design_merged.gds
string GDS_START 9317554
<< end >>
