magic
tech sky130A
magscale 1 2
timestamp 1656715967
<< error_p >>
rect -38 261 314 582
rect 27 47 79 151
rect 109 47 167 151
rect 197 47 249 151
<< nwell >>
rect -38 261 314 582
<< pwell >>
rect 1 21 275 177
rect 31 -17 65 21
<< scnmos >>
rect 79 47 109 151
rect 167 47 197 151
<< scpmoshvt >>
rect 79 339 109 497
rect 167 339 197 497
<< ndiff >>
rect 27 106 79 151
rect 27 72 35 106
rect 69 72 79 106
rect 27 47 79 72
rect 109 93 167 151
rect 109 59 121 93
rect 155 59 167 93
rect 109 47 167 59
rect 197 123 249 151
rect 197 89 207 123
rect 241 89 249 123
rect 197 47 249 89
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 339 79 375
rect 109 477 167 497
rect 109 443 121 477
rect 155 443 167 477
rect 109 409 167 443
rect 109 375 121 409
rect 155 375 167 409
rect 109 339 167 375
rect 197 477 249 497
rect 197 443 207 477
rect 241 443 249 477
rect 197 396 249 443
rect 197 362 207 396
rect 241 362 249 396
rect 197 339 249 362
<< ndiffc >>
rect 35 72 69 106
rect 121 59 155 93
rect 207 89 241 123
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 121 443 155 477
rect 121 375 155 409
rect 207 443 241 477
rect 207 362 241 396
<< poly >>
rect 79 497 109 523
rect 167 497 197 523
rect 79 324 109 339
rect 73 300 109 324
rect 73 265 103 300
rect 167 278 197 339
rect 27 249 103 265
rect 27 215 37 249
rect 71 215 103 249
rect 27 199 103 215
rect 145 262 199 278
rect 145 228 155 262
rect 189 228 199 262
rect 145 212 199 228
rect 73 190 103 199
rect 73 166 109 190
rect 79 151 109 166
rect 167 151 197 212
rect 79 21 109 47
rect 167 21 197 47
<< polycont >>
rect 37 215 71 249
rect 155 228 189 262
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 33 477 69 493
rect 33 443 35 477
rect 33 409 69 443
rect 33 375 35 409
rect 105 477 171 527
rect 105 443 121 477
rect 155 443 171 477
rect 105 409 171 443
rect 105 375 121 409
rect 155 375 171 409
rect 205 477 259 493
rect 205 443 207 477
rect 241 443 259 477
rect 205 396 259 443
rect 33 341 69 375
rect 205 362 207 396
rect 241 362 259 396
rect 33 307 168 341
rect 205 312 259 362
rect 134 278 168 307
rect 21 249 89 271
rect 21 215 37 249
rect 71 215 89 249
rect 21 197 89 215
rect 134 262 189 278
rect 134 228 155 262
rect 134 212 189 228
rect 134 161 168 212
rect 35 127 168 161
rect 223 152 259 312
rect 35 106 69 127
rect 207 123 259 152
rect 35 51 69 72
rect 105 59 121 93
rect 155 59 171 93
rect 105 17 171 59
rect 241 89 259 123
rect 207 51 259 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
<< metal1 >>
rect 0 561 276 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 496 276 527
rect 0 17 276 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 0 -48 276 -17
<< labels >>
flabel metal1 s 31 -17 65 17 0 FreeSans 200 0 0 0 VGND
port 1 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel locali s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel locali s 31 -17 65 17 0 FreeSans 200 0 0 0 VGND
port 1 nsew
flabel locali s 211 85 245 119 0 FreeSans 200 0 0 0 X
port 3 nsew
flabel locali s 211 357 245 391 0 FreeSans 200 0 0 0 X
port 3 nsew
flabel locali s 211 425 245 459 0 FreeSans 200 0 0 0 X
port 3 nsew
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 4 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 31 -17 65 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
rlabel comment s 0 0 0 0 4 buf_1
<< properties >>
string FIXED_BBOX 0 0 276 544
string GDS_END 9891810
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/design_merged.gds
string GDS_START 9866782
string path 0.000 13.600 6.900 13.600 
<< end >>
