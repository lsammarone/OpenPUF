magic
tech sky130A
timestamp 1656729169
<< metal4 >>
rect -155 459 155 500
rect -155 -459 -139 459
rect 139 -459 155 459
rect -155 -500 155 -459
<< via4 >>
rect -139 -459 139 459
<< metal5 >>
rect -155 459 155 500
rect -155 -459 -139 459
rect 139 -459 155 459
rect -155 -500 155 -459
<< properties >>
string GDS_END 9313400
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/merge/design_merged.gds
string GDS_START 9312500
<< end >>
