magic
tech sky130A
magscale 1 2
timestamp 1654904630
<< nwell >>
rect 575170 493276 580556 493654
rect 575169 492152 580556 493276
rect 574448 404400 579834 404778
rect 574447 403276 579834 404400
rect 574644 358972 580030 359350
rect 574643 357848 580030 358972
rect 575092 312804 580478 313182
rect 575091 311680 580478 312804
<< pwell >>
rect 560650 491970 565964 493466
rect 565000 491940 565964 491970
rect 560586 402828 565900 404324
rect 564936 402798 565900 402828
rect 560542 357510 565856 359006
rect 564892 357480 565856 357510
rect 560404 311202 565718 312698
rect 564754 311172 565718 311202
<< pmoslvt >>
rect 575263 492214 575463 493214
rect 575521 492214 575721 493214
rect 575779 492214 575979 493214
rect 576037 492214 576237 493214
rect 576295 492214 576495 493214
rect 576553 492214 576753 493214
rect 576811 492214 577011 493214
rect 577069 492214 577269 493214
rect 577327 492214 577527 493214
rect 577585 492214 577785 493214
rect 577843 492214 578043 493214
rect 578101 492214 578301 493214
rect 578359 492214 578559 493214
rect 578617 492214 578817 493214
rect 578875 492214 579075 493214
rect 579133 492214 579333 493214
rect 579391 492214 579591 493214
rect 579649 492214 579849 493214
rect 579907 492214 580107 493214
rect 580165 492214 580365 493214
rect 574541 403338 574741 404338
rect 574799 403338 574999 404338
rect 575057 403338 575257 404338
rect 575315 403338 575515 404338
rect 575573 403338 575773 404338
rect 575831 403338 576031 404338
rect 576089 403338 576289 404338
rect 576347 403338 576547 404338
rect 576605 403338 576805 404338
rect 576863 403338 577063 404338
rect 577121 403338 577321 404338
rect 577379 403338 577579 404338
rect 577637 403338 577837 404338
rect 577895 403338 578095 404338
rect 578153 403338 578353 404338
rect 578411 403338 578611 404338
rect 578669 403338 578869 404338
rect 578927 403338 579127 404338
rect 579185 403338 579385 404338
rect 579443 403338 579643 404338
rect 574737 357910 574937 358910
rect 574995 357910 575195 358910
rect 575253 357910 575453 358910
rect 575511 357910 575711 358910
rect 575769 357910 575969 358910
rect 576027 357910 576227 358910
rect 576285 357910 576485 358910
rect 576543 357910 576743 358910
rect 576801 357910 577001 358910
rect 577059 357910 577259 358910
rect 577317 357910 577517 358910
rect 577575 357910 577775 358910
rect 577833 357910 578033 358910
rect 578091 357910 578291 358910
rect 578349 357910 578549 358910
rect 578607 357910 578807 358910
rect 578865 357910 579065 358910
rect 579123 357910 579323 358910
rect 579381 357910 579581 358910
rect 579639 357910 579839 358910
rect 575185 311742 575385 312742
rect 575443 311742 575643 312742
rect 575701 311742 575901 312742
rect 575959 311742 576159 312742
rect 576217 311742 576417 312742
rect 576475 311742 576675 312742
rect 576733 311742 576933 312742
rect 576991 311742 577191 312742
rect 577249 311742 577449 312742
rect 577507 311742 577707 312742
rect 577765 311742 577965 312742
rect 578023 311742 578223 312742
rect 578281 311742 578481 312742
rect 578539 311742 578739 312742
rect 578797 311742 578997 312742
rect 579055 311742 579255 312742
rect 579313 311742 579513 312742
rect 579571 311742 579771 312742
rect 579829 311742 580029 312742
rect 580087 311742 580287 312742
<< nmoslvt >>
rect 560707 492440 560907 493440
rect 560965 492440 561165 493440
rect 561223 492440 561423 493440
rect 561481 492440 561681 493440
rect 561739 492440 561939 493440
rect 561997 492440 562197 493440
rect 562255 492440 562455 493440
rect 562513 492440 562713 493440
rect 562771 492440 562971 493440
rect 563029 492440 563229 493440
rect 563287 492440 563487 493440
rect 563545 492440 563745 493440
rect 563803 492440 564003 493440
rect 564061 492440 564261 493440
rect 564319 492440 564519 493440
rect 564577 492440 564777 493440
rect 564835 492440 565035 493440
rect 565093 492440 565293 493440
rect 565351 492440 565551 493440
rect 565609 492440 565809 493440
rect 560643 403298 560843 404298
rect 560901 403298 561101 404298
rect 561159 403298 561359 404298
rect 561417 403298 561617 404298
rect 561675 403298 561875 404298
rect 561933 403298 562133 404298
rect 562191 403298 562391 404298
rect 562449 403298 562649 404298
rect 562707 403298 562907 404298
rect 562965 403298 563165 404298
rect 563223 403298 563423 404298
rect 563481 403298 563681 404298
rect 563739 403298 563939 404298
rect 563997 403298 564197 404298
rect 564255 403298 564455 404298
rect 564513 403298 564713 404298
rect 564771 403298 564971 404298
rect 565029 403298 565229 404298
rect 565287 403298 565487 404298
rect 565545 403298 565745 404298
rect 560599 357980 560799 358980
rect 560857 357980 561057 358980
rect 561115 357980 561315 358980
rect 561373 357980 561573 358980
rect 561631 357980 561831 358980
rect 561889 357980 562089 358980
rect 562147 357980 562347 358980
rect 562405 357980 562605 358980
rect 562663 357980 562863 358980
rect 562921 357980 563121 358980
rect 563179 357980 563379 358980
rect 563437 357980 563637 358980
rect 563695 357980 563895 358980
rect 563953 357980 564153 358980
rect 564211 357980 564411 358980
rect 564469 357980 564669 358980
rect 564727 357980 564927 358980
rect 564985 357980 565185 358980
rect 565243 357980 565443 358980
rect 565501 357980 565701 358980
rect 560461 311672 560661 312672
rect 560719 311672 560919 312672
rect 560977 311672 561177 312672
rect 561235 311672 561435 312672
rect 561493 311672 561693 312672
rect 561751 311672 561951 312672
rect 562009 311672 562209 312672
rect 562267 311672 562467 312672
rect 562525 311672 562725 312672
rect 562783 311672 562983 312672
rect 563041 311672 563241 312672
rect 563299 311672 563499 312672
rect 563557 311672 563757 312672
rect 563815 311672 564015 312672
rect 564073 311672 564273 312672
rect 564331 311672 564531 312672
rect 564589 311672 564789 312672
rect 564847 311672 565047 312672
rect 565105 311672 565305 312672
rect 565363 311672 565563 312672
<< ndiff >>
rect 560649 493428 560707 493440
rect 560649 492452 560661 493428
rect 560695 492452 560707 493428
rect 560649 492440 560707 492452
rect 560907 493428 560965 493440
rect 560907 492452 560919 493428
rect 560953 492452 560965 493428
rect 560907 492440 560965 492452
rect 561165 493428 561223 493440
rect 561165 492452 561177 493428
rect 561211 492452 561223 493428
rect 561165 492440 561223 492452
rect 561423 493428 561481 493440
rect 561423 492452 561435 493428
rect 561469 492452 561481 493428
rect 561423 492440 561481 492452
rect 561681 493428 561739 493440
rect 561681 492452 561693 493428
rect 561727 492452 561739 493428
rect 561681 492440 561739 492452
rect 561939 493428 561997 493440
rect 561939 492452 561951 493428
rect 561985 492452 561997 493428
rect 561939 492440 561997 492452
rect 562197 493428 562255 493440
rect 562197 492452 562209 493428
rect 562243 492452 562255 493428
rect 562197 492440 562255 492452
rect 562455 493428 562513 493440
rect 562455 492452 562467 493428
rect 562501 492452 562513 493428
rect 562455 492440 562513 492452
rect 562713 493428 562771 493440
rect 562713 492452 562725 493428
rect 562759 492452 562771 493428
rect 562713 492440 562771 492452
rect 562971 493428 563029 493440
rect 562971 492452 562983 493428
rect 563017 492452 563029 493428
rect 562971 492440 563029 492452
rect 563229 493428 563287 493440
rect 563229 492452 563241 493428
rect 563275 492452 563287 493428
rect 563229 492440 563287 492452
rect 563487 493428 563545 493440
rect 563487 492452 563499 493428
rect 563533 492452 563545 493428
rect 563487 492440 563545 492452
rect 563745 493428 563803 493440
rect 563745 492452 563757 493428
rect 563791 492452 563803 493428
rect 563745 492440 563803 492452
rect 564003 493428 564061 493440
rect 564003 492452 564015 493428
rect 564049 492452 564061 493428
rect 564003 492440 564061 492452
rect 564261 493428 564319 493440
rect 564261 492452 564273 493428
rect 564307 492452 564319 493428
rect 564261 492440 564319 492452
rect 564519 493428 564577 493440
rect 564519 492452 564531 493428
rect 564565 492452 564577 493428
rect 564519 492440 564577 492452
rect 564777 493428 564835 493440
rect 564777 492452 564789 493428
rect 564823 492452 564835 493428
rect 564777 492440 564835 492452
rect 565035 493428 565093 493440
rect 565035 492452 565047 493428
rect 565081 492452 565093 493428
rect 565035 492440 565093 492452
rect 565293 493428 565351 493440
rect 565293 492452 565305 493428
rect 565339 492452 565351 493428
rect 565293 492440 565351 492452
rect 565551 493428 565609 493440
rect 565551 492452 565563 493428
rect 565597 492452 565609 493428
rect 565551 492440 565609 492452
rect 565809 493428 565867 493440
rect 565809 492452 565821 493428
rect 565855 492452 565867 493428
rect 565809 492440 565867 492452
rect 560585 404286 560643 404298
rect 560585 403310 560597 404286
rect 560631 403310 560643 404286
rect 560585 403298 560643 403310
rect 560843 404286 560901 404298
rect 560843 403310 560855 404286
rect 560889 403310 560901 404286
rect 560843 403298 560901 403310
rect 561101 404286 561159 404298
rect 561101 403310 561113 404286
rect 561147 403310 561159 404286
rect 561101 403298 561159 403310
rect 561359 404286 561417 404298
rect 561359 403310 561371 404286
rect 561405 403310 561417 404286
rect 561359 403298 561417 403310
rect 561617 404286 561675 404298
rect 561617 403310 561629 404286
rect 561663 403310 561675 404286
rect 561617 403298 561675 403310
rect 561875 404286 561933 404298
rect 561875 403310 561887 404286
rect 561921 403310 561933 404286
rect 561875 403298 561933 403310
rect 562133 404286 562191 404298
rect 562133 403310 562145 404286
rect 562179 403310 562191 404286
rect 562133 403298 562191 403310
rect 562391 404286 562449 404298
rect 562391 403310 562403 404286
rect 562437 403310 562449 404286
rect 562391 403298 562449 403310
rect 562649 404286 562707 404298
rect 562649 403310 562661 404286
rect 562695 403310 562707 404286
rect 562649 403298 562707 403310
rect 562907 404286 562965 404298
rect 562907 403310 562919 404286
rect 562953 403310 562965 404286
rect 562907 403298 562965 403310
rect 563165 404286 563223 404298
rect 563165 403310 563177 404286
rect 563211 403310 563223 404286
rect 563165 403298 563223 403310
rect 563423 404286 563481 404298
rect 563423 403310 563435 404286
rect 563469 403310 563481 404286
rect 563423 403298 563481 403310
rect 563681 404286 563739 404298
rect 563681 403310 563693 404286
rect 563727 403310 563739 404286
rect 563681 403298 563739 403310
rect 563939 404286 563997 404298
rect 563939 403310 563951 404286
rect 563985 403310 563997 404286
rect 563939 403298 563997 403310
rect 564197 404286 564255 404298
rect 564197 403310 564209 404286
rect 564243 403310 564255 404286
rect 564197 403298 564255 403310
rect 564455 404286 564513 404298
rect 564455 403310 564467 404286
rect 564501 403310 564513 404286
rect 564455 403298 564513 403310
rect 564713 404286 564771 404298
rect 564713 403310 564725 404286
rect 564759 403310 564771 404286
rect 564713 403298 564771 403310
rect 564971 404286 565029 404298
rect 564971 403310 564983 404286
rect 565017 403310 565029 404286
rect 564971 403298 565029 403310
rect 565229 404286 565287 404298
rect 565229 403310 565241 404286
rect 565275 403310 565287 404286
rect 565229 403298 565287 403310
rect 565487 404286 565545 404298
rect 565487 403310 565499 404286
rect 565533 403310 565545 404286
rect 565487 403298 565545 403310
rect 565745 404286 565803 404298
rect 565745 403310 565757 404286
rect 565791 403310 565803 404286
rect 565745 403298 565803 403310
rect 560541 358968 560599 358980
rect 560541 357992 560553 358968
rect 560587 357992 560599 358968
rect 560541 357980 560599 357992
rect 560799 358968 560857 358980
rect 560799 357992 560811 358968
rect 560845 357992 560857 358968
rect 560799 357980 560857 357992
rect 561057 358968 561115 358980
rect 561057 357992 561069 358968
rect 561103 357992 561115 358968
rect 561057 357980 561115 357992
rect 561315 358968 561373 358980
rect 561315 357992 561327 358968
rect 561361 357992 561373 358968
rect 561315 357980 561373 357992
rect 561573 358968 561631 358980
rect 561573 357992 561585 358968
rect 561619 357992 561631 358968
rect 561573 357980 561631 357992
rect 561831 358968 561889 358980
rect 561831 357992 561843 358968
rect 561877 357992 561889 358968
rect 561831 357980 561889 357992
rect 562089 358968 562147 358980
rect 562089 357992 562101 358968
rect 562135 357992 562147 358968
rect 562089 357980 562147 357992
rect 562347 358968 562405 358980
rect 562347 357992 562359 358968
rect 562393 357992 562405 358968
rect 562347 357980 562405 357992
rect 562605 358968 562663 358980
rect 562605 357992 562617 358968
rect 562651 357992 562663 358968
rect 562605 357980 562663 357992
rect 562863 358968 562921 358980
rect 562863 357992 562875 358968
rect 562909 357992 562921 358968
rect 562863 357980 562921 357992
rect 563121 358968 563179 358980
rect 563121 357992 563133 358968
rect 563167 357992 563179 358968
rect 563121 357980 563179 357992
rect 563379 358968 563437 358980
rect 563379 357992 563391 358968
rect 563425 357992 563437 358968
rect 563379 357980 563437 357992
rect 563637 358968 563695 358980
rect 563637 357992 563649 358968
rect 563683 357992 563695 358968
rect 563637 357980 563695 357992
rect 563895 358968 563953 358980
rect 563895 357992 563907 358968
rect 563941 357992 563953 358968
rect 563895 357980 563953 357992
rect 564153 358968 564211 358980
rect 564153 357992 564165 358968
rect 564199 357992 564211 358968
rect 564153 357980 564211 357992
rect 564411 358968 564469 358980
rect 564411 357992 564423 358968
rect 564457 357992 564469 358968
rect 564411 357980 564469 357992
rect 564669 358968 564727 358980
rect 564669 357992 564681 358968
rect 564715 357992 564727 358968
rect 564669 357980 564727 357992
rect 564927 358968 564985 358980
rect 564927 357992 564939 358968
rect 564973 357992 564985 358968
rect 564927 357980 564985 357992
rect 565185 358968 565243 358980
rect 565185 357992 565197 358968
rect 565231 357992 565243 358968
rect 565185 357980 565243 357992
rect 565443 358968 565501 358980
rect 565443 357992 565455 358968
rect 565489 357992 565501 358968
rect 565443 357980 565501 357992
rect 565701 358968 565759 358980
rect 565701 357992 565713 358968
rect 565747 357992 565759 358968
rect 565701 357980 565759 357992
rect 560403 312660 560461 312672
rect 560403 311684 560415 312660
rect 560449 311684 560461 312660
rect 560403 311672 560461 311684
rect 560661 312660 560719 312672
rect 560661 311684 560673 312660
rect 560707 311684 560719 312660
rect 560661 311672 560719 311684
rect 560919 312660 560977 312672
rect 560919 311684 560931 312660
rect 560965 311684 560977 312660
rect 560919 311672 560977 311684
rect 561177 312660 561235 312672
rect 561177 311684 561189 312660
rect 561223 311684 561235 312660
rect 561177 311672 561235 311684
rect 561435 312660 561493 312672
rect 561435 311684 561447 312660
rect 561481 311684 561493 312660
rect 561435 311672 561493 311684
rect 561693 312660 561751 312672
rect 561693 311684 561705 312660
rect 561739 311684 561751 312660
rect 561693 311672 561751 311684
rect 561951 312660 562009 312672
rect 561951 311684 561963 312660
rect 561997 311684 562009 312660
rect 561951 311672 562009 311684
rect 562209 312660 562267 312672
rect 562209 311684 562221 312660
rect 562255 311684 562267 312660
rect 562209 311672 562267 311684
rect 562467 312660 562525 312672
rect 562467 311684 562479 312660
rect 562513 311684 562525 312660
rect 562467 311672 562525 311684
rect 562725 312660 562783 312672
rect 562725 311684 562737 312660
rect 562771 311684 562783 312660
rect 562725 311672 562783 311684
rect 562983 312660 563041 312672
rect 562983 311684 562995 312660
rect 563029 311684 563041 312660
rect 562983 311672 563041 311684
rect 563241 312660 563299 312672
rect 563241 311684 563253 312660
rect 563287 311684 563299 312660
rect 563241 311672 563299 311684
rect 563499 312660 563557 312672
rect 563499 311684 563511 312660
rect 563545 311684 563557 312660
rect 563499 311672 563557 311684
rect 563757 312660 563815 312672
rect 563757 311684 563769 312660
rect 563803 311684 563815 312660
rect 563757 311672 563815 311684
rect 564015 312660 564073 312672
rect 564015 311684 564027 312660
rect 564061 311684 564073 312660
rect 564015 311672 564073 311684
rect 564273 312660 564331 312672
rect 564273 311684 564285 312660
rect 564319 311684 564331 312660
rect 564273 311672 564331 311684
rect 564531 312660 564589 312672
rect 564531 311684 564543 312660
rect 564577 311684 564589 312660
rect 564531 311672 564589 311684
rect 564789 312660 564847 312672
rect 564789 311684 564801 312660
rect 564835 311684 564847 312660
rect 564789 311672 564847 311684
rect 565047 312660 565105 312672
rect 565047 311684 565059 312660
rect 565093 311684 565105 312660
rect 565047 311672 565105 311684
rect 565305 312660 565363 312672
rect 565305 311684 565317 312660
rect 565351 311684 565363 312660
rect 565305 311672 565363 311684
rect 565563 312660 565621 312672
rect 565563 311684 565575 312660
rect 565609 311684 565621 312660
rect 565563 311672 565621 311684
<< pdiff >>
rect 575205 493202 575263 493214
rect 575205 492226 575217 493202
rect 575251 492226 575263 493202
rect 575205 492214 575263 492226
rect 575463 493202 575521 493214
rect 575463 492226 575475 493202
rect 575509 492226 575521 493202
rect 575463 492214 575521 492226
rect 575721 493202 575779 493214
rect 575721 492226 575733 493202
rect 575767 492226 575779 493202
rect 575721 492214 575779 492226
rect 575979 493202 576037 493214
rect 575979 492226 575991 493202
rect 576025 492226 576037 493202
rect 575979 492214 576037 492226
rect 576237 493202 576295 493214
rect 576237 492226 576249 493202
rect 576283 492226 576295 493202
rect 576237 492214 576295 492226
rect 576495 493202 576553 493214
rect 576495 492226 576507 493202
rect 576541 492226 576553 493202
rect 576495 492214 576553 492226
rect 576753 493202 576811 493214
rect 576753 492226 576765 493202
rect 576799 492226 576811 493202
rect 576753 492214 576811 492226
rect 577011 493202 577069 493214
rect 577011 492226 577023 493202
rect 577057 492226 577069 493202
rect 577011 492214 577069 492226
rect 577269 493202 577327 493214
rect 577269 492226 577281 493202
rect 577315 492226 577327 493202
rect 577269 492214 577327 492226
rect 577527 493202 577585 493214
rect 577527 492226 577539 493202
rect 577573 492226 577585 493202
rect 577527 492214 577585 492226
rect 577785 493202 577843 493214
rect 577785 492226 577797 493202
rect 577831 492226 577843 493202
rect 577785 492214 577843 492226
rect 578043 493202 578101 493214
rect 578043 492226 578055 493202
rect 578089 492226 578101 493202
rect 578043 492214 578101 492226
rect 578301 493202 578359 493214
rect 578301 492226 578313 493202
rect 578347 492226 578359 493202
rect 578301 492214 578359 492226
rect 578559 493202 578617 493214
rect 578559 492226 578571 493202
rect 578605 492226 578617 493202
rect 578559 492214 578617 492226
rect 578817 493202 578875 493214
rect 578817 492226 578829 493202
rect 578863 492226 578875 493202
rect 578817 492214 578875 492226
rect 579075 493202 579133 493214
rect 579075 492226 579087 493202
rect 579121 492226 579133 493202
rect 579075 492214 579133 492226
rect 579333 493202 579391 493214
rect 579333 492226 579345 493202
rect 579379 492226 579391 493202
rect 579333 492214 579391 492226
rect 579591 493202 579649 493214
rect 579591 492226 579603 493202
rect 579637 492226 579649 493202
rect 579591 492214 579649 492226
rect 579849 493202 579907 493214
rect 579849 492226 579861 493202
rect 579895 492226 579907 493202
rect 579849 492214 579907 492226
rect 580107 493202 580165 493214
rect 580107 492226 580119 493202
rect 580153 492226 580165 493202
rect 580107 492214 580165 492226
rect 580365 493202 580423 493214
rect 580365 492226 580377 493202
rect 580411 492226 580423 493202
rect 580365 492214 580423 492226
rect 574483 404326 574541 404338
rect 574483 403350 574495 404326
rect 574529 403350 574541 404326
rect 574483 403338 574541 403350
rect 574741 404326 574799 404338
rect 574741 403350 574753 404326
rect 574787 403350 574799 404326
rect 574741 403338 574799 403350
rect 574999 404326 575057 404338
rect 574999 403350 575011 404326
rect 575045 403350 575057 404326
rect 574999 403338 575057 403350
rect 575257 404326 575315 404338
rect 575257 403350 575269 404326
rect 575303 403350 575315 404326
rect 575257 403338 575315 403350
rect 575515 404326 575573 404338
rect 575515 403350 575527 404326
rect 575561 403350 575573 404326
rect 575515 403338 575573 403350
rect 575773 404326 575831 404338
rect 575773 403350 575785 404326
rect 575819 403350 575831 404326
rect 575773 403338 575831 403350
rect 576031 404326 576089 404338
rect 576031 403350 576043 404326
rect 576077 403350 576089 404326
rect 576031 403338 576089 403350
rect 576289 404326 576347 404338
rect 576289 403350 576301 404326
rect 576335 403350 576347 404326
rect 576289 403338 576347 403350
rect 576547 404326 576605 404338
rect 576547 403350 576559 404326
rect 576593 403350 576605 404326
rect 576547 403338 576605 403350
rect 576805 404326 576863 404338
rect 576805 403350 576817 404326
rect 576851 403350 576863 404326
rect 576805 403338 576863 403350
rect 577063 404326 577121 404338
rect 577063 403350 577075 404326
rect 577109 403350 577121 404326
rect 577063 403338 577121 403350
rect 577321 404326 577379 404338
rect 577321 403350 577333 404326
rect 577367 403350 577379 404326
rect 577321 403338 577379 403350
rect 577579 404326 577637 404338
rect 577579 403350 577591 404326
rect 577625 403350 577637 404326
rect 577579 403338 577637 403350
rect 577837 404326 577895 404338
rect 577837 403350 577849 404326
rect 577883 403350 577895 404326
rect 577837 403338 577895 403350
rect 578095 404326 578153 404338
rect 578095 403350 578107 404326
rect 578141 403350 578153 404326
rect 578095 403338 578153 403350
rect 578353 404326 578411 404338
rect 578353 403350 578365 404326
rect 578399 403350 578411 404326
rect 578353 403338 578411 403350
rect 578611 404326 578669 404338
rect 578611 403350 578623 404326
rect 578657 403350 578669 404326
rect 578611 403338 578669 403350
rect 578869 404326 578927 404338
rect 578869 403350 578881 404326
rect 578915 403350 578927 404326
rect 578869 403338 578927 403350
rect 579127 404326 579185 404338
rect 579127 403350 579139 404326
rect 579173 403350 579185 404326
rect 579127 403338 579185 403350
rect 579385 404326 579443 404338
rect 579385 403350 579397 404326
rect 579431 403350 579443 404326
rect 579385 403338 579443 403350
rect 579643 404326 579701 404338
rect 579643 403350 579655 404326
rect 579689 403350 579701 404326
rect 579643 403338 579701 403350
rect 574679 358898 574737 358910
rect 574679 357922 574691 358898
rect 574725 357922 574737 358898
rect 574679 357910 574737 357922
rect 574937 358898 574995 358910
rect 574937 357922 574949 358898
rect 574983 357922 574995 358898
rect 574937 357910 574995 357922
rect 575195 358898 575253 358910
rect 575195 357922 575207 358898
rect 575241 357922 575253 358898
rect 575195 357910 575253 357922
rect 575453 358898 575511 358910
rect 575453 357922 575465 358898
rect 575499 357922 575511 358898
rect 575453 357910 575511 357922
rect 575711 358898 575769 358910
rect 575711 357922 575723 358898
rect 575757 357922 575769 358898
rect 575711 357910 575769 357922
rect 575969 358898 576027 358910
rect 575969 357922 575981 358898
rect 576015 357922 576027 358898
rect 575969 357910 576027 357922
rect 576227 358898 576285 358910
rect 576227 357922 576239 358898
rect 576273 357922 576285 358898
rect 576227 357910 576285 357922
rect 576485 358898 576543 358910
rect 576485 357922 576497 358898
rect 576531 357922 576543 358898
rect 576485 357910 576543 357922
rect 576743 358898 576801 358910
rect 576743 357922 576755 358898
rect 576789 357922 576801 358898
rect 576743 357910 576801 357922
rect 577001 358898 577059 358910
rect 577001 357922 577013 358898
rect 577047 357922 577059 358898
rect 577001 357910 577059 357922
rect 577259 358898 577317 358910
rect 577259 357922 577271 358898
rect 577305 357922 577317 358898
rect 577259 357910 577317 357922
rect 577517 358898 577575 358910
rect 577517 357922 577529 358898
rect 577563 357922 577575 358898
rect 577517 357910 577575 357922
rect 577775 358898 577833 358910
rect 577775 357922 577787 358898
rect 577821 357922 577833 358898
rect 577775 357910 577833 357922
rect 578033 358898 578091 358910
rect 578033 357922 578045 358898
rect 578079 357922 578091 358898
rect 578033 357910 578091 357922
rect 578291 358898 578349 358910
rect 578291 357922 578303 358898
rect 578337 357922 578349 358898
rect 578291 357910 578349 357922
rect 578549 358898 578607 358910
rect 578549 357922 578561 358898
rect 578595 357922 578607 358898
rect 578549 357910 578607 357922
rect 578807 358898 578865 358910
rect 578807 357922 578819 358898
rect 578853 357922 578865 358898
rect 578807 357910 578865 357922
rect 579065 358898 579123 358910
rect 579065 357922 579077 358898
rect 579111 357922 579123 358898
rect 579065 357910 579123 357922
rect 579323 358898 579381 358910
rect 579323 357922 579335 358898
rect 579369 357922 579381 358898
rect 579323 357910 579381 357922
rect 579581 358898 579639 358910
rect 579581 357922 579593 358898
rect 579627 357922 579639 358898
rect 579581 357910 579639 357922
rect 579839 358898 579897 358910
rect 579839 357922 579851 358898
rect 579885 357922 579897 358898
rect 579839 357910 579897 357922
rect 575127 312730 575185 312742
rect 575127 311754 575139 312730
rect 575173 311754 575185 312730
rect 575127 311742 575185 311754
rect 575385 312730 575443 312742
rect 575385 311754 575397 312730
rect 575431 311754 575443 312730
rect 575385 311742 575443 311754
rect 575643 312730 575701 312742
rect 575643 311754 575655 312730
rect 575689 311754 575701 312730
rect 575643 311742 575701 311754
rect 575901 312730 575959 312742
rect 575901 311754 575913 312730
rect 575947 311754 575959 312730
rect 575901 311742 575959 311754
rect 576159 312730 576217 312742
rect 576159 311754 576171 312730
rect 576205 311754 576217 312730
rect 576159 311742 576217 311754
rect 576417 312730 576475 312742
rect 576417 311754 576429 312730
rect 576463 311754 576475 312730
rect 576417 311742 576475 311754
rect 576675 312730 576733 312742
rect 576675 311754 576687 312730
rect 576721 311754 576733 312730
rect 576675 311742 576733 311754
rect 576933 312730 576991 312742
rect 576933 311754 576945 312730
rect 576979 311754 576991 312730
rect 576933 311742 576991 311754
rect 577191 312730 577249 312742
rect 577191 311754 577203 312730
rect 577237 311754 577249 312730
rect 577191 311742 577249 311754
rect 577449 312730 577507 312742
rect 577449 311754 577461 312730
rect 577495 311754 577507 312730
rect 577449 311742 577507 311754
rect 577707 312730 577765 312742
rect 577707 311754 577719 312730
rect 577753 311754 577765 312730
rect 577707 311742 577765 311754
rect 577965 312730 578023 312742
rect 577965 311754 577977 312730
rect 578011 311754 578023 312730
rect 577965 311742 578023 311754
rect 578223 312730 578281 312742
rect 578223 311754 578235 312730
rect 578269 311754 578281 312730
rect 578223 311742 578281 311754
rect 578481 312730 578539 312742
rect 578481 311754 578493 312730
rect 578527 311754 578539 312730
rect 578481 311742 578539 311754
rect 578739 312730 578797 312742
rect 578739 311754 578751 312730
rect 578785 311754 578797 312730
rect 578739 311742 578797 311754
rect 578997 312730 579055 312742
rect 578997 311754 579009 312730
rect 579043 311754 579055 312730
rect 578997 311742 579055 311754
rect 579255 312730 579313 312742
rect 579255 311754 579267 312730
rect 579301 311754 579313 312730
rect 579255 311742 579313 311754
rect 579513 312730 579571 312742
rect 579513 311754 579525 312730
rect 579559 311754 579571 312730
rect 579513 311742 579571 311754
rect 579771 312730 579829 312742
rect 579771 311754 579783 312730
rect 579817 311754 579829 312730
rect 579771 311742 579829 311754
rect 580029 312730 580087 312742
rect 580029 311754 580041 312730
rect 580075 311754 580087 312730
rect 580029 311742 580087 311754
rect 580287 312730 580345 312742
rect 580287 311754 580299 312730
rect 580333 311754 580345 312730
rect 580287 311742 580345 311754
<< ndiffc >>
rect 560661 492452 560695 493428
rect 560919 492452 560953 493428
rect 561177 492452 561211 493428
rect 561435 492452 561469 493428
rect 561693 492452 561727 493428
rect 561951 492452 561985 493428
rect 562209 492452 562243 493428
rect 562467 492452 562501 493428
rect 562725 492452 562759 493428
rect 562983 492452 563017 493428
rect 563241 492452 563275 493428
rect 563499 492452 563533 493428
rect 563757 492452 563791 493428
rect 564015 492452 564049 493428
rect 564273 492452 564307 493428
rect 564531 492452 564565 493428
rect 564789 492452 564823 493428
rect 565047 492452 565081 493428
rect 565305 492452 565339 493428
rect 565563 492452 565597 493428
rect 565821 492452 565855 493428
rect 560597 403310 560631 404286
rect 560855 403310 560889 404286
rect 561113 403310 561147 404286
rect 561371 403310 561405 404286
rect 561629 403310 561663 404286
rect 561887 403310 561921 404286
rect 562145 403310 562179 404286
rect 562403 403310 562437 404286
rect 562661 403310 562695 404286
rect 562919 403310 562953 404286
rect 563177 403310 563211 404286
rect 563435 403310 563469 404286
rect 563693 403310 563727 404286
rect 563951 403310 563985 404286
rect 564209 403310 564243 404286
rect 564467 403310 564501 404286
rect 564725 403310 564759 404286
rect 564983 403310 565017 404286
rect 565241 403310 565275 404286
rect 565499 403310 565533 404286
rect 565757 403310 565791 404286
rect 560553 357992 560587 358968
rect 560811 357992 560845 358968
rect 561069 357992 561103 358968
rect 561327 357992 561361 358968
rect 561585 357992 561619 358968
rect 561843 357992 561877 358968
rect 562101 357992 562135 358968
rect 562359 357992 562393 358968
rect 562617 357992 562651 358968
rect 562875 357992 562909 358968
rect 563133 357992 563167 358968
rect 563391 357992 563425 358968
rect 563649 357992 563683 358968
rect 563907 357992 563941 358968
rect 564165 357992 564199 358968
rect 564423 357992 564457 358968
rect 564681 357992 564715 358968
rect 564939 357992 564973 358968
rect 565197 357992 565231 358968
rect 565455 357992 565489 358968
rect 565713 357992 565747 358968
rect 560415 311684 560449 312660
rect 560673 311684 560707 312660
rect 560931 311684 560965 312660
rect 561189 311684 561223 312660
rect 561447 311684 561481 312660
rect 561705 311684 561739 312660
rect 561963 311684 561997 312660
rect 562221 311684 562255 312660
rect 562479 311684 562513 312660
rect 562737 311684 562771 312660
rect 562995 311684 563029 312660
rect 563253 311684 563287 312660
rect 563511 311684 563545 312660
rect 563769 311684 563803 312660
rect 564027 311684 564061 312660
rect 564285 311684 564319 312660
rect 564543 311684 564577 312660
rect 564801 311684 564835 312660
rect 565059 311684 565093 312660
rect 565317 311684 565351 312660
rect 565575 311684 565609 312660
<< pdiffc >>
rect 575217 492226 575251 493202
rect 575475 492226 575509 493202
rect 575733 492226 575767 493202
rect 575991 492226 576025 493202
rect 576249 492226 576283 493202
rect 576507 492226 576541 493202
rect 576765 492226 576799 493202
rect 577023 492226 577057 493202
rect 577281 492226 577315 493202
rect 577539 492226 577573 493202
rect 577797 492226 577831 493202
rect 578055 492226 578089 493202
rect 578313 492226 578347 493202
rect 578571 492226 578605 493202
rect 578829 492226 578863 493202
rect 579087 492226 579121 493202
rect 579345 492226 579379 493202
rect 579603 492226 579637 493202
rect 579861 492226 579895 493202
rect 580119 492226 580153 493202
rect 580377 492226 580411 493202
rect 574495 403350 574529 404326
rect 574753 403350 574787 404326
rect 575011 403350 575045 404326
rect 575269 403350 575303 404326
rect 575527 403350 575561 404326
rect 575785 403350 575819 404326
rect 576043 403350 576077 404326
rect 576301 403350 576335 404326
rect 576559 403350 576593 404326
rect 576817 403350 576851 404326
rect 577075 403350 577109 404326
rect 577333 403350 577367 404326
rect 577591 403350 577625 404326
rect 577849 403350 577883 404326
rect 578107 403350 578141 404326
rect 578365 403350 578399 404326
rect 578623 403350 578657 404326
rect 578881 403350 578915 404326
rect 579139 403350 579173 404326
rect 579397 403350 579431 404326
rect 579655 403350 579689 404326
rect 574691 357922 574725 358898
rect 574949 357922 574983 358898
rect 575207 357922 575241 358898
rect 575465 357922 575499 358898
rect 575723 357922 575757 358898
rect 575981 357922 576015 358898
rect 576239 357922 576273 358898
rect 576497 357922 576531 358898
rect 576755 357922 576789 358898
rect 577013 357922 577047 358898
rect 577271 357922 577305 358898
rect 577529 357922 577563 358898
rect 577787 357922 577821 358898
rect 578045 357922 578079 358898
rect 578303 357922 578337 358898
rect 578561 357922 578595 358898
rect 578819 357922 578853 358898
rect 579077 357922 579111 358898
rect 579335 357922 579369 358898
rect 579593 357922 579627 358898
rect 579851 357922 579885 358898
rect 575139 311754 575173 312730
rect 575397 311754 575431 312730
rect 575655 311754 575689 312730
rect 575913 311754 575947 312730
rect 576171 311754 576205 312730
rect 576429 311754 576463 312730
rect 576687 311754 576721 312730
rect 576945 311754 576979 312730
rect 577203 311754 577237 312730
rect 577461 311754 577495 312730
rect 577719 311754 577753 312730
rect 577977 311754 578011 312730
rect 578235 311754 578269 312730
rect 578493 311754 578527 312730
rect 578751 311754 578785 312730
rect 579009 311754 579043 312730
rect 579267 311754 579301 312730
rect 579525 311754 579559 312730
rect 579783 311754 579817 312730
rect 580041 311754 580075 312730
rect 580299 311754 580333 312730
<< psubdiff >>
rect 565886 492100 565926 492140
rect 562148 492068 562268 492070
rect 562148 492032 562184 492068
rect 562228 492032 562268 492068
rect 562148 492020 562268 492032
rect 563448 492068 563568 492070
rect 563448 492032 563484 492068
rect 563528 492032 563568 492068
rect 563448 492020 563568 492032
rect 564748 492068 564868 492070
rect 564748 492032 564784 492068
rect 564828 492032 564868 492068
rect 564748 492020 564868 492032
rect 565886 492020 565926 492060
rect 565822 402958 565862 402998
rect 562084 402926 562204 402928
rect 562084 402890 562120 402926
rect 562164 402890 562204 402926
rect 562084 402878 562204 402890
rect 563384 402926 563504 402928
rect 563384 402890 563420 402926
rect 563464 402890 563504 402926
rect 563384 402878 563504 402890
rect 564684 402926 564804 402928
rect 564684 402890 564720 402926
rect 564764 402890 564804 402926
rect 564684 402878 564804 402890
rect 565822 402878 565862 402918
rect 565778 357640 565818 357680
rect 562040 357608 562160 357610
rect 562040 357572 562076 357608
rect 562120 357572 562160 357608
rect 562040 357560 562160 357572
rect 563340 357608 563460 357610
rect 563340 357572 563376 357608
rect 563420 357572 563460 357608
rect 563340 357560 563460 357572
rect 564640 357608 564760 357610
rect 564640 357572 564676 357608
rect 564720 357572 564760 357608
rect 564640 357560 564760 357572
rect 565778 357560 565818 357600
rect 565640 311332 565680 311372
rect 561902 311300 562022 311302
rect 561902 311264 561938 311300
rect 561982 311264 562022 311300
rect 561902 311252 562022 311264
rect 563202 311300 563322 311302
rect 563202 311264 563238 311300
rect 563282 311264 563322 311300
rect 563202 311252 563322 311264
rect 564502 311300 564622 311302
rect 564502 311264 564538 311300
rect 564582 311264 564622 311300
rect 564502 311252 564622 311264
rect 565640 311252 565680 311292
<< nsubdiff >>
rect 576740 493522 576860 493524
rect 576740 493486 576776 493522
rect 576820 493486 576860 493522
rect 576740 493484 576860 493486
rect 578040 493522 578160 493524
rect 578040 493486 578076 493522
rect 578120 493486 578160 493522
rect 578040 493484 578160 493486
rect 579340 493522 579460 493524
rect 579340 493486 579376 493522
rect 579420 493486 579460 493522
rect 579340 493484 579460 493486
rect 580478 493474 580518 493514
rect 580478 493394 580518 493434
rect 576018 404646 576138 404648
rect 576018 404610 576054 404646
rect 576098 404610 576138 404646
rect 576018 404608 576138 404610
rect 577318 404646 577438 404648
rect 577318 404610 577354 404646
rect 577398 404610 577438 404646
rect 577318 404608 577438 404610
rect 578618 404646 578738 404648
rect 578618 404610 578654 404646
rect 578698 404610 578738 404646
rect 578618 404608 578738 404610
rect 579756 404598 579796 404638
rect 579756 404518 579796 404558
rect 576214 359218 576334 359220
rect 576214 359182 576250 359218
rect 576294 359182 576334 359218
rect 576214 359180 576334 359182
rect 577514 359218 577634 359220
rect 577514 359182 577550 359218
rect 577594 359182 577634 359218
rect 577514 359180 577634 359182
rect 578814 359218 578934 359220
rect 578814 359182 578850 359218
rect 578894 359182 578934 359218
rect 578814 359180 578934 359182
rect 579952 359170 579992 359210
rect 579952 359090 579992 359130
rect 576662 313050 576782 313052
rect 576662 313014 576698 313050
rect 576742 313014 576782 313050
rect 576662 313012 576782 313014
rect 577962 313050 578082 313052
rect 577962 313014 577998 313050
rect 578042 313014 578082 313050
rect 577962 313012 578082 313014
rect 579262 313050 579382 313052
rect 579262 313014 579298 313050
rect 579342 313014 579382 313050
rect 579262 313012 579382 313014
rect 580400 313002 580440 313042
rect 580400 312922 580440 312962
<< psubdiffcont >>
rect 562184 492032 562228 492068
rect 563484 492032 563528 492068
rect 564784 492032 564828 492068
rect 565886 492060 565926 492100
rect 562120 402890 562164 402926
rect 563420 402890 563464 402926
rect 564720 402890 564764 402926
rect 565822 402918 565862 402958
rect 562076 357572 562120 357608
rect 563376 357572 563420 357608
rect 564676 357572 564720 357608
rect 565778 357600 565818 357640
rect 561938 311264 561982 311300
rect 563238 311264 563282 311300
rect 564538 311264 564582 311300
rect 565640 311292 565680 311332
<< nsubdiffcont >>
rect 576776 493486 576820 493522
rect 578076 493486 578120 493522
rect 579376 493486 579420 493522
rect 580478 493434 580518 493474
rect 576054 404610 576098 404646
rect 577354 404610 577398 404646
rect 578654 404610 578698 404646
rect 579756 404558 579796 404598
rect 576250 359182 576294 359218
rect 577550 359182 577594 359218
rect 578850 359182 578894 359218
rect 579952 359130 579992 359170
rect 576698 313014 576742 313050
rect 577998 313014 578042 313050
rect 579298 313014 579342 313050
rect 580400 312962 580440 313002
<< poly >>
rect 560707 493440 560907 493466
rect 560965 493440 561165 493466
rect 561223 493440 561423 493466
rect 561481 493440 561681 493466
rect 561739 493440 561939 493466
rect 561997 493440 562197 493466
rect 562255 493440 562455 493466
rect 562513 493440 562713 493466
rect 562771 493440 562971 493466
rect 563029 493440 563229 493466
rect 563287 493440 563487 493466
rect 563545 493440 563745 493466
rect 563803 493440 564003 493466
rect 564061 493440 564261 493466
rect 564319 493440 564519 493466
rect 564577 493440 564777 493466
rect 564835 493440 565035 493466
rect 565093 493440 565293 493466
rect 565351 493440 565551 493466
rect 565609 493440 565809 493466
rect 575263 493214 575463 493240
rect 575521 493214 575721 493240
rect 575779 493214 575979 493240
rect 576037 493214 576237 493240
rect 576295 493214 576495 493240
rect 576553 493214 576753 493240
rect 576811 493214 577011 493240
rect 577069 493214 577269 493240
rect 577327 493214 577527 493240
rect 577585 493214 577785 493240
rect 577843 493214 578043 493240
rect 578101 493214 578301 493240
rect 578359 493214 578559 493240
rect 578617 493214 578817 493240
rect 578875 493214 579075 493240
rect 579133 493214 579333 493240
rect 579391 493214 579591 493240
rect 579649 493214 579849 493240
rect 579907 493214 580107 493240
rect 580165 493214 580365 493240
rect 560707 492414 560907 492440
rect 560965 492414 561165 492440
rect 561223 492414 561423 492440
rect 561481 492414 561681 492440
rect 561739 492414 561939 492440
rect 561997 492414 562197 492440
rect 562255 492414 562455 492440
rect 562513 492414 562713 492440
rect 562771 492414 562971 492440
rect 563029 492414 563229 492440
rect 563287 492414 563487 492440
rect 563545 492414 563745 492440
rect 563803 492414 564003 492440
rect 564061 492414 564261 492440
rect 564319 492414 564519 492440
rect 564577 492414 564777 492440
rect 564835 492414 565035 492440
rect 565093 492414 565293 492440
rect 565351 492414 565551 492440
rect 565609 492414 565809 492440
rect 560762 492224 560882 492414
rect 561018 492224 561138 492414
rect 561274 492224 561394 492414
rect 561530 492224 561650 492414
rect 561786 492224 561906 492414
rect 562042 492224 562162 492414
rect 562298 492224 562418 492414
rect 562554 492224 562674 492414
rect 562810 492224 562930 492414
rect 563066 492224 563186 492414
rect 563322 492224 563442 492414
rect 563578 492224 563698 492414
rect 563834 492224 563954 492414
rect 564090 492224 564210 492414
rect 564346 492224 564466 492414
rect 564602 492224 564722 492414
rect 564858 492224 564978 492414
rect 565114 492224 565234 492414
rect 565370 492224 565490 492414
rect 565626 492224 565746 492414
rect 560650 492204 565786 492224
rect 560650 492144 560836 492204
rect 560896 492144 561036 492204
rect 561096 492144 561236 492204
rect 561296 492144 561436 492204
rect 561496 492144 561636 492204
rect 561696 492144 561836 492204
rect 561896 492144 562036 492204
rect 562096 492144 562236 492204
rect 562296 492144 562436 492204
rect 562496 492144 562636 492204
rect 562696 492144 562836 492204
rect 562896 492144 563036 492204
rect 563096 492144 563236 492204
rect 563296 492144 563436 492204
rect 563496 492144 563636 492204
rect 563696 492144 563836 492204
rect 563896 492144 564036 492204
rect 564096 492144 564236 492204
rect 564296 492144 564436 492204
rect 564496 492144 564636 492204
rect 564696 492144 564836 492204
rect 564896 492144 565036 492204
rect 565096 492144 565236 492204
rect 565296 492144 565436 492204
rect 565496 492144 565636 492204
rect 565696 492144 565786 492204
rect 575263 492188 575463 492214
rect 575521 492188 575721 492214
rect 575779 492188 575979 492214
rect 576037 492188 576237 492214
rect 576295 492188 576495 492214
rect 576553 492188 576753 492214
rect 576811 492188 577011 492214
rect 577069 492188 577269 492214
rect 577327 492188 577527 492214
rect 577585 492188 577785 492214
rect 577843 492188 578043 492214
rect 578101 492188 578301 492214
rect 578359 492188 578559 492214
rect 578617 492188 578817 492214
rect 578875 492188 579075 492214
rect 579133 492188 579333 492214
rect 579391 492188 579591 492214
rect 579649 492188 579849 492214
rect 579907 492188 580107 492214
rect 580165 492188 580365 492214
rect 560650 492124 565786 492144
rect 575334 491942 575454 492188
rect 575590 491942 575710 492188
rect 575846 491942 575966 492188
rect 576102 491942 576222 492188
rect 576358 491942 576478 492188
rect 576614 491942 576734 492188
rect 576870 491942 576990 492188
rect 577126 491942 577246 492188
rect 577382 491942 577502 492188
rect 577638 491942 577758 492188
rect 577894 491942 578014 492188
rect 578150 491942 578270 492188
rect 578406 491942 578526 492188
rect 578662 491942 578782 492188
rect 578918 491942 579038 492188
rect 579174 491942 579294 492188
rect 579430 491942 579550 492188
rect 579686 491942 579806 492188
rect 579942 491942 580062 492188
rect 580198 491942 580318 492188
rect 575170 491922 580458 491942
rect 575170 491862 575228 491922
rect 575288 491862 575428 491922
rect 575488 491862 575628 491922
rect 575688 491862 575828 491922
rect 575888 491862 576028 491922
rect 576088 491862 576228 491922
rect 576288 491862 576428 491922
rect 576488 491862 576628 491922
rect 576688 491862 576828 491922
rect 576888 491862 577028 491922
rect 577088 491862 577228 491922
rect 577288 491862 577428 491922
rect 577488 491862 577628 491922
rect 577688 491862 577828 491922
rect 577888 491862 578028 491922
rect 578088 491862 578228 491922
rect 578288 491862 578428 491922
rect 578488 491862 578628 491922
rect 578688 491862 578828 491922
rect 578888 491862 579028 491922
rect 579088 491862 579228 491922
rect 579288 491862 579428 491922
rect 579488 491862 579628 491922
rect 579688 491862 579828 491922
rect 579888 491862 580028 491922
rect 580088 491862 580228 491922
rect 580288 491862 580458 491922
rect 575170 491842 580458 491862
rect 574541 404338 574741 404364
rect 574799 404338 574999 404364
rect 575057 404338 575257 404364
rect 575315 404338 575515 404364
rect 575573 404338 575773 404364
rect 575831 404338 576031 404364
rect 576089 404338 576289 404364
rect 576347 404338 576547 404364
rect 576605 404338 576805 404364
rect 576863 404338 577063 404364
rect 577121 404338 577321 404364
rect 577379 404338 577579 404364
rect 577637 404338 577837 404364
rect 577895 404338 578095 404364
rect 578153 404338 578353 404364
rect 578411 404338 578611 404364
rect 578669 404338 578869 404364
rect 578927 404338 579127 404364
rect 579185 404338 579385 404364
rect 579443 404338 579643 404364
rect 560643 404298 560843 404324
rect 560901 404298 561101 404324
rect 561159 404298 561359 404324
rect 561417 404298 561617 404324
rect 561675 404298 561875 404324
rect 561933 404298 562133 404324
rect 562191 404298 562391 404324
rect 562449 404298 562649 404324
rect 562707 404298 562907 404324
rect 562965 404298 563165 404324
rect 563223 404298 563423 404324
rect 563481 404298 563681 404324
rect 563739 404298 563939 404324
rect 563997 404298 564197 404324
rect 564255 404298 564455 404324
rect 564513 404298 564713 404324
rect 564771 404298 564971 404324
rect 565029 404298 565229 404324
rect 565287 404298 565487 404324
rect 565545 404298 565745 404324
rect 574541 403312 574741 403338
rect 574799 403312 574999 403338
rect 575057 403312 575257 403338
rect 575315 403312 575515 403338
rect 575573 403312 575773 403338
rect 575831 403312 576031 403338
rect 576089 403312 576289 403338
rect 576347 403312 576547 403338
rect 576605 403312 576805 403338
rect 576863 403312 577063 403338
rect 577121 403312 577321 403338
rect 577379 403312 577579 403338
rect 577637 403312 577837 403338
rect 577895 403312 578095 403338
rect 578153 403312 578353 403338
rect 578411 403312 578611 403338
rect 578669 403312 578869 403338
rect 578927 403312 579127 403338
rect 579185 403312 579385 403338
rect 579443 403312 579643 403338
rect 560643 403272 560843 403298
rect 560901 403272 561101 403298
rect 561159 403272 561359 403298
rect 561417 403272 561617 403298
rect 561675 403272 561875 403298
rect 561933 403272 562133 403298
rect 562191 403272 562391 403298
rect 562449 403272 562649 403298
rect 562707 403272 562907 403298
rect 562965 403272 563165 403298
rect 563223 403272 563423 403298
rect 563481 403272 563681 403298
rect 563739 403272 563939 403298
rect 563997 403272 564197 403298
rect 564255 403272 564455 403298
rect 564513 403272 564713 403298
rect 564771 403272 564971 403298
rect 565029 403272 565229 403298
rect 565287 403272 565487 403298
rect 565545 403272 565745 403298
rect 560698 403082 560818 403272
rect 560954 403082 561074 403272
rect 561210 403082 561330 403272
rect 561466 403082 561586 403272
rect 561722 403082 561842 403272
rect 561978 403082 562098 403272
rect 562234 403082 562354 403272
rect 562490 403082 562610 403272
rect 562746 403082 562866 403272
rect 563002 403082 563122 403272
rect 563258 403082 563378 403272
rect 563514 403082 563634 403272
rect 563770 403082 563890 403272
rect 564026 403082 564146 403272
rect 564282 403082 564402 403272
rect 564538 403082 564658 403272
rect 564794 403082 564914 403272
rect 565050 403082 565170 403272
rect 565306 403082 565426 403272
rect 565562 403082 565682 403272
rect 560586 403062 565722 403082
rect 574612 403066 574732 403312
rect 574868 403066 574988 403312
rect 575124 403066 575244 403312
rect 575380 403066 575500 403312
rect 575636 403066 575756 403312
rect 575892 403066 576012 403312
rect 576148 403066 576268 403312
rect 576404 403066 576524 403312
rect 576660 403066 576780 403312
rect 576916 403066 577036 403312
rect 577172 403066 577292 403312
rect 577428 403066 577548 403312
rect 577684 403066 577804 403312
rect 577940 403066 578060 403312
rect 578196 403066 578316 403312
rect 578452 403066 578572 403312
rect 578708 403066 578828 403312
rect 578964 403066 579084 403312
rect 579220 403066 579340 403312
rect 579476 403066 579596 403312
rect 560586 403002 560772 403062
rect 560832 403002 560972 403062
rect 561032 403002 561172 403062
rect 561232 403002 561372 403062
rect 561432 403002 561572 403062
rect 561632 403002 561772 403062
rect 561832 403002 561972 403062
rect 562032 403002 562172 403062
rect 562232 403002 562372 403062
rect 562432 403002 562572 403062
rect 562632 403002 562772 403062
rect 562832 403002 562972 403062
rect 563032 403002 563172 403062
rect 563232 403002 563372 403062
rect 563432 403002 563572 403062
rect 563632 403002 563772 403062
rect 563832 403002 563972 403062
rect 564032 403002 564172 403062
rect 564232 403002 564372 403062
rect 564432 403002 564572 403062
rect 564632 403002 564772 403062
rect 564832 403002 564972 403062
rect 565032 403002 565172 403062
rect 565232 403002 565372 403062
rect 565432 403002 565572 403062
rect 565632 403002 565722 403062
rect 560586 402982 565722 403002
rect 574448 403046 579736 403066
rect 574448 402986 574506 403046
rect 574566 402986 574706 403046
rect 574766 402986 574906 403046
rect 574966 402986 575106 403046
rect 575166 402986 575306 403046
rect 575366 402986 575506 403046
rect 575566 402986 575706 403046
rect 575766 402986 575906 403046
rect 575966 402986 576106 403046
rect 576166 402986 576306 403046
rect 576366 402986 576506 403046
rect 576566 402986 576706 403046
rect 576766 402986 576906 403046
rect 576966 402986 577106 403046
rect 577166 402986 577306 403046
rect 577366 402986 577506 403046
rect 577566 402986 577706 403046
rect 577766 402986 577906 403046
rect 577966 402986 578106 403046
rect 578166 402986 578306 403046
rect 578366 402986 578506 403046
rect 578566 402986 578706 403046
rect 578766 402986 578906 403046
rect 578966 402986 579106 403046
rect 579166 402986 579306 403046
rect 579366 402986 579506 403046
rect 579566 402986 579736 403046
rect 574448 402966 579736 402986
rect 560599 358980 560799 359006
rect 560857 358980 561057 359006
rect 561115 358980 561315 359006
rect 561373 358980 561573 359006
rect 561631 358980 561831 359006
rect 561889 358980 562089 359006
rect 562147 358980 562347 359006
rect 562405 358980 562605 359006
rect 562663 358980 562863 359006
rect 562921 358980 563121 359006
rect 563179 358980 563379 359006
rect 563437 358980 563637 359006
rect 563695 358980 563895 359006
rect 563953 358980 564153 359006
rect 564211 358980 564411 359006
rect 564469 358980 564669 359006
rect 564727 358980 564927 359006
rect 564985 358980 565185 359006
rect 565243 358980 565443 359006
rect 565501 358980 565701 359006
rect 574737 358910 574937 358936
rect 574995 358910 575195 358936
rect 575253 358910 575453 358936
rect 575511 358910 575711 358936
rect 575769 358910 575969 358936
rect 576027 358910 576227 358936
rect 576285 358910 576485 358936
rect 576543 358910 576743 358936
rect 576801 358910 577001 358936
rect 577059 358910 577259 358936
rect 577317 358910 577517 358936
rect 577575 358910 577775 358936
rect 577833 358910 578033 358936
rect 578091 358910 578291 358936
rect 578349 358910 578549 358936
rect 578607 358910 578807 358936
rect 578865 358910 579065 358936
rect 579123 358910 579323 358936
rect 579381 358910 579581 358936
rect 579639 358910 579839 358936
rect 560599 357954 560799 357980
rect 560857 357954 561057 357980
rect 561115 357954 561315 357980
rect 561373 357954 561573 357980
rect 561631 357954 561831 357980
rect 561889 357954 562089 357980
rect 562147 357954 562347 357980
rect 562405 357954 562605 357980
rect 562663 357954 562863 357980
rect 562921 357954 563121 357980
rect 563179 357954 563379 357980
rect 563437 357954 563637 357980
rect 563695 357954 563895 357980
rect 563953 357954 564153 357980
rect 564211 357954 564411 357980
rect 564469 357954 564669 357980
rect 564727 357954 564927 357980
rect 564985 357954 565185 357980
rect 565243 357954 565443 357980
rect 565501 357954 565701 357980
rect 560654 357764 560774 357954
rect 560910 357764 561030 357954
rect 561166 357764 561286 357954
rect 561422 357764 561542 357954
rect 561678 357764 561798 357954
rect 561934 357764 562054 357954
rect 562190 357764 562310 357954
rect 562446 357764 562566 357954
rect 562702 357764 562822 357954
rect 562958 357764 563078 357954
rect 563214 357764 563334 357954
rect 563470 357764 563590 357954
rect 563726 357764 563846 357954
rect 563982 357764 564102 357954
rect 564238 357764 564358 357954
rect 564494 357764 564614 357954
rect 564750 357764 564870 357954
rect 565006 357764 565126 357954
rect 565262 357764 565382 357954
rect 565518 357764 565638 357954
rect 574737 357884 574937 357910
rect 574995 357884 575195 357910
rect 575253 357884 575453 357910
rect 575511 357884 575711 357910
rect 575769 357884 575969 357910
rect 576027 357884 576227 357910
rect 576285 357884 576485 357910
rect 576543 357884 576743 357910
rect 576801 357884 577001 357910
rect 577059 357884 577259 357910
rect 577317 357884 577517 357910
rect 577575 357884 577775 357910
rect 577833 357884 578033 357910
rect 578091 357884 578291 357910
rect 578349 357884 578549 357910
rect 578607 357884 578807 357910
rect 578865 357884 579065 357910
rect 579123 357884 579323 357910
rect 579381 357884 579581 357910
rect 579639 357884 579839 357910
rect 560542 357744 565678 357764
rect 560542 357684 560728 357744
rect 560788 357684 560928 357744
rect 560988 357684 561128 357744
rect 561188 357684 561328 357744
rect 561388 357684 561528 357744
rect 561588 357684 561728 357744
rect 561788 357684 561928 357744
rect 561988 357684 562128 357744
rect 562188 357684 562328 357744
rect 562388 357684 562528 357744
rect 562588 357684 562728 357744
rect 562788 357684 562928 357744
rect 562988 357684 563128 357744
rect 563188 357684 563328 357744
rect 563388 357684 563528 357744
rect 563588 357684 563728 357744
rect 563788 357684 563928 357744
rect 563988 357684 564128 357744
rect 564188 357684 564328 357744
rect 564388 357684 564528 357744
rect 564588 357684 564728 357744
rect 564788 357684 564928 357744
rect 564988 357684 565128 357744
rect 565188 357684 565328 357744
rect 565388 357684 565528 357744
rect 565588 357684 565678 357744
rect 560542 357664 565678 357684
rect 574808 357638 574928 357884
rect 575064 357638 575184 357884
rect 575320 357638 575440 357884
rect 575576 357638 575696 357884
rect 575832 357638 575952 357884
rect 576088 357638 576208 357884
rect 576344 357638 576464 357884
rect 576600 357638 576720 357884
rect 576856 357638 576976 357884
rect 577112 357638 577232 357884
rect 577368 357638 577488 357884
rect 577624 357638 577744 357884
rect 577880 357638 578000 357884
rect 578136 357638 578256 357884
rect 578392 357638 578512 357884
rect 578648 357638 578768 357884
rect 578904 357638 579024 357884
rect 579160 357638 579280 357884
rect 579416 357638 579536 357884
rect 579672 357638 579792 357884
rect 574644 357618 579932 357638
rect 574644 357558 574702 357618
rect 574762 357558 574902 357618
rect 574962 357558 575102 357618
rect 575162 357558 575302 357618
rect 575362 357558 575502 357618
rect 575562 357558 575702 357618
rect 575762 357558 575902 357618
rect 575962 357558 576102 357618
rect 576162 357558 576302 357618
rect 576362 357558 576502 357618
rect 576562 357558 576702 357618
rect 576762 357558 576902 357618
rect 576962 357558 577102 357618
rect 577162 357558 577302 357618
rect 577362 357558 577502 357618
rect 577562 357558 577702 357618
rect 577762 357558 577902 357618
rect 577962 357558 578102 357618
rect 578162 357558 578302 357618
rect 578362 357558 578502 357618
rect 578562 357558 578702 357618
rect 578762 357558 578902 357618
rect 578962 357558 579102 357618
rect 579162 357558 579302 357618
rect 579362 357558 579502 357618
rect 579562 357558 579702 357618
rect 579762 357558 579932 357618
rect 574644 357538 579932 357558
rect 575185 312742 575385 312768
rect 575443 312742 575643 312768
rect 575701 312742 575901 312768
rect 575959 312742 576159 312768
rect 576217 312742 576417 312768
rect 576475 312742 576675 312768
rect 576733 312742 576933 312768
rect 576991 312742 577191 312768
rect 577249 312742 577449 312768
rect 577507 312742 577707 312768
rect 577765 312742 577965 312768
rect 578023 312742 578223 312768
rect 578281 312742 578481 312768
rect 578539 312742 578739 312768
rect 578797 312742 578997 312768
rect 579055 312742 579255 312768
rect 579313 312742 579513 312768
rect 579571 312742 579771 312768
rect 579829 312742 580029 312768
rect 580087 312742 580287 312768
rect 560461 312672 560661 312698
rect 560719 312672 560919 312698
rect 560977 312672 561177 312698
rect 561235 312672 561435 312698
rect 561493 312672 561693 312698
rect 561751 312672 561951 312698
rect 562009 312672 562209 312698
rect 562267 312672 562467 312698
rect 562525 312672 562725 312698
rect 562783 312672 562983 312698
rect 563041 312672 563241 312698
rect 563299 312672 563499 312698
rect 563557 312672 563757 312698
rect 563815 312672 564015 312698
rect 564073 312672 564273 312698
rect 564331 312672 564531 312698
rect 564589 312672 564789 312698
rect 564847 312672 565047 312698
rect 565105 312672 565305 312698
rect 565363 312672 565563 312698
rect 575185 311716 575385 311742
rect 575443 311716 575643 311742
rect 575701 311716 575901 311742
rect 575959 311716 576159 311742
rect 576217 311716 576417 311742
rect 576475 311716 576675 311742
rect 576733 311716 576933 311742
rect 576991 311716 577191 311742
rect 577249 311716 577449 311742
rect 577507 311716 577707 311742
rect 577765 311716 577965 311742
rect 578023 311716 578223 311742
rect 578281 311716 578481 311742
rect 578539 311716 578739 311742
rect 578797 311716 578997 311742
rect 579055 311716 579255 311742
rect 579313 311716 579513 311742
rect 579571 311716 579771 311742
rect 579829 311716 580029 311742
rect 580087 311716 580287 311742
rect 560461 311646 560661 311672
rect 560719 311646 560919 311672
rect 560977 311646 561177 311672
rect 561235 311646 561435 311672
rect 561493 311646 561693 311672
rect 561751 311646 561951 311672
rect 562009 311646 562209 311672
rect 562267 311646 562467 311672
rect 562525 311646 562725 311672
rect 562783 311646 562983 311672
rect 563041 311646 563241 311672
rect 563299 311646 563499 311672
rect 563557 311646 563757 311672
rect 563815 311646 564015 311672
rect 564073 311646 564273 311672
rect 564331 311646 564531 311672
rect 564589 311646 564789 311672
rect 564847 311646 565047 311672
rect 565105 311646 565305 311672
rect 565363 311646 565563 311672
rect 560516 311456 560636 311646
rect 560772 311456 560892 311646
rect 561028 311456 561148 311646
rect 561284 311456 561404 311646
rect 561540 311456 561660 311646
rect 561796 311456 561916 311646
rect 562052 311456 562172 311646
rect 562308 311456 562428 311646
rect 562564 311456 562684 311646
rect 562820 311456 562940 311646
rect 563076 311456 563196 311646
rect 563332 311456 563452 311646
rect 563588 311456 563708 311646
rect 563844 311456 563964 311646
rect 564100 311456 564220 311646
rect 564356 311456 564476 311646
rect 564612 311456 564732 311646
rect 564868 311456 564988 311646
rect 565124 311456 565244 311646
rect 565380 311456 565500 311646
rect 575256 311470 575376 311716
rect 575512 311470 575632 311716
rect 575768 311470 575888 311716
rect 576024 311470 576144 311716
rect 576280 311470 576400 311716
rect 576536 311470 576656 311716
rect 576792 311470 576912 311716
rect 577048 311470 577168 311716
rect 577304 311470 577424 311716
rect 577560 311470 577680 311716
rect 577816 311470 577936 311716
rect 578072 311470 578192 311716
rect 578328 311470 578448 311716
rect 578584 311470 578704 311716
rect 578840 311470 578960 311716
rect 579096 311470 579216 311716
rect 579352 311470 579472 311716
rect 579608 311470 579728 311716
rect 579864 311470 579984 311716
rect 580120 311470 580240 311716
rect 560404 311436 565540 311456
rect 560404 311376 560590 311436
rect 560650 311376 560790 311436
rect 560850 311376 560990 311436
rect 561050 311376 561190 311436
rect 561250 311376 561390 311436
rect 561450 311376 561590 311436
rect 561650 311376 561790 311436
rect 561850 311376 561990 311436
rect 562050 311376 562190 311436
rect 562250 311376 562390 311436
rect 562450 311376 562590 311436
rect 562650 311376 562790 311436
rect 562850 311376 562990 311436
rect 563050 311376 563190 311436
rect 563250 311376 563390 311436
rect 563450 311376 563590 311436
rect 563650 311376 563790 311436
rect 563850 311376 563990 311436
rect 564050 311376 564190 311436
rect 564250 311376 564390 311436
rect 564450 311376 564590 311436
rect 564650 311376 564790 311436
rect 564850 311376 564990 311436
rect 565050 311376 565190 311436
rect 565250 311376 565390 311436
rect 565450 311376 565540 311436
rect 560404 311356 565540 311376
rect 575092 311450 580380 311470
rect 575092 311390 575150 311450
rect 575210 311390 575350 311450
rect 575410 311390 575550 311450
rect 575610 311390 575750 311450
rect 575810 311390 575950 311450
rect 576010 311390 576150 311450
rect 576210 311390 576350 311450
rect 576410 311390 576550 311450
rect 576610 311390 576750 311450
rect 576810 311390 576950 311450
rect 577010 311390 577150 311450
rect 577210 311390 577350 311450
rect 577410 311390 577550 311450
rect 577610 311390 577750 311450
rect 577810 311390 577950 311450
rect 578010 311390 578150 311450
rect 578210 311390 578350 311450
rect 578410 311390 578550 311450
rect 578610 311390 578750 311450
rect 578810 311390 578950 311450
rect 579010 311390 579150 311450
rect 579210 311390 579350 311450
rect 579410 311390 579550 311450
rect 579610 311390 579750 311450
rect 579810 311390 579950 311450
rect 580010 311390 580150 311450
rect 580210 311390 580380 311450
rect 575092 311370 580380 311390
<< polycont >>
rect 560836 492144 560896 492204
rect 561036 492144 561096 492204
rect 561236 492144 561296 492204
rect 561436 492144 561496 492204
rect 561636 492144 561696 492204
rect 561836 492144 561896 492204
rect 562036 492144 562096 492204
rect 562236 492144 562296 492204
rect 562436 492144 562496 492204
rect 562636 492144 562696 492204
rect 562836 492144 562896 492204
rect 563036 492144 563096 492204
rect 563236 492144 563296 492204
rect 563436 492144 563496 492204
rect 563636 492144 563696 492204
rect 563836 492144 563896 492204
rect 564036 492144 564096 492204
rect 564236 492144 564296 492204
rect 564436 492144 564496 492204
rect 564636 492144 564696 492204
rect 564836 492144 564896 492204
rect 565036 492144 565096 492204
rect 565236 492144 565296 492204
rect 565436 492144 565496 492204
rect 565636 492144 565696 492204
rect 575228 491862 575288 491922
rect 575428 491862 575488 491922
rect 575628 491862 575688 491922
rect 575828 491862 575888 491922
rect 576028 491862 576088 491922
rect 576228 491862 576288 491922
rect 576428 491862 576488 491922
rect 576628 491862 576688 491922
rect 576828 491862 576888 491922
rect 577028 491862 577088 491922
rect 577228 491862 577288 491922
rect 577428 491862 577488 491922
rect 577628 491862 577688 491922
rect 577828 491862 577888 491922
rect 578028 491862 578088 491922
rect 578228 491862 578288 491922
rect 578428 491862 578488 491922
rect 578628 491862 578688 491922
rect 578828 491862 578888 491922
rect 579028 491862 579088 491922
rect 579228 491862 579288 491922
rect 579428 491862 579488 491922
rect 579628 491862 579688 491922
rect 579828 491862 579888 491922
rect 580028 491862 580088 491922
rect 580228 491862 580288 491922
rect 560772 403002 560832 403062
rect 560972 403002 561032 403062
rect 561172 403002 561232 403062
rect 561372 403002 561432 403062
rect 561572 403002 561632 403062
rect 561772 403002 561832 403062
rect 561972 403002 562032 403062
rect 562172 403002 562232 403062
rect 562372 403002 562432 403062
rect 562572 403002 562632 403062
rect 562772 403002 562832 403062
rect 562972 403002 563032 403062
rect 563172 403002 563232 403062
rect 563372 403002 563432 403062
rect 563572 403002 563632 403062
rect 563772 403002 563832 403062
rect 563972 403002 564032 403062
rect 564172 403002 564232 403062
rect 564372 403002 564432 403062
rect 564572 403002 564632 403062
rect 564772 403002 564832 403062
rect 564972 403002 565032 403062
rect 565172 403002 565232 403062
rect 565372 403002 565432 403062
rect 565572 403002 565632 403062
rect 574506 402986 574566 403046
rect 574706 402986 574766 403046
rect 574906 402986 574966 403046
rect 575106 402986 575166 403046
rect 575306 402986 575366 403046
rect 575506 402986 575566 403046
rect 575706 402986 575766 403046
rect 575906 402986 575966 403046
rect 576106 402986 576166 403046
rect 576306 402986 576366 403046
rect 576506 402986 576566 403046
rect 576706 402986 576766 403046
rect 576906 402986 576966 403046
rect 577106 402986 577166 403046
rect 577306 402986 577366 403046
rect 577506 402986 577566 403046
rect 577706 402986 577766 403046
rect 577906 402986 577966 403046
rect 578106 402986 578166 403046
rect 578306 402986 578366 403046
rect 578506 402986 578566 403046
rect 578706 402986 578766 403046
rect 578906 402986 578966 403046
rect 579106 402986 579166 403046
rect 579306 402986 579366 403046
rect 579506 402986 579566 403046
rect 560728 357684 560788 357744
rect 560928 357684 560988 357744
rect 561128 357684 561188 357744
rect 561328 357684 561388 357744
rect 561528 357684 561588 357744
rect 561728 357684 561788 357744
rect 561928 357684 561988 357744
rect 562128 357684 562188 357744
rect 562328 357684 562388 357744
rect 562528 357684 562588 357744
rect 562728 357684 562788 357744
rect 562928 357684 562988 357744
rect 563128 357684 563188 357744
rect 563328 357684 563388 357744
rect 563528 357684 563588 357744
rect 563728 357684 563788 357744
rect 563928 357684 563988 357744
rect 564128 357684 564188 357744
rect 564328 357684 564388 357744
rect 564528 357684 564588 357744
rect 564728 357684 564788 357744
rect 564928 357684 564988 357744
rect 565128 357684 565188 357744
rect 565328 357684 565388 357744
rect 565528 357684 565588 357744
rect 574702 357558 574762 357618
rect 574902 357558 574962 357618
rect 575102 357558 575162 357618
rect 575302 357558 575362 357618
rect 575502 357558 575562 357618
rect 575702 357558 575762 357618
rect 575902 357558 575962 357618
rect 576102 357558 576162 357618
rect 576302 357558 576362 357618
rect 576502 357558 576562 357618
rect 576702 357558 576762 357618
rect 576902 357558 576962 357618
rect 577102 357558 577162 357618
rect 577302 357558 577362 357618
rect 577502 357558 577562 357618
rect 577702 357558 577762 357618
rect 577902 357558 577962 357618
rect 578102 357558 578162 357618
rect 578302 357558 578362 357618
rect 578502 357558 578562 357618
rect 578702 357558 578762 357618
rect 578902 357558 578962 357618
rect 579102 357558 579162 357618
rect 579302 357558 579362 357618
rect 579502 357558 579562 357618
rect 579702 357558 579762 357618
rect 560590 311376 560650 311436
rect 560790 311376 560850 311436
rect 560990 311376 561050 311436
rect 561190 311376 561250 311436
rect 561390 311376 561450 311436
rect 561590 311376 561650 311436
rect 561790 311376 561850 311436
rect 561990 311376 562050 311436
rect 562190 311376 562250 311436
rect 562390 311376 562450 311436
rect 562590 311376 562650 311436
rect 562790 311376 562850 311436
rect 562990 311376 563050 311436
rect 563190 311376 563250 311436
rect 563390 311376 563450 311436
rect 563590 311376 563650 311436
rect 563790 311376 563850 311436
rect 563990 311376 564050 311436
rect 564190 311376 564250 311436
rect 564390 311376 564450 311436
rect 564590 311376 564650 311436
rect 564790 311376 564850 311436
rect 564990 311376 565050 311436
rect 565190 311376 565250 311436
rect 565390 311376 565450 311436
rect 575150 311390 575210 311450
rect 575350 311390 575410 311450
rect 575550 311390 575610 311450
rect 575750 311390 575810 311450
rect 575950 311390 576010 311450
rect 576150 311390 576210 311450
rect 576350 311390 576410 311450
rect 576550 311390 576610 311450
rect 576750 311390 576810 311450
rect 576950 311390 577010 311450
rect 577150 311390 577210 311450
rect 577350 311390 577410 311450
rect 577550 311390 577610 311450
rect 577750 311390 577810 311450
rect 577950 311390 578010 311450
rect 578150 311390 578210 311450
rect 578350 311390 578410 311450
rect 578550 311390 578610 311450
rect 578750 311390 578810 311450
rect 578950 311390 579010 311450
rect 579150 311390 579210 311450
rect 579350 311390 579410 311450
rect 579550 311390 579610 311450
rect 579750 311390 579810 311450
rect 579950 311390 580010 311450
rect 580150 311390 580210 311450
<< locali >>
rect 560650 493790 560836 493850
rect 560896 493790 561036 493850
rect 561096 493790 561236 493850
rect 561296 493790 561436 493850
rect 561496 493790 561636 493850
rect 561696 493790 561836 493850
rect 561896 493790 562036 493850
rect 562096 493790 562236 493850
rect 562296 493790 562436 493850
rect 562496 493790 562636 493850
rect 562696 493790 562836 493850
rect 562896 493790 563036 493850
rect 563096 493790 563236 493850
rect 563296 493790 563436 493850
rect 563496 493790 563636 493850
rect 563696 493790 563836 493850
rect 563896 493790 564036 493850
rect 564096 493790 564236 493850
rect 564296 493790 564436 493850
rect 564496 493790 564636 493850
rect 564696 493790 564836 493850
rect 564896 493790 565036 493850
rect 565096 493790 565236 493850
rect 565296 493790 565436 493850
rect 565496 493790 565636 493850
rect 565696 493790 565964 493850
rect 560388 493690 560448 493692
rect 560388 493630 565866 493690
rect 560388 492522 560482 493630
rect 560342 492504 560482 492522
rect 560330 492482 560482 492504
rect 560330 492332 560340 492482
rect 560472 492332 560482 492482
rect 560661 493428 560695 493444
rect 560661 492436 560695 492452
rect 560919 493428 560953 493630
rect 560919 492436 560953 492452
rect 561177 493428 561211 493444
rect 561177 492370 561211 492452
rect 561435 493428 561469 493630
rect 561435 492436 561469 492452
rect 561693 493428 561727 493444
rect 561693 492370 561727 492452
rect 561951 493428 561985 493630
rect 561951 492436 561985 492452
rect 562209 493428 562243 493444
rect 562209 492370 562243 492452
rect 562467 493428 562501 493630
rect 562467 492436 562501 492452
rect 562725 493428 562759 493444
rect 562725 492370 562759 492452
rect 562983 493428 563017 493630
rect 562983 492436 563017 492452
rect 563241 493428 563275 493444
rect 563241 492370 563275 492452
rect 563499 493428 563533 493630
rect 563499 492436 563533 492452
rect 563757 493428 563791 493444
rect 563757 492370 563791 492452
rect 564015 493428 564049 493630
rect 564015 492436 564049 492452
rect 564273 493428 564307 493444
rect 564273 492370 564307 492452
rect 564531 493428 564565 493630
rect 564531 492436 564565 492452
rect 564789 493428 564823 493444
rect 564789 492370 564823 492452
rect 565047 493428 565081 493630
rect 565047 492436 565081 492452
rect 565305 493428 565339 493444
rect 565305 492370 565339 492452
rect 565563 493428 565597 493630
rect 575170 493564 575228 493624
rect 575288 493564 575428 493624
rect 575488 493564 575628 493624
rect 575688 493564 575828 493624
rect 575888 493564 576028 493624
rect 576088 493564 576228 493624
rect 576288 493564 576428 493624
rect 576488 493564 576628 493624
rect 576688 493564 576828 493624
rect 576888 493564 577028 493624
rect 577088 493564 577228 493624
rect 577288 493564 577428 493624
rect 577488 493564 577628 493624
rect 577688 493564 577828 493624
rect 577888 493564 578028 493624
rect 578088 493564 578228 493624
rect 578288 493564 578428 493624
rect 578488 493564 578628 493624
rect 578688 493564 578828 493624
rect 578888 493564 579028 493624
rect 579088 493564 579228 493624
rect 579288 493564 579428 493624
rect 579488 493564 579628 493624
rect 579688 493564 579828 493624
rect 579888 493564 580028 493624
rect 580088 493564 580228 493624
rect 580288 493564 580556 493624
rect 576720 493522 576880 493564
rect 576720 493486 576776 493522
rect 576820 493486 576880 493522
rect 576720 493484 576880 493486
rect 578020 493522 578180 493564
rect 578020 493486 578076 493522
rect 578120 493486 578180 493522
rect 578020 493484 578180 493486
rect 579320 493522 579480 493564
rect 579320 493486 579376 493522
rect 579420 493486 579480 493522
rect 579320 493484 579480 493486
rect 580468 493474 580528 493564
rect 574980 493444 575040 493446
rect 565563 492436 565597 492452
rect 565821 493428 565855 493444
rect 565821 492444 565855 492452
rect 574980 493404 580398 493444
rect 580468 493434 580478 493474
rect 580518 493434 580528 493474
rect 574980 493384 580396 493404
rect 565821 492424 565880 492444
rect 565821 492370 566074 492424
rect 560330 492312 560482 492332
rect 560388 492204 560482 492312
rect 560648 492320 566074 492370
rect 566234 492320 566240 492424
rect 560648 492310 566240 492320
rect 560388 492144 560836 492204
rect 560896 492144 561036 492204
rect 561096 492144 561236 492204
rect 561296 492144 561436 492204
rect 561496 492144 561636 492204
rect 561696 492144 561836 492204
rect 561896 492144 562036 492204
rect 562096 492144 562236 492204
rect 562296 492144 562436 492204
rect 562496 492144 562636 492204
rect 562696 492144 562836 492204
rect 562896 492144 563036 492204
rect 563096 492144 563236 492204
rect 563296 492144 563436 492204
rect 563496 492144 563636 492204
rect 563696 492144 563836 492204
rect 563896 492144 564036 492204
rect 564096 492144 564236 492204
rect 564296 492144 564436 492204
rect 564496 492144 564636 492204
rect 564696 492144 564836 492204
rect 564896 492144 565036 492204
rect 565096 492144 565236 492204
rect 565296 492144 565436 492204
rect 565496 492144 565636 492204
rect 565696 492144 565786 492204
rect 565876 492100 565936 492180
rect 562128 492068 562288 492090
rect 562128 492032 562184 492068
rect 562228 492032 562288 492068
rect 562128 491970 562288 492032
rect 563428 492068 563588 492090
rect 563428 492032 563484 492068
rect 563528 492032 563588 492068
rect 563428 491970 563588 492032
rect 564728 492068 564888 492090
rect 564728 492032 564784 492068
rect 564828 492032 564888 492068
rect 564728 491970 564888 492032
rect 565876 492060 565886 492100
rect 565926 492060 565936 492100
rect 565876 491970 565936 492060
rect 574980 492038 575040 493384
rect 575217 493202 575251 493218
rect 575217 492084 575251 492226
rect 575475 493202 575509 493384
rect 575475 492210 575509 492226
rect 575733 493202 575767 493218
rect 575733 492084 575767 492226
rect 575991 493202 576025 493384
rect 575991 492210 576025 492226
rect 576249 493202 576283 493218
rect 576249 492084 576283 492226
rect 576507 493202 576541 493384
rect 576507 492210 576541 492226
rect 576765 493202 576799 493218
rect 576765 492084 576799 492226
rect 577023 493202 577057 493384
rect 577023 492210 577057 492226
rect 577281 493202 577315 493218
rect 577281 492084 577315 492226
rect 577539 493202 577573 493384
rect 577539 492210 577573 492226
rect 577797 493202 577831 493218
rect 577797 492084 577831 492226
rect 578055 493202 578089 493384
rect 578055 492210 578089 492226
rect 578313 493202 578347 493218
rect 578313 492084 578347 492226
rect 578571 493202 578605 493384
rect 578571 492210 578605 492226
rect 578829 493202 578863 493218
rect 578829 492084 578863 492226
rect 579087 493202 579121 493384
rect 579087 492210 579121 492226
rect 579345 493202 579379 493218
rect 579345 492084 579379 492226
rect 579603 493202 579637 493384
rect 579603 492210 579637 492226
rect 579861 493202 579895 493218
rect 579861 492084 579895 492226
rect 580119 493202 580153 493384
rect 580468 493354 580528 493434
rect 580119 492210 580153 492226
rect 580377 493202 580411 493218
rect 580377 492208 580411 492226
rect 580414 492118 580642 492128
rect 580414 492084 580542 492118
rect 574924 491984 575040 492038
rect 575164 492030 580542 492084
rect 580632 492030 580642 492118
rect 575164 492024 580642 492030
rect 560650 491910 560836 491970
rect 560896 491910 561036 491970
rect 561096 491910 561236 491970
rect 561296 491910 561436 491970
rect 561496 491910 561636 491970
rect 561696 491910 561836 491970
rect 561896 491910 562036 491970
rect 562096 491910 562236 491970
rect 562296 491910 562436 491970
rect 562496 491910 562636 491970
rect 562696 491910 562836 491970
rect 562896 491910 563036 491970
rect 563096 491910 563236 491970
rect 563296 491910 563436 491970
rect 563496 491910 563636 491970
rect 563696 491910 563836 491970
rect 563896 491910 564036 491970
rect 564096 491910 564236 491970
rect 564296 491910 564436 491970
rect 564496 491910 564636 491970
rect 564696 491910 564836 491970
rect 564896 491910 565036 491970
rect 565096 491910 565236 491970
rect 565296 491910 565436 491970
rect 565496 491910 565636 491970
rect 565696 491910 565964 491970
rect 574924 491880 574934 491984
rect 575026 491922 575040 491984
rect 575026 491880 575228 491922
rect 574924 491864 575228 491880
rect 574962 491862 575228 491864
rect 575288 491862 575428 491922
rect 575488 491862 575628 491922
rect 575688 491862 575828 491922
rect 575888 491862 576028 491922
rect 576088 491862 576228 491922
rect 576288 491862 576428 491922
rect 576488 491862 576628 491922
rect 576688 491862 576828 491922
rect 576888 491862 577028 491922
rect 577088 491862 577228 491922
rect 577288 491862 577428 491922
rect 577488 491862 577628 491922
rect 577688 491862 577828 491922
rect 577888 491862 578028 491922
rect 578088 491862 578228 491922
rect 578288 491862 578428 491922
rect 578488 491862 578628 491922
rect 578688 491862 578828 491922
rect 578888 491862 579028 491922
rect 579088 491862 579228 491922
rect 579288 491862 579428 491922
rect 579488 491862 579628 491922
rect 579688 491862 579828 491922
rect 579888 491862 580028 491922
rect 580088 491862 580228 491922
rect 580288 491862 580458 491922
rect 575170 491684 575228 491744
rect 575288 491684 575428 491744
rect 575488 491684 575628 491744
rect 575688 491684 575828 491744
rect 575888 491684 576028 491744
rect 576088 491684 576228 491744
rect 576288 491684 576428 491744
rect 576488 491684 576628 491744
rect 576688 491684 576828 491744
rect 576888 491684 577028 491744
rect 577088 491684 577228 491744
rect 577288 491684 577428 491744
rect 577488 491684 577628 491744
rect 577688 491684 577828 491744
rect 577888 491684 578028 491744
rect 578088 491684 578228 491744
rect 578288 491684 578428 491744
rect 578488 491684 578628 491744
rect 578688 491684 578828 491744
rect 578888 491684 579028 491744
rect 579088 491684 579228 491744
rect 579288 491684 579428 491744
rect 579488 491684 579628 491744
rect 579688 491684 579828 491744
rect 579888 491684 580028 491744
rect 580088 491684 580228 491744
rect 580288 491684 580556 491744
rect 560586 404648 560772 404708
rect 560832 404648 560972 404708
rect 561032 404648 561172 404708
rect 561232 404648 561372 404708
rect 561432 404648 561572 404708
rect 561632 404648 561772 404708
rect 561832 404648 561972 404708
rect 562032 404648 562172 404708
rect 562232 404648 562372 404708
rect 562432 404648 562572 404708
rect 562632 404648 562772 404708
rect 562832 404648 562972 404708
rect 563032 404648 563172 404708
rect 563232 404648 563372 404708
rect 563432 404648 563572 404708
rect 563632 404648 563772 404708
rect 563832 404648 563972 404708
rect 564032 404648 564172 404708
rect 564232 404648 564372 404708
rect 564432 404648 564572 404708
rect 564632 404648 564772 404708
rect 564832 404648 564972 404708
rect 565032 404648 565172 404708
rect 565232 404648 565372 404708
rect 565432 404648 565572 404708
rect 565632 404648 565900 404708
rect 574448 404688 574506 404748
rect 574566 404688 574706 404748
rect 574766 404688 574906 404748
rect 574966 404688 575106 404748
rect 575166 404688 575306 404748
rect 575366 404688 575506 404748
rect 575566 404688 575706 404748
rect 575766 404688 575906 404748
rect 575966 404688 576106 404748
rect 576166 404688 576306 404748
rect 576366 404688 576506 404748
rect 576566 404688 576706 404748
rect 576766 404688 576906 404748
rect 576966 404688 577106 404748
rect 577166 404688 577306 404748
rect 577366 404688 577506 404748
rect 577566 404688 577706 404748
rect 577766 404688 577906 404748
rect 577966 404688 578106 404748
rect 578166 404688 578306 404748
rect 578366 404688 578506 404748
rect 578566 404688 578706 404748
rect 578766 404688 578906 404748
rect 578966 404688 579106 404748
rect 579166 404688 579306 404748
rect 579366 404688 579506 404748
rect 579566 404688 579834 404748
rect 575998 404646 576158 404688
rect 575998 404610 576054 404646
rect 576098 404610 576158 404646
rect 575998 404608 576158 404610
rect 577298 404646 577458 404688
rect 577298 404610 577354 404646
rect 577398 404610 577458 404646
rect 577298 404608 577458 404610
rect 578598 404646 578758 404688
rect 578598 404610 578654 404646
rect 578698 404610 578758 404646
rect 578598 404608 578758 404610
rect 579746 404598 579806 404688
rect 574258 404568 574318 404570
rect 560324 404548 560384 404550
rect 560324 404488 565802 404548
rect 574258 404528 579676 404568
rect 579746 404558 579756 404598
rect 579796 404558 579806 404598
rect 574258 404508 579674 404528
rect 560324 403380 560418 404488
rect 560278 403362 560418 403380
rect 560266 403340 560418 403362
rect 560266 403190 560276 403340
rect 560408 403190 560418 403340
rect 560597 404286 560631 404302
rect 560597 403294 560631 403310
rect 560855 404286 560889 404488
rect 560855 403294 560889 403310
rect 561113 404286 561147 404302
rect 561113 403228 561147 403310
rect 561371 404286 561405 404488
rect 561371 403294 561405 403310
rect 561629 404286 561663 404302
rect 561629 403228 561663 403310
rect 561887 404286 561921 404488
rect 561887 403294 561921 403310
rect 562145 404286 562179 404302
rect 562145 403228 562179 403310
rect 562403 404286 562437 404488
rect 562403 403294 562437 403310
rect 562661 404286 562695 404302
rect 562661 403228 562695 403310
rect 562919 404286 562953 404488
rect 562919 403294 562953 403310
rect 563177 404286 563211 404302
rect 563177 403228 563211 403310
rect 563435 404286 563469 404488
rect 563435 403294 563469 403310
rect 563693 404286 563727 404302
rect 563693 403228 563727 403310
rect 563951 404286 563985 404488
rect 563951 403294 563985 403310
rect 564209 404286 564243 404302
rect 564209 403228 564243 403310
rect 564467 404286 564501 404488
rect 564467 403294 564501 403310
rect 564725 404286 564759 404302
rect 564725 403228 564759 403310
rect 564983 404286 565017 404488
rect 564983 403294 565017 403310
rect 565241 404286 565275 404302
rect 565241 403228 565275 403310
rect 565499 404286 565533 404488
rect 565499 403294 565533 403310
rect 565757 404286 565791 404302
rect 565757 403302 565791 403310
rect 565757 403282 565816 403302
rect 565757 403228 566010 403282
rect 560266 403170 560418 403190
rect 560324 403062 560418 403170
rect 560584 403178 566010 403228
rect 566170 403178 566176 403282
rect 560584 403168 566176 403178
rect 574258 403162 574318 404508
rect 574495 404326 574529 404342
rect 574495 403208 574529 403350
rect 574753 404326 574787 404508
rect 574753 403334 574787 403350
rect 575011 404326 575045 404342
rect 575011 403208 575045 403350
rect 575269 404326 575303 404508
rect 575269 403334 575303 403350
rect 575527 404326 575561 404342
rect 575527 403208 575561 403350
rect 575785 404326 575819 404508
rect 575785 403334 575819 403350
rect 576043 404326 576077 404342
rect 576043 403208 576077 403350
rect 576301 404326 576335 404508
rect 576301 403334 576335 403350
rect 576559 404326 576593 404342
rect 576559 403208 576593 403350
rect 576817 404326 576851 404508
rect 576817 403334 576851 403350
rect 577075 404326 577109 404342
rect 577075 403208 577109 403350
rect 577333 404326 577367 404508
rect 577333 403334 577367 403350
rect 577591 404326 577625 404342
rect 577591 403208 577625 403350
rect 577849 404326 577883 404508
rect 577849 403334 577883 403350
rect 578107 404326 578141 404342
rect 578107 403208 578141 403350
rect 578365 404326 578399 404508
rect 578365 403334 578399 403350
rect 578623 404326 578657 404342
rect 578623 403208 578657 403350
rect 578881 404326 578915 404508
rect 578881 403334 578915 403350
rect 579139 404326 579173 404342
rect 579139 403208 579173 403350
rect 579397 404326 579431 404508
rect 579746 404478 579806 404558
rect 579397 403334 579431 403350
rect 579655 404326 579689 404342
rect 579655 403332 579689 403350
rect 579692 403242 579920 403252
rect 579692 403208 579820 403242
rect 574202 403108 574318 403162
rect 574442 403154 579820 403208
rect 579910 403154 579920 403242
rect 574442 403148 579920 403154
rect 560324 403002 560772 403062
rect 560832 403002 560972 403062
rect 561032 403002 561172 403062
rect 561232 403002 561372 403062
rect 561432 403002 561572 403062
rect 561632 403002 561772 403062
rect 561832 403002 561972 403062
rect 562032 403002 562172 403062
rect 562232 403002 562372 403062
rect 562432 403002 562572 403062
rect 562632 403002 562772 403062
rect 562832 403002 562972 403062
rect 563032 403002 563172 403062
rect 563232 403002 563372 403062
rect 563432 403002 563572 403062
rect 563632 403002 563772 403062
rect 563832 403002 563972 403062
rect 564032 403002 564172 403062
rect 564232 403002 564372 403062
rect 564432 403002 564572 403062
rect 564632 403002 564772 403062
rect 564832 403002 564972 403062
rect 565032 403002 565172 403062
rect 565232 403002 565372 403062
rect 565432 403002 565572 403062
rect 565632 403002 565722 403062
rect 565812 402958 565872 403038
rect 574202 403004 574212 403108
rect 574304 403046 574318 403108
rect 574304 403004 574506 403046
rect 574202 402988 574506 403004
rect 574240 402986 574506 402988
rect 574566 402986 574706 403046
rect 574766 402986 574906 403046
rect 574966 402986 575106 403046
rect 575166 402986 575306 403046
rect 575366 402986 575506 403046
rect 575566 402986 575706 403046
rect 575766 402986 575906 403046
rect 575966 402986 576106 403046
rect 576166 402986 576306 403046
rect 576366 402986 576506 403046
rect 576566 402986 576706 403046
rect 576766 402986 576906 403046
rect 576966 402986 577106 403046
rect 577166 402986 577306 403046
rect 577366 402986 577506 403046
rect 577566 402986 577706 403046
rect 577766 402986 577906 403046
rect 577966 402986 578106 403046
rect 578166 402986 578306 403046
rect 578366 402986 578506 403046
rect 578566 402986 578706 403046
rect 578766 402986 578906 403046
rect 578966 402986 579106 403046
rect 579166 402986 579306 403046
rect 579366 402986 579506 403046
rect 579566 402986 579736 403046
rect 562064 402926 562224 402948
rect 562064 402890 562120 402926
rect 562164 402890 562224 402926
rect 562064 402828 562224 402890
rect 563364 402926 563524 402948
rect 563364 402890 563420 402926
rect 563464 402890 563524 402926
rect 563364 402828 563524 402890
rect 564664 402926 564824 402948
rect 564664 402890 564720 402926
rect 564764 402890 564824 402926
rect 564664 402828 564824 402890
rect 565812 402918 565822 402958
rect 565862 402918 565872 402958
rect 565812 402828 565872 402918
rect 560586 402768 560772 402828
rect 560832 402768 560972 402828
rect 561032 402768 561172 402828
rect 561232 402768 561372 402828
rect 561432 402768 561572 402828
rect 561632 402768 561772 402828
rect 561832 402768 561972 402828
rect 562032 402768 562172 402828
rect 562232 402768 562372 402828
rect 562432 402768 562572 402828
rect 562632 402768 562772 402828
rect 562832 402768 562972 402828
rect 563032 402768 563172 402828
rect 563232 402768 563372 402828
rect 563432 402768 563572 402828
rect 563632 402768 563772 402828
rect 563832 402768 563972 402828
rect 564032 402768 564172 402828
rect 564232 402768 564372 402828
rect 564432 402768 564572 402828
rect 564632 402768 564772 402828
rect 564832 402768 564972 402828
rect 565032 402768 565172 402828
rect 565232 402768 565372 402828
rect 565432 402768 565572 402828
rect 565632 402768 565900 402828
rect 574448 402808 574506 402868
rect 574566 402808 574706 402868
rect 574766 402808 574906 402868
rect 574966 402808 575106 402868
rect 575166 402808 575306 402868
rect 575366 402808 575506 402868
rect 575566 402808 575706 402868
rect 575766 402808 575906 402868
rect 575966 402808 576106 402868
rect 576166 402808 576306 402868
rect 576366 402808 576506 402868
rect 576566 402808 576706 402868
rect 576766 402808 576906 402868
rect 576966 402808 577106 402868
rect 577166 402808 577306 402868
rect 577366 402808 577506 402868
rect 577566 402808 577706 402868
rect 577766 402808 577906 402868
rect 577966 402808 578106 402868
rect 578166 402808 578306 402868
rect 578366 402808 578506 402868
rect 578566 402808 578706 402868
rect 578766 402808 578906 402868
rect 578966 402808 579106 402868
rect 579166 402808 579306 402868
rect 579366 402808 579506 402868
rect 579566 402808 579834 402868
rect 560542 359330 560728 359390
rect 560788 359330 560928 359390
rect 560988 359330 561128 359390
rect 561188 359330 561328 359390
rect 561388 359330 561528 359390
rect 561588 359330 561728 359390
rect 561788 359330 561928 359390
rect 561988 359330 562128 359390
rect 562188 359330 562328 359390
rect 562388 359330 562528 359390
rect 562588 359330 562728 359390
rect 562788 359330 562928 359390
rect 562988 359330 563128 359390
rect 563188 359330 563328 359390
rect 563388 359330 563528 359390
rect 563588 359330 563728 359390
rect 563788 359330 563928 359390
rect 563988 359330 564128 359390
rect 564188 359330 564328 359390
rect 564388 359330 564528 359390
rect 564588 359330 564728 359390
rect 564788 359330 564928 359390
rect 564988 359330 565128 359390
rect 565188 359330 565328 359390
rect 565388 359330 565528 359390
rect 565588 359330 565856 359390
rect 574644 359260 574702 359320
rect 574762 359260 574902 359320
rect 574962 359260 575102 359320
rect 575162 359260 575302 359320
rect 575362 359260 575502 359320
rect 575562 359260 575702 359320
rect 575762 359260 575902 359320
rect 575962 359260 576102 359320
rect 576162 359260 576302 359320
rect 576362 359260 576502 359320
rect 576562 359260 576702 359320
rect 576762 359260 576902 359320
rect 576962 359260 577102 359320
rect 577162 359260 577302 359320
rect 577362 359260 577502 359320
rect 577562 359260 577702 359320
rect 577762 359260 577902 359320
rect 577962 359260 578102 359320
rect 578162 359260 578302 359320
rect 578362 359260 578502 359320
rect 578562 359260 578702 359320
rect 578762 359260 578902 359320
rect 578962 359260 579102 359320
rect 579162 359260 579302 359320
rect 579362 359260 579502 359320
rect 579562 359260 579702 359320
rect 579762 359260 580030 359320
rect 560280 359230 560340 359232
rect 560280 359170 565758 359230
rect 576194 359218 576354 359260
rect 576194 359182 576250 359218
rect 576294 359182 576354 359218
rect 576194 359180 576354 359182
rect 577494 359218 577654 359260
rect 577494 359182 577550 359218
rect 577594 359182 577654 359218
rect 577494 359180 577654 359182
rect 578794 359218 578954 359260
rect 578794 359182 578850 359218
rect 578894 359182 578954 359218
rect 578794 359180 578954 359182
rect 579942 359170 580002 359260
rect 560280 358062 560374 359170
rect 560234 358044 560374 358062
rect 560222 358022 560374 358044
rect 560222 357872 560232 358022
rect 560364 357872 560374 358022
rect 560553 358968 560587 358984
rect 560553 357976 560587 357992
rect 560811 358968 560845 359170
rect 560811 357976 560845 357992
rect 561069 358968 561103 358984
rect 561069 357910 561103 357992
rect 561327 358968 561361 359170
rect 561327 357976 561361 357992
rect 561585 358968 561619 358984
rect 561585 357910 561619 357992
rect 561843 358968 561877 359170
rect 561843 357976 561877 357992
rect 562101 358968 562135 358984
rect 562101 357910 562135 357992
rect 562359 358968 562393 359170
rect 562359 357976 562393 357992
rect 562617 358968 562651 358984
rect 562617 357910 562651 357992
rect 562875 358968 562909 359170
rect 562875 357976 562909 357992
rect 563133 358968 563167 358984
rect 563133 357910 563167 357992
rect 563391 358968 563425 359170
rect 563391 357976 563425 357992
rect 563649 358968 563683 358984
rect 563649 357910 563683 357992
rect 563907 358968 563941 359170
rect 563907 357976 563941 357992
rect 564165 358968 564199 358984
rect 564165 357910 564199 357992
rect 564423 358968 564457 359170
rect 564423 357976 564457 357992
rect 564681 358968 564715 358984
rect 564681 357910 564715 357992
rect 564939 358968 564973 359170
rect 564939 357976 564973 357992
rect 565197 358968 565231 358984
rect 565197 357910 565231 357992
rect 565455 358968 565489 359170
rect 574454 359140 574514 359142
rect 574454 359100 579872 359140
rect 579942 359130 579952 359170
rect 579992 359130 580002 359170
rect 574454 359080 579870 359100
rect 565455 357976 565489 357992
rect 565713 358968 565747 358984
rect 565713 357984 565747 357992
rect 565713 357964 565772 357984
rect 565713 357910 565966 357964
rect 560222 357852 560374 357872
rect 560280 357744 560374 357852
rect 560540 357860 565966 357910
rect 566126 357860 566132 357964
rect 560540 357850 566132 357860
rect 560280 357684 560728 357744
rect 560788 357684 560928 357744
rect 560988 357684 561128 357744
rect 561188 357684 561328 357744
rect 561388 357684 561528 357744
rect 561588 357684 561728 357744
rect 561788 357684 561928 357744
rect 561988 357684 562128 357744
rect 562188 357684 562328 357744
rect 562388 357684 562528 357744
rect 562588 357684 562728 357744
rect 562788 357684 562928 357744
rect 562988 357684 563128 357744
rect 563188 357684 563328 357744
rect 563388 357684 563528 357744
rect 563588 357684 563728 357744
rect 563788 357684 563928 357744
rect 563988 357684 564128 357744
rect 564188 357684 564328 357744
rect 564388 357684 564528 357744
rect 564588 357684 564728 357744
rect 564788 357684 564928 357744
rect 564988 357684 565128 357744
rect 565188 357684 565328 357744
rect 565388 357684 565528 357744
rect 565588 357684 565678 357744
rect 574454 357734 574514 359080
rect 574691 358898 574725 358914
rect 574691 357780 574725 357922
rect 574949 358898 574983 359080
rect 574949 357906 574983 357922
rect 575207 358898 575241 358914
rect 575207 357780 575241 357922
rect 575465 358898 575499 359080
rect 575465 357906 575499 357922
rect 575723 358898 575757 358914
rect 575723 357780 575757 357922
rect 575981 358898 576015 359080
rect 575981 357906 576015 357922
rect 576239 358898 576273 358914
rect 576239 357780 576273 357922
rect 576497 358898 576531 359080
rect 576497 357906 576531 357922
rect 576755 358898 576789 358914
rect 576755 357780 576789 357922
rect 577013 358898 577047 359080
rect 577013 357906 577047 357922
rect 577271 358898 577305 358914
rect 577271 357780 577305 357922
rect 577529 358898 577563 359080
rect 577529 357906 577563 357922
rect 577787 358898 577821 358914
rect 577787 357780 577821 357922
rect 578045 358898 578079 359080
rect 578045 357906 578079 357922
rect 578303 358898 578337 358914
rect 578303 357780 578337 357922
rect 578561 358898 578595 359080
rect 578561 357906 578595 357922
rect 578819 358898 578853 358914
rect 578819 357780 578853 357922
rect 579077 358898 579111 359080
rect 579077 357906 579111 357922
rect 579335 358898 579369 358914
rect 579335 357780 579369 357922
rect 579593 358898 579627 359080
rect 579942 359050 580002 359130
rect 579593 357906 579627 357922
rect 579851 358898 579885 358914
rect 579851 357904 579885 357922
rect 579888 357814 580116 357824
rect 579888 357780 580016 357814
rect 565768 357640 565828 357720
rect 562020 357608 562180 357630
rect 562020 357572 562076 357608
rect 562120 357572 562180 357608
rect 562020 357510 562180 357572
rect 563320 357608 563480 357630
rect 563320 357572 563376 357608
rect 563420 357572 563480 357608
rect 563320 357510 563480 357572
rect 564620 357608 564780 357630
rect 564620 357572 564676 357608
rect 564720 357572 564780 357608
rect 564620 357510 564780 357572
rect 565768 357600 565778 357640
rect 565818 357600 565828 357640
rect 565768 357510 565828 357600
rect 574398 357680 574514 357734
rect 574638 357726 580016 357780
rect 580106 357726 580116 357814
rect 574638 357720 580116 357726
rect 574398 357576 574408 357680
rect 574500 357618 574514 357680
rect 574500 357576 574702 357618
rect 574398 357560 574702 357576
rect 574436 357558 574702 357560
rect 574762 357558 574902 357618
rect 574962 357558 575102 357618
rect 575162 357558 575302 357618
rect 575362 357558 575502 357618
rect 575562 357558 575702 357618
rect 575762 357558 575902 357618
rect 575962 357558 576102 357618
rect 576162 357558 576302 357618
rect 576362 357558 576502 357618
rect 576562 357558 576702 357618
rect 576762 357558 576902 357618
rect 576962 357558 577102 357618
rect 577162 357558 577302 357618
rect 577362 357558 577502 357618
rect 577562 357558 577702 357618
rect 577762 357558 577902 357618
rect 577962 357558 578102 357618
rect 578162 357558 578302 357618
rect 578362 357558 578502 357618
rect 578562 357558 578702 357618
rect 578762 357558 578902 357618
rect 578962 357558 579102 357618
rect 579162 357558 579302 357618
rect 579362 357558 579502 357618
rect 579562 357558 579702 357618
rect 579762 357558 579932 357618
rect 560542 357450 560728 357510
rect 560788 357450 560928 357510
rect 560988 357450 561128 357510
rect 561188 357450 561328 357510
rect 561388 357450 561528 357510
rect 561588 357450 561728 357510
rect 561788 357450 561928 357510
rect 561988 357450 562128 357510
rect 562188 357450 562328 357510
rect 562388 357450 562528 357510
rect 562588 357450 562728 357510
rect 562788 357450 562928 357510
rect 562988 357450 563128 357510
rect 563188 357450 563328 357510
rect 563388 357450 563528 357510
rect 563588 357450 563728 357510
rect 563788 357450 563928 357510
rect 563988 357450 564128 357510
rect 564188 357450 564328 357510
rect 564388 357450 564528 357510
rect 564588 357450 564728 357510
rect 564788 357450 564928 357510
rect 564988 357450 565128 357510
rect 565188 357450 565328 357510
rect 565388 357450 565528 357510
rect 565588 357450 565856 357510
rect 574644 357380 574702 357440
rect 574762 357380 574902 357440
rect 574962 357380 575102 357440
rect 575162 357380 575302 357440
rect 575362 357380 575502 357440
rect 575562 357380 575702 357440
rect 575762 357380 575902 357440
rect 575962 357380 576102 357440
rect 576162 357380 576302 357440
rect 576362 357380 576502 357440
rect 576562 357380 576702 357440
rect 576762 357380 576902 357440
rect 576962 357380 577102 357440
rect 577162 357380 577302 357440
rect 577362 357380 577502 357440
rect 577562 357380 577702 357440
rect 577762 357380 577902 357440
rect 577962 357380 578102 357440
rect 578162 357380 578302 357440
rect 578362 357380 578502 357440
rect 578562 357380 578702 357440
rect 578762 357380 578902 357440
rect 578962 357380 579102 357440
rect 579162 357380 579302 357440
rect 579362 357380 579502 357440
rect 579562 357380 579702 357440
rect 579762 357380 580030 357440
rect 575092 313092 575150 313152
rect 575210 313092 575350 313152
rect 575410 313092 575550 313152
rect 575610 313092 575750 313152
rect 575810 313092 575950 313152
rect 576010 313092 576150 313152
rect 576210 313092 576350 313152
rect 576410 313092 576550 313152
rect 576610 313092 576750 313152
rect 576810 313092 576950 313152
rect 577010 313092 577150 313152
rect 577210 313092 577350 313152
rect 577410 313092 577550 313152
rect 577610 313092 577750 313152
rect 577810 313092 577950 313152
rect 578010 313092 578150 313152
rect 578210 313092 578350 313152
rect 578410 313092 578550 313152
rect 578610 313092 578750 313152
rect 578810 313092 578950 313152
rect 579010 313092 579150 313152
rect 579210 313092 579350 313152
rect 579410 313092 579550 313152
rect 579610 313092 579750 313152
rect 579810 313092 579950 313152
rect 580010 313092 580150 313152
rect 580210 313092 580478 313152
rect 560404 313022 560590 313082
rect 560650 313022 560790 313082
rect 560850 313022 560990 313082
rect 561050 313022 561190 313082
rect 561250 313022 561390 313082
rect 561450 313022 561590 313082
rect 561650 313022 561790 313082
rect 561850 313022 561990 313082
rect 562050 313022 562190 313082
rect 562250 313022 562390 313082
rect 562450 313022 562590 313082
rect 562650 313022 562790 313082
rect 562850 313022 562990 313082
rect 563050 313022 563190 313082
rect 563250 313022 563390 313082
rect 563450 313022 563590 313082
rect 563650 313022 563790 313082
rect 563850 313022 563990 313082
rect 564050 313022 564190 313082
rect 564250 313022 564390 313082
rect 564450 313022 564590 313082
rect 564650 313022 564790 313082
rect 564850 313022 564990 313082
rect 565050 313022 565190 313082
rect 565250 313022 565390 313082
rect 565450 313022 565718 313082
rect 576642 313050 576802 313092
rect 576642 313014 576698 313050
rect 576742 313014 576802 313050
rect 576642 313012 576802 313014
rect 577942 313050 578102 313092
rect 577942 313014 577998 313050
rect 578042 313014 578102 313050
rect 577942 313012 578102 313014
rect 579242 313050 579402 313092
rect 579242 313014 579298 313050
rect 579342 313014 579402 313050
rect 579242 313012 579402 313014
rect 580390 313002 580450 313092
rect 574902 312972 574962 312974
rect 574902 312932 580320 312972
rect 580390 312962 580400 313002
rect 580440 312962 580450 313002
rect 560142 312922 560202 312924
rect 560142 312862 565620 312922
rect 574902 312912 580318 312932
rect 560142 311754 560236 312862
rect 560096 311736 560236 311754
rect 560084 311714 560236 311736
rect 560084 311564 560094 311714
rect 560226 311564 560236 311714
rect 560415 312660 560449 312676
rect 560415 311668 560449 311684
rect 560673 312660 560707 312862
rect 560673 311668 560707 311684
rect 560931 312660 560965 312676
rect 560931 311602 560965 311684
rect 561189 312660 561223 312862
rect 561189 311668 561223 311684
rect 561447 312660 561481 312676
rect 561447 311602 561481 311684
rect 561705 312660 561739 312862
rect 561705 311668 561739 311684
rect 561963 312660 561997 312676
rect 561963 311602 561997 311684
rect 562221 312660 562255 312862
rect 562221 311668 562255 311684
rect 562479 312660 562513 312676
rect 562479 311602 562513 311684
rect 562737 312660 562771 312862
rect 562737 311668 562771 311684
rect 562995 312660 563029 312676
rect 562995 311602 563029 311684
rect 563253 312660 563287 312862
rect 563253 311668 563287 311684
rect 563511 312660 563545 312676
rect 563511 311602 563545 311684
rect 563769 312660 563803 312862
rect 563769 311668 563803 311684
rect 564027 312660 564061 312676
rect 564027 311602 564061 311684
rect 564285 312660 564319 312862
rect 564285 311668 564319 311684
rect 564543 312660 564577 312676
rect 564543 311602 564577 311684
rect 564801 312660 564835 312862
rect 564801 311668 564835 311684
rect 565059 312660 565093 312676
rect 565059 311602 565093 311684
rect 565317 312660 565351 312862
rect 565317 311668 565351 311684
rect 565575 312660 565609 312676
rect 565575 311676 565609 311684
rect 565575 311656 565634 311676
rect 565575 311602 565828 311656
rect 560084 311544 560236 311564
rect 560142 311436 560236 311544
rect 560402 311552 565828 311602
rect 565988 311552 565994 311656
rect 574902 311566 574962 312912
rect 575139 312730 575173 312746
rect 575139 311612 575173 311754
rect 575397 312730 575431 312912
rect 575397 311738 575431 311754
rect 575655 312730 575689 312746
rect 575655 311612 575689 311754
rect 575913 312730 575947 312912
rect 575913 311738 575947 311754
rect 576171 312730 576205 312746
rect 576171 311612 576205 311754
rect 576429 312730 576463 312912
rect 576429 311738 576463 311754
rect 576687 312730 576721 312746
rect 576687 311612 576721 311754
rect 576945 312730 576979 312912
rect 576945 311738 576979 311754
rect 577203 312730 577237 312746
rect 577203 311612 577237 311754
rect 577461 312730 577495 312912
rect 577461 311738 577495 311754
rect 577719 312730 577753 312746
rect 577719 311612 577753 311754
rect 577977 312730 578011 312912
rect 577977 311738 578011 311754
rect 578235 312730 578269 312746
rect 578235 311612 578269 311754
rect 578493 312730 578527 312912
rect 578493 311738 578527 311754
rect 578751 312730 578785 312746
rect 578751 311612 578785 311754
rect 579009 312730 579043 312912
rect 579009 311738 579043 311754
rect 579267 312730 579301 312746
rect 579267 311612 579301 311754
rect 579525 312730 579559 312912
rect 579525 311738 579559 311754
rect 579783 312730 579817 312746
rect 579783 311612 579817 311754
rect 580041 312730 580075 312912
rect 580390 312882 580450 312962
rect 580041 311738 580075 311754
rect 580299 312730 580333 312746
rect 580299 311736 580333 311754
rect 580336 311646 580564 311656
rect 580336 311612 580464 311646
rect 560402 311542 565994 311552
rect 574846 311512 574962 311566
rect 575086 311558 580464 311612
rect 580554 311558 580564 311646
rect 575086 311552 580564 311558
rect 560142 311376 560590 311436
rect 560650 311376 560790 311436
rect 560850 311376 560990 311436
rect 561050 311376 561190 311436
rect 561250 311376 561390 311436
rect 561450 311376 561590 311436
rect 561650 311376 561790 311436
rect 561850 311376 561990 311436
rect 562050 311376 562190 311436
rect 562250 311376 562390 311436
rect 562450 311376 562590 311436
rect 562650 311376 562790 311436
rect 562850 311376 562990 311436
rect 563050 311376 563190 311436
rect 563250 311376 563390 311436
rect 563450 311376 563590 311436
rect 563650 311376 563790 311436
rect 563850 311376 563990 311436
rect 564050 311376 564190 311436
rect 564250 311376 564390 311436
rect 564450 311376 564590 311436
rect 564650 311376 564790 311436
rect 564850 311376 564990 311436
rect 565050 311376 565190 311436
rect 565250 311376 565390 311436
rect 565450 311376 565540 311436
rect 565630 311332 565690 311412
rect 574846 311408 574856 311512
rect 574948 311450 574962 311512
rect 574948 311408 575150 311450
rect 574846 311392 575150 311408
rect 574884 311390 575150 311392
rect 575210 311390 575350 311450
rect 575410 311390 575550 311450
rect 575610 311390 575750 311450
rect 575810 311390 575950 311450
rect 576010 311390 576150 311450
rect 576210 311390 576350 311450
rect 576410 311390 576550 311450
rect 576610 311390 576750 311450
rect 576810 311390 576950 311450
rect 577010 311390 577150 311450
rect 577210 311390 577350 311450
rect 577410 311390 577550 311450
rect 577610 311390 577750 311450
rect 577810 311390 577950 311450
rect 578010 311390 578150 311450
rect 578210 311390 578350 311450
rect 578410 311390 578550 311450
rect 578610 311390 578750 311450
rect 578810 311390 578950 311450
rect 579010 311390 579150 311450
rect 579210 311390 579350 311450
rect 579410 311390 579550 311450
rect 579610 311390 579750 311450
rect 579810 311390 579950 311450
rect 580010 311390 580150 311450
rect 580210 311390 580380 311450
rect 561882 311300 562042 311322
rect 561882 311264 561938 311300
rect 561982 311264 562042 311300
rect 561882 311202 562042 311264
rect 563182 311300 563342 311322
rect 563182 311264 563238 311300
rect 563282 311264 563342 311300
rect 563182 311202 563342 311264
rect 564482 311300 564642 311322
rect 564482 311264 564538 311300
rect 564582 311264 564642 311300
rect 564482 311202 564642 311264
rect 565630 311292 565640 311332
rect 565680 311292 565690 311332
rect 565630 311202 565690 311292
rect 575092 311212 575150 311272
rect 575210 311212 575350 311272
rect 575410 311212 575550 311272
rect 575610 311212 575750 311272
rect 575810 311212 575950 311272
rect 576010 311212 576150 311272
rect 576210 311212 576350 311272
rect 576410 311212 576550 311272
rect 576610 311212 576750 311272
rect 576810 311212 576950 311272
rect 577010 311212 577150 311272
rect 577210 311212 577350 311272
rect 577410 311212 577550 311272
rect 577610 311212 577750 311272
rect 577810 311212 577950 311272
rect 578010 311212 578150 311272
rect 578210 311212 578350 311272
rect 578410 311212 578550 311272
rect 578610 311212 578750 311272
rect 578810 311212 578950 311272
rect 579010 311212 579150 311272
rect 579210 311212 579350 311272
rect 579410 311212 579550 311272
rect 579610 311212 579750 311272
rect 579810 311212 579950 311272
rect 580010 311212 580150 311272
rect 580210 311212 580478 311272
rect 560404 311142 560590 311202
rect 560650 311142 560790 311202
rect 560850 311142 560990 311202
rect 561050 311142 561190 311202
rect 561250 311142 561390 311202
rect 561450 311142 561590 311202
rect 561650 311142 561790 311202
rect 561850 311142 561990 311202
rect 562050 311142 562190 311202
rect 562250 311142 562390 311202
rect 562450 311142 562590 311202
rect 562650 311142 562790 311202
rect 562850 311142 562990 311202
rect 563050 311142 563190 311202
rect 563250 311142 563390 311202
rect 563450 311142 563590 311202
rect 563650 311142 563790 311202
rect 563850 311142 563990 311202
rect 564050 311142 564190 311202
rect 564250 311142 564390 311202
rect 564450 311142 564590 311202
rect 564650 311142 564790 311202
rect 564850 311142 564990 311202
rect 565050 311142 565190 311202
rect 565250 311142 565390 311202
rect 565450 311142 565718 311202
<< viali >>
rect 560836 493790 560896 493850
rect 561036 493790 561096 493850
rect 561236 493790 561296 493850
rect 561436 493790 561496 493850
rect 561636 493790 561696 493850
rect 561836 493790 561896 493850
rect 562036 493790 562096 493850
rect 562236 493790 562296 493850
rect 562436 493790 562496 493850
rect 562636 493790 562696 493850
rect 562836 493790 562896 493850
rect 563036 493790 563096 493850
rect 563236 493790 563296 493850
rect 563436 493790 563496 493850
rect 563636 493790 563696 493850
rect 563836 493790 563896 493850
rect 564036 493790 564096 493850
rect 564236 493790 564296 493850
rect 564436 493790 564496 493850
rect 564636 493790 564696 493850
rect 564836 493790 564896 493850
rect 565036 493790 565096 493850
rect 565236 493790 565296 493850
rect 565436 493790 565496 493850
rect 565636 493790 565696 493850
rect 560340 492332 560472 492482
rect 560661 492452 560695 493428
rect 560919 492452 560953 493428
rect 561177 492452 561211 493428
rect 561435 492452 561469 493428
rect 561693 492452 561727 493428
rect 561951 492452 561985 493428
rect 562209 492452 562243 493428
rect 562467 492452 562501 493428
rect 562725 492452 562759 493428
rect 562983 492452 563017 493428
rect 563241 492452 563275 493428
rect 563499 492452 563533 493428
rect 563757 492452 563791 493428
rect 564015 492452 564049 493428
rect 564273 492452 564307 493428
rect 564531 492452 564565 493428
rect 564789 492452 564823 493428
rect 565047 492452 565081 493428
rect 565305 492452 565339 493428
rect 575228 493564 575288 493624
rect 575428 493564 575488 493624
rect 575628 493564 575688 493624
rect 575828 493564 575888 493624
rect 576028 493564 576088 493624
rect 576228 493564 576288 493624
rect 576428 493564 576488 493624
rect 576628 493564 576688 493624
rect 576828 493564 576888 493624
rect 577028 493564 577088 493624
rect 577228 493564 577288 493624
rect 577428 493564 577488 493624
rect 577628 493564 577688 493624
rect 577828 493564 577888 493624
rect 578028 493564 578088 493624
rect 578228 493564 578288 493624
rect 578428 493564 578488 493624
rect 578628 493564 578688 493624
rect 578828 493564 578888 493624
rect 579028 493564 579088 493624
rect 579228 493564 579288 493624
rect 579428 493564 579488 493624
rect 579628 493564 579688 493624
rect 579828 493564 579888 493624
rect 580028 493564 580088 493624
rect 580228 493564 580288 493624
rect 565563 492452 565597 493428
rect 565821 492452 565855 493428
rect 566074 492320 566234 492428
rect 575217 492226 575251 493202
rect 575475 492226 575509 493202
rect 575733 492226 575767 493202
rect 575991 492226 576025 493202
rect 576249 492226 576283 493202
rect 576507 492226 576541 493202
rect 576765 492226 576799 493202
rect 577023 492226 577057 493202
rect 577281 492226 577315 493202
rect 577539 492226 577573 493202
rect 577797 492226 577831 493202
rect 578055 492226 578089 493202
rect 578313 492226 578347 493202
rect 578571 492226 578605 493202
rect 578829 492226 578863 493202
rect 579087 492226 579121 493202
rect 579345 492226 579379 493202
rect 579603 492226 579637 493202
rect 579861 492226 579895 493202
rect 580119 492226 580153 493202
rect 580377 492226 580411 493202
rect 580542 492030 580632 492118
rect 560836 491910 560896 491970
rect 561036 491910 561096 491970
rect 561236 491910 561296 491970
rect 561436 491910 561496 491970
rect 561636 491910 561696 491970
rect 561836 491910 561896 491970
rect 562036 491910 562096 491970
rect 562236 491910 562296 491970
rect 562436 491910 562496 491970
rect 562636 491910 562696 491970
rect 562836 491910 562896 491970
rect 563036 491910 563096 491970
rect 563236 491910 563296 491970
rect 563436 491910 563496 491970
rect 563636 491910 563696 491970
rect 563836 491910 563896 491970
rect 564036 491910 564096 491970
rect 564236 491910 564296 491970
rect 564436 491910 564496 491970
rect 564636 491910 564696 491970
rect 564836 491910 564896 491970
rect 565036 491910 565096 491970
rect 565236 491910 565296 491970
rect 565436 491910 565496 491970
rect 565636 491910 565696 491970
rect 574934 491880 575026 491984
rect 575228 491684 575288 491744
rect 575428 491684 575488 491744
rect 575628 491684 575688 491744
rect 575828 491684 575888 491744
rect 576028 491684 576088 491744
rect 576228 491684 576288 491744
rect 576428 491684 576488 491744
rect 576628 491684 576688 491744
rect 576828 491684 576888 491744
rect 577028 491684 577088 491744
rect 577228 491684 577288 491744
rect 577428 491684 577488 491744
rect 577628 491684 577688 491744
rect 577828 491684 577888 491744
rect 578028 491684 578088 491744
rect 578228 491684 578288 491744
rect 578428 491684 578488 491744
rect 578628 491684 578688 491744
rect 578828 491684 578888 491744
rect 579028 491684 579088 491744
rect 579228 491684 579288 491744
rect 579428 491684 579488 491744
rect 579628 491684 579688 491744
rect 579828 491684 579888 491744
rect 580028 491684 580088 491744
rect 580228 491684 580288 491744
rect 560772 404648 560832 404708
rect 560972 404648 561032 404708
rect 561172 404648 561232 404708
rect 561372 404648 561432 404708
rect 561572 404648 561632 404708
rect 561772 404648 561832 404708
rect 561972 404648 562032 404708
rect 562172 404648 562232 404708
rect 562372 404648 562432 404708
rect 562572 404648 562632 404708
rect 562772 404648 562832 404708
rect 562972 404648 563032 404708
rect 563172 404648 563232 404708
rect 563372 404648 563432 404708
rect 563572 404648 563632 404708
rect 563772 404648 563832 404708
rect 563972 404648 564032 404708
rect 564172 404648 564232 404708
rect 564372 404648 564432 404708
rect 564572 404648 564632 404708
rect 564772 404648 564832 404708
rect 564972 404648 565032 404708
rect 565172 404648 565232 404708
rect 565372 404648 565432 404708
rect 565572 404648 565632 404708
rect 574506 404688 574566 404748
rect 574706 404688 574766 404748
rect 574906 404688 574966 404748
rect 575106 404688 575166 404748
rect 575306 404688 575366 404748
rect 575506 404688 575566 404748
rect 575706 404688 575766 404748
rect 575906 404688 575966 404748
rect 576106 404688 576166 404748
rect 576306 404688 576366 404748
rect 576506 404688 576566 404748
rect 576706 404688 576766 404748
rect 576906 404688 576966 404748
rect 577106 404688 577166 404748
rect 577306 404688 577366 404748
rect 577506 404688 577566 404748
rect 577706 404688 577766 404748
rect 577906 404688 577966 404748
rect 578106 404688 578166 404748
rect 578306 404688 578366 404748
rect 578506 404688 578566 404748
rect 578706 404688 578766 404748
rect 578906 404688 578966 404748
rect 579106 404688 579166 404748
rect 579306 404688 579366 404748
rect 579506 404688 579566 404748
rect 560276 403190 560408 403340
rect 560597 403310 560631 404286
rect 560855 403310 560889 404286
rect 561113 403310 561147 404286
rect 561371 403310 561405 404286
rect 561629 403310 561663 404286
rect 561887 403310 561921 404286
rect 562145 403310 562179 404286
rect 562403 403310 562437 404286
rect 562661 403310 562695 404286
rect 562919 403310 562953 404286
rect 563177 403310 563211 404286
rect 563435 403310 563469 404286
rect 563693 403310 563727 404286
rect 563951 403310 563985 404286
rect 564209 403310 564243 404286
rect 564467 403310 564501 404286
rect 564725 403310 564759 404286
rect 564983 403310 565017 404286
rect 565241 403310 565275 404286
rect 565499 403310 565533 404286
rect 565757 403310 565791 404286
rect 566010 403178 566170 403286
rect 574495 403350 574529 404326
rect 574753 403350 574787 404326
rect 575011 403350 575045 404326
rect 575269 403350 575303 404326
rect 575527 403350 575561 404326
rect 575785 403350 575819 404326
rect 576043 403350 576077 404326
rect 576301 403350 576335 404326
rect 576559 403350 576593 404326
rect 576817 403350 576851 404326
rect 577075 403350 577109 404326
rect 577333 403350 577367 404326
rect 577591 403350 577625 404326
rect 577849 403350 577883 404326
rect 578107 403350 578141 404326
rect 578365 403350 578399 404326
rect 578623 403350 578657 404326
rect 578881 403350 578915 404326
rect 579139 403350 579173 404326
rect 579397 403350 579431 404326
rect 579655 403350 579689 404326
rect 579820 403154 579910 403242
rect 574212 403004 574304 403108
rect 560772 402768 560832 402828
rect 560972 402768 561032 402828
rect 561172 402768 561232 402828
rect 561372 402768 561432 402828
rect 561572 402768 561632 402828
rect 561772 402768 561832 402828
rect 561972 402768 562032 402828
rect 562172 402768 562232 402828
rect 562372 402768 562432 402828
rect 562572 402768 562632 402828
rect 562772 402768 562832 402828
rect 562972 402768 563032 402828
rect 563172 402768 563232 402828
rect 563372 402768 563432 402828
rect 563572 402768 563632 402828
rect 563772 402768 563832 402828
rect 563972 402768 564032 402828
rect 564172 402768 564232 402828
rect 564372 402768 564432 402828
rect 564572 402768 564632 402828
rect 564772 402768 564832 402828
rect 564972 402768 565032 402828
rect 565172 402768 565232 402828
rect 565372 402768 565432 402828
rect 565572 402768 565632 402828
rect 574506 402808 574566 402868
rect 574706 402808 574766 402868
rect 574906 402808 574966 402868
rect 575106 402808 575166 402868
rect 575306 402808 575366 402868
rect 575506 402808 575566 402868
rect 575706 402808 575766 402868
rect 575906 402808 575966 402868
rect 576106 402808 576166 402868
rect 576306 402808 576366 402868
rect 576506 402808 576566 402868
rect 576706 402808 576766 402868
rect 576906 402808 576966 402868
rect 577106 402808 577166 402868
rect 577306 402808 577366 402868
rect 577506 402808 577566 402868
rect 577706 402808 577766 402868
rect 577906 402808 577966 402868
rect 578106 402808 578166 402868
rect 578306 402808 578366 402868
rect 578506 402808 578566 402868
rect 578706 402808 578766 402868
rect 578906 402808 578966 402868
rect 579106 402808 579166 402868
rect 579306 402808 579366 402868
rect 579506 402808 579566 402868
rect 560728 359330 560788 359390
rect 560928 359330 560988 359390
rect 561128 359330 561188 359390
rect 561328 359330 561388 359390
rect 561528 359330 561588 359390
rect 561728 359330 561788 359390
rect 561928 359330 561988 359390
rect 562128 359330 562188 359390
rect 562328 359330 562388 359390
rect 562528 359330 562588 359390
rect 562728 359330 562788 359390
rect 562928 359330 562988 359390
rect 563128 359330 563188 359390
rect 563328 359330 563388 359390
rect 563528 359330 563588 359390
rect 563728 359330 563788 359390
rect 563928 359330 563988 359390
rect 564128 359330 564188 359390
rect 564328 359330 564388 359390
rect 564528 359330 564588 359390
rect 564728 359330 564788 359390
rect 564928 359330 564988 359390
rect 565128 359330 565188 359390
rect 565328 359330 565388 359390
rect 565528 359330 565588 359390
rect 574702 359260 574762 359320
rect 574902 359260 574962 359320
rect 575102 359260 575162 359320
rect 575302 359260 575362 359320
rect 575502 359260 575562 359320
rect 575702 359260 575762 359320
rect 575902 359260 575962 359320
rect 576102 359260 576162 359320
rect 576302 359260 576362 359320
rect 576502 359260 576562 359320
rect 576702 359260 576762 359320
rect 576902 359260 576962 359320
rect 577102 359260 577162 359320
rect 577302 359260 577362 359320
rect 577502 359260 577562 359320
rect 577702 359260 577762 359320
rect 577902 359260 577962 359320
rect 578102 359260 578162 359320
rect 578302 359260 578362 359320
rect 578502 359260 578562 359320
rect 578702 359260 578762 359320
rect 578902 359260 578962 359320
rect 579102 359260 579162 359320
rect 579302 359260 579362 359320
rect 579502 359260 579562 359320
rect 579702 359260 579762 359320
rect 560232 357872 560364 358022
rect 560553 357992 560587 358968
rect 560811 357992 560845 358968
rect 561069 357992 561103 358968
rect 561327 357992 561361 358968
rect 561585 357992 561619 358968
rect 561843 357992 561877 358968
rect 562101 357992 562135 358968
rect 562359 357992 562393 358968
rect 562617 357992 562651 358968
rect 562875 357992 562909 358968
rect 563133 357992 563167 358968
rect 563391 357992 563425 358968
rect 563649 357992 563683 358968
rect 563907 357992 563941 358968
rect 564165 357992 564199 358968
rect 564423 357992 564457 358968
rect 564681 357992 564715 358968
rect 564939 357992 564973 358968
rect 565197 357992 565231 358968
rect 565455 357992 565489 358968
rect 565713 357992 565747 358968
rect 565966 357860 566126 357968
rect 574691 357922 574725 358898
rect 574949 357922 574983 358898
rect 575207 357922 575241 358898
rect 575465 357922 575499 358898
rect 575723 357922 575757 358898
rect 575981 357922 576015 358898
rect 576239 357922 576273 358898
rect 576497 357922 576531 358898
rect 576755 357922 576789 358898
rect 577013 357922 577047 358898
rect 577271 357922 577305 358898
rect 577529 357922 577563 358898
rect 577787 357922 577821 358898
rect 578045 357922 578079 358898
rect 578303 357922 578337 358898
rect 578561 357922 578595 358898
rect 578819 357922 578853 358898
rect 579077 357922 579111 358898
rect 579335 357922 579369 358898
rect 579593 357922 579627 358898
rect 579851 357922 579885 358898
rect 580016 357726 580106 357814
rect 574408 357576 574500 357680
rect 560728 357450 560788 357510
rect 560928 357450 560988 357510
rect 561128 357450 561188 357510
rect 561328 357450 561388 357510
rect 561528 357450 561588 357510
rect 561728 357450 561788 357510
rect 561928 357450 561988 357510
rect 562128 357450 562188 357510
rect 562328 357450 562388 357510
rect 562528 357450 562588 357510
rect 562728 357450 562788 357510
rect 562928 357450 562988 357510
rect 563128 357450 563188 357510
rect 563328 357450 563388 357510
rect 563528 357450 563588 357510
rect 563728 357450 563788 357510
rect 563928 357450 563988 357510
rect 564128 357450 564188 357510
rect 564328 357450 564388 357510
rect 564528 357450 564588 357510
rect 564728 357450 564788 357510
rect 564928 357450 564988 357510
rect 565128 357450 565188 357510
rect 565328 357450 565388 357510
rect 565528 357450 565588 357510
rect 574702 357380 574762 357440
rect 574902 357380 574962 357440
rect 575102 357380 575162 357440
rect 575302 357380 575362 357440
rect 575502 357380 575562 357440
rect 575702 357380 575762 357440
rect 575902 357380 575962 357440
rect 576102 357380 576162 357440
rect 576302 357380 576362 357440
rect 576502 357380 576562 357440
rect 576702 357380 576762 357440
rect 576902 357380 576962 357440
rect 577102 357380 577162 357440
rect 577302 357380 577362 357440
rect 577502 357380 577562 357440
rect 577702 357380 577762 357440
rect 577902 357380 577962 357440
rect 578102 357380 578162 357440
rect 578302 357380 578362 357440
rect 578502 357380 578562 357440
rect 578702 357380 578762 357440
rect 578902 357380 578962 357440
rect 579102 357380 579162 357440
rect 579302 357380 579362 357440
rect 579502 357380 579562 357440
rect 579702 357380 579762 357440
rect 575150 313092 575210 313152
rect 575350 313092 575410 313152
rect 575550 313092 575610 313152
rect 575750 313092 575810 313152
rect 575950 313092 576010 313152
rect 576150 313092 576210 313152
rect 576350 313092 576410 313152
rect 576550 313092 576610 313152
rect 576750 313092 576810 313152
rect 576950 313092 577010 313152
rect 577150 313092 577210 313152
rect 577350 313092 577410 313152
rect 577550 313092 577610 313152
rect 577750 313092 577810 313152
rect 577950 313092 578010 313152
rect 578150 313092 578210 313152
rect 578350 313092 578410 313152
rect 578550 313092 578610 313152
rect 578750 313092 578810 313152
rect 578950 313092 579010 313152
rect 579150 313092 579210 313152
rect 579350 313092 579410 313152
rect 579550 313092 579610 313152
rect 579750 313092 579810 313152
rect 579950 313092 580010 313152
rect 580150 313092 580210 313152
rect 560590 313022 560650 313082
rect 560790 313022 560850 313082
rect 560990 313022 561050 313082
rect 561190 313022 561250 313082
rect 561390 313022 561450 313082
rect 561590 313022 561650 313082
rect 561790 313022 561850 313082
rect 561990 313022 562050 313082
rect 562190 313022 562250 313082
rect 562390 313022 562450 313082
rect 562590 313022 562650 313082
rect 562790 313022 562850 313082
rect 562990 313022 563050 313082
rect 563190 313022 563250 313082
rect 563390 313022 563450 313082
rect 563590 313022 563650 313082
rect 563790 313022 563850 313082
rect 563990 313022 564050 313082
rect 564190 313022 564250 313082
rect 564390 313022 564450 313082
rect 564590 313022 564650 313082
rect 564790 313022 564850 313082
rect 564990 313022 565050 313082
rect 565190 313022 565250 313082
rect 565390 313022 565450 313082
rect 560094 311564 560226 311714
rect 560415 311684 560449 312660
rect 560673 311684 560707 312660
rect 560931 311684 560965 312660
rect 561189 311684 561223 312660
rect 561447 311684 561481 312660
rect 561705 311684 561739 312660
rect 561963 311684 561997 312660
rect 562221 311684 562255 312660
rect 562479 311684 562513 312660
rect 562737 311684 562771 312660
rect 562995 311684 563029 312660
rect 563253 311684 563287 312660
rect 563511 311684 563545 312660
rect 563769 311684 563803 312660
rect 564027 311684 564061 312660
rect 564285 311684 564319 312660
rect 564543 311684 564577 312660
rect 564801 311684 564835 312660
rect 565059 311684 565093 312660
rect 565317 311684 565351 312660
rect 565575 311684 565609 312660
rect 565828 311552 565988 311660
rect 575139 311754 575173 312730
rect 575397 311754 575431 312730
rect 575655 311754 575689 312730
rect 575913 311754 575947 312730
rect 576171 311754 576205 312730
rect 576429 311754 576463 312730
rect 576687 311754 576721 312730
rect 576945 311754 576979 312730
rect 577203 311754 577237 312730
rect 577461 311754 577495 312730
rect 577719 311754 577753 312730
rect 577977 311754 578011 312730
rect 578235 311754 578269 312730
rect 578493 311754 578527 312730
rect 578751 311754 578785 312730
rect 579009 311754 579043 312730
rect 579267 311754 579301 312730
rect 579525 311754 579559 312730
rect 579783 311754 579817 312730
rect 580041 311754 580075 312730
rect 580299 311754 580333 312730
rect 580464 311558 580554 311646
rect 574856 311408 574948 311512
rect 575150 311212 575210 311272
rect 575350 311212 575410 311272
rect 575550 311212 575610 311272
rect 575750 311212 575810 311272
rect 575950 311212 576010 311272
rect 576150 311212 576210 311272
rect 576350 311212 576410 311272
rect 576550 311212 576610 311272
rect 576750 311212 576810 311272
rect 576950 311212 577010 311272
rect 577150 311212 577210 311272
rect 577350 311212 577410 311272
rect 577550 311212 577610 311272
rect 577750 311212 577810 311272
rect 577950 311212 578010 311272
rect 578150 311212 578210 311272
rect 578350 311212 578410 311272
rect 578550 311212 578610 311272
rect 578750 311212 578810 311272
rect 578950 311212 579010 311272
rect 579150 311212 579210 311272
rect 579350 311212 579410 311272
rect 579550 311212 579610 311272
rect 579750 311212 579810 311272
rect 579950 311212 580010 311272
rect 580150 311212 580210 311272
rect 560590 311142 560650 311202
rect 560790 311142 560850 311202
rect 560990 311142 561050 311202
rect 561190 311142 561250 311202
rect 561390 311142 561450 311202
rect 561590 311142 561650 311202
rect 561790 311142 561850 311202
rect 561990 311142 562050 311202
rect 562190 311142 562250 311202
rect 562390 311142 562450 311202
rect 562590 311142 562650 311202
rect 562790 311142 562850 311202
rect 562990 311142 563050 311202
rect 563190 311142 563250 311202
rect 563390 311142 563450 311202
rect 563590 311142 563650 311202
rect 563790 311142 563850 311202
rect 563990 311142 564050 311202
rect 564190 311142 564250 311202
rect 564390 311142 564450 311202
rect 564590 311142 564650 311202
rect 564790 311142 564850 311202
rect 564990 311142 565050 311202
rect 565190 311142 565250 311202
rect 565390 311142 565450 311202
<< metal1 >>
rect 573584 494882 573796 494888
rect 565696 494762 573796 494882
rect 565696 493880 565816 494762
rect 566176 494126 566186 494310
rect 566408 494126 566418 494310
rect 560650 493850 565964 493880
rect 560650 493790 560836 493850
rect 560896 493790 561036 493850
rect 561096 493790 561236 493850
rect 561296 493790 561436 493850
rect 561496 493790 561636 493850
rect 561696 493790 561836 493850
rect 561896 493790 562036 493850
rect 562096 493790 562236 493850
rect 562296 493790 562436 493850
rect 562496 493790 562636 493850
rect 562696 493790 562836 493850
rect 562896 493790 563036 493850
rect 563096 493790 563236 493850
rect 563296 493790 563436 493850
rect 563496 493790 563636 493850
rect 563696 493790 563836 493850
rect 563896 493790 564036 493850
rect 564096 493790 564236 493850
rect 564296 493790 564436 493850
rect 564496 493790 564636 493850
rect 564696 493790 564836 493850
rect 564896 493790 565036 493850
rect 565096 493790 565236 493850
rect 565296 493790 565436 493850
rect 565496 493790 565636 493850
rect 565696 493790 565964 493850
rect 560650 493760 565964 493790
rect 560655 493428 560701 493440
rect 559792 492548 560110 492554
rect 559788 492536 560448 492548
rect 559788 492324 559802 492536
rect 560012 492512 560448 492536
rect 560012 492482 560486 492512
rect 560012 492332 560340 492482
rect 560472 492332 560486 492482
rect 560655 492452 560661 493428
rect 560695 492452 560701 493428
rect 560655 492440 560701 492452
rect 560913 493428 560959 493440
rect 560913 492452 560919 493428
rect 560953 492452 560959 493428
rect 560913 492440 560959 492452
rect 561171 493428 561217 493440
rect 561171 492452 561177 493428
rect 561211 492452 561217 493428
rect 561171 492440 561217 492452
rect 561429 493428 561475 493440
rect 561429 492452 561435 493428
rect 561469 492452 561475 493428
rect 561429 492440 561475 492452
rect 561687 493428 561733 493440
rect 561687 492452 561693 493428
rect 561727 492452 561733 493428
rect 561687 492440 561733 492452
rect 561945 493428 561991 493440
rect 561945 492452 561951 493428
rect 561985 492452 561991 493428
rect 561945 492440 561991 492452
rect 562203 493428 562249 493440
rect 562203 492452 562209 493428
rect 562243 492452 562249 493428
rect 562203 492440 562249 492452
rect 562461 493428 562507 493440
rect 562461 492452 562467 493428
rect 562501 492452 562507 493428
rect 562461 492440 562507 492452
rect 562719 493428 562765 493440
rect 562719 492452 562725 493428
rect 562759 492452 562765 493428
rect 562719 492440 562765 492452
rect 562977 493428 563023 493440
rect 562977 492452 562983 493428
rect 563017 492452 563023 493428
rect 562977 492440 563023 492452
rect 563235 493428 563281 493440
rect 563235 492452 563241 493428
rect 563275 492452 563281 493428
rect 563235 492440 563281 492452
rect 563493 493428 563539 493440
rect 563493 492452 563499 493428
rect 563533 492452 563539 493428
rect 563493 492440 563539 492452
rect 563751 493428 563797 493440
rect 563751 492452 563757 493428
rect 563791 492452 563797 493428
rect 563751 492440 563797 492452
rect 564009 493428 564055 493440
rect 564009 492452 564015 493428
rect 564049 492452 564055 493428
rect 564009 492440 564055 492452
rect 564267 493428 564313 493440
rect 564267 492452 564273 493428
rect 564307 492452 564313 493428
rect 564267 492440 564313 492452
rect 564525 493428 564571 493440
rect 564525 492452 564531 493428
rect 564565 492452 564571 493428
rect 564525 492440 564571 492452
rect 564783 493428 564829 493440
rect 564783 492452 564789 493428
rect 564823 492452 564829 493428
rect 564783 492440 564829 492452
rect 565041 493428 565087 493440
rect 565041 492452 565047 493428
rect 565081 492452 565087 493428
rect 565041 492440 565087 492452
rect 565299 493428 565345 493440
rect 565299 492452 565305 493428
rect 565339 492452 565345 493428
rect 565299 492440 565345 492452
rect 565557 493428 565603 493440
rect 565557 492452 565563 493428
rect 565597 492452 565603 493428
rect 565557 492440 565603 492452
rect 565815 493428 565861 493440
rect 565815 492452 565821 493428
rect 565855 492452 565861 493428
rect 566196 492512 566404 494126
rect 573584 493658 573796 494762
rect 580846 494136 580856 494348
rect 581040 494136 581050 494348
rect 573584 493654 573980 493658
rect 565815 492440 565861 492452
rect 566034 492452 566404 492512
rect 573576 493624 580556 493654
rect 573576 493564 575228 493624
rect 575288 493564 575428 493624
rect 575488 493564 575628 493624
rect 575688 493564 575828 493624
rect 575888 493564 576028 493624
rect 576088 493564 576228 493624
rect 576288 493564 576428 493624
rect 576488 493564 576628 493624
rect 576688 493564 576828 493624
rect 576888 493564 577028 493624
rect 577088 493564 577228 493624
rect 577288 493564 577428 493624
rect 577488 493564 577628 493624
rect 577688 493564 577828 493624
rect 577888 493564 578028 493624
rect 578088 493564 578228 493624
rect 578288 493564 578428 493624
rect 578488 493564 578628 493624
rect 578688 493564 578828 493624
rect 578888 493564 579028 493624
rect 579088 493564 579228 493624
rect 579288 493564 579428 493624
rect 579488 493564 579628 493624
rect 579688 493564 579828 493624
rect 579888 493564 580028 493624
rect 580088 493564 580228 493624
rect 580288 493564 580556 493624
rect 573576 493534 580556 493564
rect 560012 492324 560486 492332
rect 559788 492304 560486 492324
rect 566034 492428 566526 492452
rect 566034 492320 566074 492428
rect 566234 492320 566526 492428
rect 566034 492304 566526 492320
rect 559788 492000 559996 492304
rect 573576 492196 573796 493534
rect 575211 493202 575257 493214
rect 575211 492226 575217 493202
rect 575251 492226 575257 493202
rect 575211 492214 575257 492226
rect 575469 493202 575515 493214
rect 575469 492226 575475 493202
rect 575509 492226 575515 493202
rect 575469 492214 575515 492226
rect 575727 493202 575773 493214
rect 575727 492226 575733 493202
rect 575767 492226 575773 493202
rect 575727 492214 575773 492226
rect 575985 493202 576031 493214
rect 575985 492226 575991 493202
rect 576025 492226 576031 493202
rect 575985 492214 576031 492226
rect 576243 493202 576289 493214
rect 576243 492226 576249 493202
rect 576283 492226 576289 493202
rect 576243 492214 576289 492226
rect 576501 493202 576547 493214
rect 576501 492226 576507 493202
rect 576541 492226 576547 493202
rect 576501 492214 576547 492226
rect 576759 493202 576805 493214
rect 576759 492226 576765 493202
rect 576799 492226 576805 493202
rect 576759 492214 576805 492226
rect 577017 493202 577063 493214
rect 577017 492226 577023 493202
rect 577057 492226 577063 493202
rect 577017 492214 577063 492226
rect 577275 493202 577321 493214
rect 577275 492226 577281 493202
rect 577315 492226 577321 493202
rect 577275 492214 577321 492226
rect 577533 493202 577579 493214
rect 577533 492226 577539 493202
rect 577573 492226 577579 493202
rect 577533 492214 577579 492226
rect 577791 493202 577837 493214
rect 577791 492226 577797 493202
rect 577831 492226 577837 493202
rect 577791 492214 577837 492226
rect 578049 493202 578095 493214
rect 578049 492226 578055 493202
rect 578089 492226 578095 493202
rect 578049 492214 578095 492226
rect 578307 493202 578353 493214
rect 578307 492226 578313 493202
rect 578347 492226 578353 493202
rect 578307 492214 578353 492226
rect 578565 493202 578611 493214
rect 578565 492226 578571 493202
rect 578605 492226 578611 493202
rect 578565 492214 578611 492226
rect 578823 493202 578869 493214
rect 578823 492226 578829 493202
rect 578863 492226 578869 493202
rect 578823 492214 578869 492226
rect 579081 493202 579127 493214
rect 579081 492226 579087 493202
rect 579121 492226 579127 493202
rect 579081 492214 579127 492226
rect 579339 493202 579385 493214
rect 579339 492226 579345 493202
rect 579379 492226 579385 493202
rect 579339 492214 579385 492226
rect 579597 493202 579643 493214
rect 579597 492226 579603 493202
rect 579637 492226 579643 493202
rect 579597 492214 579643 492226
rect 579855 493202 579901 493214
rect 579855 492226 579861 493202
rect 579895 492226 579901 493202
rect 579855 492214 579901 492226
rect 580113 493202 580159 493214
rect 580113 492226 580119 493202
rect 580153 492226 580159 493202
rect 580113 492214 580159 492226
rect 580371 493202 580417 493214
rect 580371 492226 580377 493202
rect 580411 492226 580417 493202
rect 580371 492214 580417 492226
rect 573506 492160 573954 492196
rect 559788 491970 565964 492000
rect 559788 491910 560836 491970
rect 560896 491910 561036 491970
rect 561096 491910 561236 491970
rect 561296 491910 561436 491970
rect 561496 491910 561636 491970
rect 561696 491910 561836 491970
rect 561896 491910 562036 491970
rect 562096 491910 562236 491970
rect 562296 491910 562436 491970
rect 562496 491910 562636 491970
rect 562696 491910 562836 491970
rect 562896 491910 563036 491970
rect 563096 491910 563236 491970
rect 563296 491910 563436 491970
rect 563496 491910 563636 491970
rect 563696 491910 563836 491970
rect 563896 491910 564036 491970
rect 564096 491910 564236 491970
rect 564296 491910 564436 491970
rect 564496 491910 564636 491970
rect 564696 491910 564836 491970
rect 564896 491910 565036 491970
rect 565096 491910 565236 491970
rect 565296 491910 565436 491970
rect 565496 491910 565636 491970
rect 565696 491910 565964 491970
rect 559788 491884 565964 491910
rect 559834 491880 565964 491884
rect 573506 491888 573564 492160
rect 573874 492076 573954 492160
rect 580852 492130 581040 494136
rect 580530 492118 581040 492130
rect 573874 491984 575038 492076
rect 580530 492030 580542 492118
rect 580632 492030 581040 492118
rect 580530 492026 581040 492030
rect 580530 492024 580644 492026
rect 573874 491888 574934 491984
rect 573506 491880 574934 491888
rect 575026 491948 575038 491984
rect 575026 491880 575034 491948
rect 565726 491604 565846 491880
rect 573506 491868 575034 491880
rect 575170 491744 580556 491774
rect 575170 491684 575228 491744
rect 575288 491684 575428 491744
rect 575488 491684 575628 491744
rect 575688 491684 575828 491744
rect 575888 491684 576028 491744
rect 576088 491684 576228 491744
rect 576288 491684 576428 491744
rect 576488 491684 576628 491744
rect 576688 491684 576828 491744
rect 576888 491684 577028 491744
rect 577088 491684 577228 491744
rect 577288 491684 577428 491744
rect 577488 491684 577628 491744
rect 577688 491684 577828 491744
rect 577888 491684 578028 491744
rect 578088 491684 578228 491744
rect 578288 491684 578428 491744
rect 578488 491684 578628 491744
rect 578688 491684 578828 491744
rect 578888 491684 579028 491744
rect 579088 491684 579228 491744
rect 579288 491684 579428 491744
rect 579488 491684 579628 491744
rect 579688 491684 579828 491744
rect 579888 491684 580028 491744
rect 580088 491684 580228 491744
rect 580288 491684 580556 491744
rect 575170 491654 580556 491684
rect 575288 491604 575408 491654
rect 565726 491484 575408 491604
rect 560592 406072 573714 406192
rect 560592 404738 560712 406072
rect 566254 405476 566462 405488
rect 566246 405258 566256 405476
rect 566462 405258 566472 405476
rect 560586 404708 565944 404738
rect 560586 404648 560772 404708
rect 560832 404648 560972 404708
rect 561032 404648 561172 404708
rect 561232 404648 561372 404708
rect 561432 404648 561572 404708
rect 561632 404648 561772 404708
rect 561832 404648 561972 404708
rect 562032 404648 562172 404708
rect 562232 404648 562372 404708
rect 562432 404648 562572 404708
rect 562632 404648 562772 404708
rect 562832 404648 562972 404708
rect 563032 404648 563172 404708
rect 563232 404648 563372 404708
rect 563432 404648 563572 404708
rect 563632 404648 563772 404708
rect 563832 404648 563972 404708
rect 564032 404648 564172 404708
rect 564232 404648 564372 404708
rect 564432 404648 564572 404708
rect 564632 404648 564772 404708
rect 564832 404648 564972 404708
rect 565032 404648 565172 404708
rect 565232 404648 565372 404708
rect 565432 404648 565572 404708
rect 565632 404648 565944 404708
rect 560586 404618 565944 404648
rect 560591 404286 560637 404298
rect 559706 403370 560120 403492
rect 559706 403368 560422 403370
rect 559706 403280 559736 403368
rect 559704 403192 559736 403280
rect 559926 403340 560422 403368
rect 559926 403192 560276 403340
rect 559704 403190 560276 403192
rect 560408 403190 560422 403340
rect 560591 403310 560597 404286
rect 560631 403310 560637 404286
rect 560591 403298 560637 403310
rect 560849 404286 560895 404298
rect 560849 403310 560855 404286
rect 560889 403310 560895 404286
rect 560849 403298 560895 403310
rect 561107 404286 561153 404298
rect 561107 403310 561113 404286
rect 561147 403310 561153 404286
rect 561107 403298 561153 403310
rect 561365 404286 561411 404298
rect 561365 403310 561371 404286
rect 561405 403310 561411 404286
rect 561365 403298 561411 403310
rect 561623 404286 561669 404298
rect 561623 403310 561629 404286
rect 561663 403310 561669 404286
rect 561623 403298 561669 403310
rect 561881 404286 561927 404298
rect 561881 403310 561887 404286
rect 561921 403310 561927 404286
rect 561881 403298 561927 403310
rect 562139 404286 562185 404298
rect 562139 403310 562145 404286
rect 562179 403310 562185 404286
rect 562139 403298 562185 403310
rect 562397 404286 562443 404298
rect 562397 403310 562403 404286
rect 562437 403310 562443 404286
rect 562397 403298 562443 403310
rect 562655 404286 562701 404298
rect 562655 403310 562661 404286
rect 562695 403310 562701 404286
rect 562655 403298 562701 403310
rect 562913 404286 562959 404298
rect 562913 403310 562919 404286
rect 562953 403310 562959 404286
rect 562913 403298 562959 403310
rect 563171 404286 563217 404298
rect 563171 403310 563177 404286
rect 563211 403310 563217 404286
rect 563171 403298 563217 403310
rect 563429 404286 563475 404298
rect 563429 403310 563435 404286
rect 563469 403310 563475 404286
rect 563429 403298 563475 403310
rect 563687 404286 563733 404298
rect 563687 403310 563693 404286
rect 563727 403310 563733 404286
rect 563687 403298 563733 403310
rect 563945 404286 563991 404298
rect 563945 403310 563951 404286
rect 563985 403310 563991 404286
rect 563945 403298 563991 403310
rect 564203 404286 564249 404298
rect 564203 403310 564209 404286
rect 564243 403310 564249 404286
rect 564203 403298 564249 403310
rect 564461 404286 564507 404298
rect 564461 403310 564467 404286
rect 564501 403310 564507 404286
rect 564461 403298 564507 403310
rect 564719 404286 564765 404298
rect 564719 403310 564725 404286
rect 564759 403310 564765 404286
rect 564719 403298 564765 403310
rect 564977 404286 565023 404298
rect 564977 403310 564983 404286
rect 565017 403310 565023 404286
rect 564977 403298 565023 403310
rect 565235 404286 565281 404298
rect 565235 403310 565241 404286
rect 565275 403310 565281 404286
rect 565235 403298 565281 403310
rect 565493 404286 565539 404298
rect 565493 403310 565499 404286
rect 565533 403310 565539 404286
rect 565493 403298 565539 403310
rect 565751 404286 565797 404298
rect 565751 403310 565757 404286
rect 565791 403310 565797 404286
rect 566254 403310 566462 405258
rect 573512 404778 573714 406072
rect 580076 405402 580180 405420
rect 580064 405292 580074 405402
rect 580182 405292 580192 405402
rect 573512 404748 579834 404778
rect 573512 404688 574506 404748
rect 574566 404688 574706 404748
rect 574766 404688 574906 404748
rect 574966 404688 575106 404748
rect 575166 404688 575306 404748
rect 575366 404688 575506 404748
rect 575566 404688 575706 404748
rect 575766 404688 575906 404748
rect 575966 404688 576106 404748
rect 576166 404688 576306 404748
rect 576366 404688 576506 404748
rect 576566 404688 576706 404748
rect 576766 404688 576906 404748
rect 576966 404688 577106 404748
rect 577166 404688 577306 404748
rect 577366 404688 577506 404748
rect 577566 404688 577706 404748
rect 577766 404688 577906 404748
rect 577966 404688 578106 404748
rect 578166 404688 578306 404748
rect 578366 404688 578506 404748
rect 578566 404688 578706 404748
rect 578766 404688 578906 404748
rect 578966 404688 579106 404748
rect 579166 404688 579306 404748
rect 579366 404688 579506 404748
rect 579566 404688 579834 404748
rect 573512 404658 579834 404688
rect 573512 403353 573672 404658
rect 574489 404326 574535 404338
rect 565751 403298 565797 403310
rect 559704 403162 560422 403190
rect 565994 403286 566462 403310
rect 565994 403178 566010 403286
rect 566170 403178 566462 403286
rect 565994 403162 566462 403178
rect 573509 403312 574144 403353
rect 574489 403350 574495 404326
rect 574529 403350 574535 404326
rect 574489 403338 574535 403350
rect 574747 404326 574793 404338
rect 574747 403350 574753 404326
rect 574787 403350 574793 404326
rect 574747 403338 574793 403350
rect 575005 404326 575051 404338
rect 575005 403350 575011 404326
rect 575045 403350 575051 404326
rect 575005 403338 575051 403350
rect 575263 404326 575309 404338
rect 575263 403350 575269 404326
rect 575303 403350 575309 404326
rect 575263 403338 575309 403350
rect 575521 404326 575567 404338
rect 575521 403350 575527 404326
rect 575561 403350 575567 404326
rect 575521 403338 575567 403350
rect 575779 404326 575825 404338
rect 575779 403350 575785 404326
rect 575819 403350 575825 404326
rect 575779 403338 575825 403350
rect 576037 404326 576083 404338
rect 576037 403350 576043 404326
rect 576077 403350 576083 404326
rect 576037 403338 576083 403350
rect 576295 404326 576341 404338
rect 576295 403350 576301 404326
rect 576335 403350 576341 404326
rect 576295 403338 576341 403350
rect 576553 404326 576599 404338
rect 576553 403350 576559 404326
rect 576593 403350 576599 404326
rect 576553 403338 576599 403350
rect 576811 404326 576857 404338
rect 576811 403350 576817 404326
rect 576851 403350 576857 404326
rect 576811 403338 576857 403350
rect 577069 404326 577115 404338
rect 577069 403350 577075 404326
rect 577109 403350 577115 404326
rect 577069 403338 577115 403350
rect 577327 404326 577373 404338
rect 577327 403350 577333 404326
rect 577367 403350 577373 404326
rect 577327 403338 577373 403350
rect 577585 404326 577631 404338
rect 577585 403350 577591 404326
rect 577625 403350 577631 404326
rect 577585 403338 577631 403350
rect 577843 404326 577889 404338
rect 577843 403350 577849 404326
rect 577883 403350 577889 404326
rect 577843 403338 577889 403350
rect 578101 404326 578147 404338
rect 578101 403350 578107 404326
rect 578141 403350 578147 404326
rect 578101 403338 578147 403350
rect 578359 404326 578405 404338
rect 578359 403350 578365 404326
rect 578399 403350 578405 404326
rect 578359 403338 578405 403350
rect 578617 404326 578663 404338
rect 578617 403350 578623 404326
rect 578657 403350 578663 404326
rect 578617 403338 578663 403350
rect 578875 404326 578921 404338
rect 578875 403350 578881 404326
rect 578915 403350 578921 404326
rect 578875 403338 578921 403350
rect 579133 404326 579179 404338
rect 579133 403350 579139 404326
rect 579173 403350 579179 404326
rect 579133 403338 579179 403350
rect 579391 404326 579437 404338
rect 579391 403350 579397 404326
rect 579431 403350 579437 404326
rect 579391 403338 579437 403350
rect 579649 404326 579695 404338
rect 579649 403350 579655 404326
rect 579689 403350 579695 404326
rect 579649 403338 579695 403350
rect 559704 402858 560146 403162
rect 573509 403107 573538 403312
rect 573510 402980 573538 403107
rect 573888 403120 574144 403312
rect 580076 403254 580180 405292
rect 579808 403242 580180 403254
rect 579808 403154 579820 403242
rect 579910 403154 580180 403242
rect 579808 403150 580180 403154
rect 579808 403148 579922 403150
rect 573888 403108 574312 403120
rect 573888 403004 574212 403108
rect 574304 403004 574312 403108
rect 573888 402992 574312 403004
rect 573888 402980 574196 402992
rect 573510 402956 574196 402980
rect 574448 402868 579834 402898
rect 574448 402858 574506 402868
rect 559704 402828 574506 402858
rect 559704 402768 560772 402828
rect 560832 402768 560972 402828
rect 561032 402768 561172 402828
rect 561232 402768 561372 402828
rect 561432 402768 561572 402828
rect 561632 402768 561772 402828
rect 561832 402768 561972 402828
rect 562032 402768 562172 402828
rect 562232 402768 562372 402828
rect 562432 402768 562572 402828
rect 562632 402768 562772 402828
rect 562832 402768 562972 402828
rect 563032 402768 563172 402828
rect 563232 402768 563372 402828
rect 563432 402768 563572 402828
rect 563632 402768 563772 402828
rect 563832 402768 563972 402828
rect 564032 402768 564172 402828
rect 564232 402768 564372 402828
rect 564432 402768 564572 402828
rect 564632 402768 564772 402828
rect 564832 402768 564972 402828
rect 565032 402768 565172 402828
rect 565232 402768 565372 402828
rect 565432 402768 565572 402828
rect 565632 402808 574506 402828
rect 574566 402808 574706 402868
rect 574766 402808 574906 402868
rect 574966 402808 575106 402868
rect 575166 402808 575306 402868
rect 575366 402808 575506 402868
rect 575566 402808 575706 402868
rect 575766 402808 575906 402868
rect 575966 402808 576106 402868
rect 576166 402808 576306 402868
rect 576366 402808 576506 402868
rect 576566 402808 576706 402868
rect 576766 402808 576906 402868
rect 576966 402808 577106 402868
rect 577166 402808 577306 402868
rect 577366 402808 577506 402868
rect 577566 402808 577706 402868
rect 577766 402808 577906 402868
rect 577966 402808 578106 402868
rect 578166 402808 578306 402868
rect 578366 402808 578506 402868
rect 578566 402808 578706 402868
rect 578766 402808 578906 402868
rect 578966 402808 579106 402868
rect 579166 402808 579306 402868
rect 579366 402808 579506 402868
rect 579566 402808 579834 402868
rect 565632 402778 579834 402808
rect 565632 402768 574718 402778
rect 559704 402738 574718 402768
rect 565736 360464 573796 360584
rect 565736 359420 565856 360464
rect 566270 359978 566494 360002
rect 566264 359786 566274 359978
rect 566500 359786 566510 359978
rect 560542 359390 565856 359420
rect 560542 359330 560728 359390
rect 560788 359330 560928 359390
rect 560988 359330 561128 359390
rect 561188 359330 561328 359390
rect 561388 359330 561528 359390
rect 561588 359330 561728 359390
rect 561788 359330 561928 359390
rect 561988 359330 562128 359390
rect 562188 359330 562328 359390
rect 562388 359330 562528 359390
rect 562588 359330 562728 359390
rect 562788 359330 562928 359390
rect 562988 359330 563128 359390
rect 563188 359330 563328 359390
rect 563388 359330 563528 359390
rect 563588 359330 563728 359390
rect 563788 359330 563928 359390
rect 563988 359330 564128 359390
rect 564188 359330 564328 359390
rect 564388 359330 564528 359390
rect 564588 359330 564728 359390
rect 564788 359330 564928 359390
rect 564988 359330 565128 359390
rect 565188 359330 565328 359390
rect 565388 359330 565528 359390
rect 565588 359330 565856 359390
rect 560542 359300 565856 359330
rect 560547 358968 560593 358980
rect 559702 357844 559712 358052
rect 559920 358022 560378 358052
rect 559920 357872 560232 358022
rect 560364 357872 560378 358022
rect 560547 357992 560553 358968
rect 560587 357992 560593 358968
rect 560547 357980 560593 357992
rect 560805 358968 560851 358980
rect 560805 357992 560811 358968
rect 560845 357992 560851 358968
rect 560805 357980 560851 357992
rect 561063 358968 561109 358980
rect 561063 357992 561069 358968
rect 561103 357992 561109 358968
rect 561063 357980 561109 357992
rect 561321 358968 561367 358980
rect 561321 357992 561327 358968
rect 561361 357992 561367 358968
rect 561321 357980 561367 357992
rect 561579 358968 561625 358980
rect 561579 357992 561585 358968
rect 561619 357992 561625 358968
rect 561579 357980 561625 357992
rect 561837 358968 561883 358980
rect 561837 357992 561843 358968
rect 561877 357992 561883 358968
rect 561837 357980 561883 357992
rect 562095 358968 562141 358980
rect 562095 357992 562101 358968
rect 562135 357992 562141 358968
rect 562095 357980 562141 357992
rect 562353 358968 562399 358980
rect 562353 357992 562359 358968
rect 562393 357992 562399 358968
rect 562353 357980 562399 357992
rect 562611 358968 562657 358980
rect 562611 357992 562617 358968
rect 562651 357992 562657 358968
rect 562611 357980 562657 357992
rect 562869 358968 562915 358980
rect 562869 357992 562875 358968
rect 562909 357992 562915 358968
rect 562869 357980 562915 357992
rect 563127 358968 563173 358980
rect 563127 357992 563133 358968
rect 563167 357992 563173 358968
rect 563127 357980 563173 357992
rect 563385 358968 563431 358980
rect 563385 357992 563391 358968
rect 563425 357992 563431 358968
rect 563385 357980 563431 357992
rect 563643 358968 563689 358980
rect 563643 357992 563649 358968
rect 563683 357992 563689 358968
rect 563643 357980 563689 357992
rect 563901 358968 563947 358980
rect 563901 357992 563907 358968
rect 563941 357992 563947 358968
rect 563901 357980 563947 357992
rect 564159 358968 564205 358980
rect 564159 357992 564165 358968
rect 564199 357992 564205 358968
rect 564159 357980 564205 357992
rect 564417 358968 564463 358980
rect 564417 357992 564423 358968
rect 564457 357992 564463 358968
rect 564417 357980 564463 357992
rect 564675 358968 564721 358980
rect 564675 357992 564681 358968
rect 564715 357992 564721 358968
rect 564675 357980 564721 357992
rect 564933 358968 564979 358980
rect 564933 357992 564939 358968
rect 564973 357992 564979 358968
rect 564933 357980 564979 357992
rect 565191 358968 565237 358980
rect 565191 357992 565197 358968
rect 565231 357992 565237 358968
rect 565191 357980 565237 357992
rect 565449 358968 565495 358980
rect 565449 357992 565455 358968
rect 565489 357992 565495 358968
rect 565449 357980 565495 357992
rect 565707 358968 565753 358980
rect 565707 357992 565713 358968
rect 565747 357992 565753 358968
rect 566270 357992 566494 359786
rect 573588 359350 573796 360464
rect 580252 359906 580356 359934
rect 580242 359786 580252 359906
rect 580358 359786 580368 359906
rect 573588 359320 580030 359350
rect 573588 359260 574702 359320
rect 574762 359260 574902 359320
rect 574962 359260 575102 359320
rect 575162 359260 575302 359320
rect 575362 359260 575502 359320
rect 575562 359260 575702 359320
rect 575762 359260 575902 359320
rect 575962 359260 576102 359320
rect 576162 359260 576302 359320
rect 576362 359260 576502 359320
rect 576562 359260 576702 359320
rect 576762 359260 576902 359320
rect 576962 359260 577102 359320
rect 577162 359260 577302 359320
rect 577362 359260 577502 359320
rect 577562 359260 577702 359320
rect 577762 359260 577902 359320
rect 577962 359260 578102 359320
rect 578162 359260 578302 359320
rect 578362 359260 578502 359320
rect 578562 359260 578702 359320
rect 578762 359260 578902 359320
rect 578962 359260 579102 359320
rect 579162 359260 579302 359320
rect 579362 359260 579502 359320
rect 579562 359260 579702 359320
rect 579762 359260 580030 359320
rect 573588 359256 580030 359260
rect 565707 357980 565753 357992
rect 559920 357844 560378 357872
rect 565950 357968 566494 357992
rect 565950 357860 565966 357968
rect 566126 357860 566494 357968
rect 573590 359230 580030 359256
rect 573590 357965 573828 359230
rect 565950 357846 566494 357860
rect 573509 357959 573828 357965
rect 574685 358898 574731 358910
rect 573509 357920 573911 357959
rect 565950 357844 566418 357846
rect 559732 357540 559928 357844
rect 573509 357594 573540 357920
rect 573878 357810 573911 357920
rect 574685 357922 574691 358898
rect 574725 357922 574731 358898
rect 574685 357910 574731 357922
rect 574943 358898 574989 358910
rect 574943 357922 574949 358898
rect 574983 357922 574989 358898
rect 574943 357910 574989 357922
rect 575201 358898 575247 358910
rect 575201 357922 575207 358898
rect 575241 357922 575247 358898
rect 575201 357910 575247 357922
rect 575459 358898 575505 358910
rect 575459 357922 575465 358898
rect 575499 357922 575505 358898
rect 575459 357910 575505 357922
rect 575717 358898 575763 358910
rect 575717 357922 575723 358898
rect 575757 357922 575763 358898
rect 575717 357910 575763 357922
rect 575975 358898 576021 358910
rect 575975 357922 575981 358898
rect 576015 357922 576021 358898
rect 575975 357910 576021 357922
rect 576233 358898 576279 358910
rect 576233 357922 576239 358898
rect 576273 357922 576279 358898
rect 576233 357910 576279 357922
rect 576491 358898 576537 358910
rect 576491 357922 576497 358898
rect 576531 357922 576537 358898
rect 576491 357910 576537 357922
rect 576749 358898 576795 358910
rect 576749 357922 576755 358898
rect 576789 357922 576795 358898
rect 576749 357910 576795 357922
rect 577007 358898 577053 358910
rect 577007 357922 577013 358898
rect 577047 357922 577053 358898
rect 577007 357910 577053 357922
rect 577265 358898 577311 358910
rect 577265 357922 577271 358898
rect 577305 357922 577311 358898
rect 577265 357910 577311 357922
rect 577523 358898 577569 358910
rect 577523 357922 577529 358898
rect 577563 357922 577569 358898
rect 577523 357910 577569 357922
rect 577781 358898 577827 358910
rect 577781 357922 577787 358898
rect 577821 357922 577827 358898
rect 577781 357910 577827 357922
rect 578039 358898 578085 358910
rect 578039 357922 578045 358898
rect 578079 357922 578085 358898
rect 578039 357910 578085 357922
rect 578297 358898 578343 358910
rect 578297 357922 578303 358898
rect 578337 357922 578343 358898
rect 578297 357910 578343 357922
rect 578555 358898 578601 358910
rect 578555 357922 578561 358898
rect 578595 357922 578601 358898
rect 578555 357910 578601 357922
rect 578813 358898 578859 358910
rect 578813 357922 578819 358898
rect 578853 357922 578859 358898
rect 578813 357910 578859 357922
rect 579071 358898 579117 358910
rect 579071 357922 579077 358898
rect 579111 357922 579117 358898
rect 579071 357910 579117 357922
rect 579329 358898 579375 358910
rect 579329 357922 579335 358898
rect 579369 357922 579375 358898
rect 579329 357910 579375 357922
rect 579587 358898 579633 358910
rect 579587 357922 579593 358898
rect 579627 357922 579633 358898
rect 579587 357910 579633 357922
rect 579845 358898 579891 358910
rect 579845 357922 579851 358898
rect 579885 357922 579891 358898
rect 579845 357910 579891 357922
rect 580252 357826 580356 359786
rect 580004 357814 580356 357826
rect 573878 357682 574512 357810
rect 580004 357726 580016 357814
rect 580106 357726 580356 357814
rect 580004 357722 580356 357726
rect 580004 357720 580118 357722
rect 573878 357680 574508 357682
rect 573878 357594 574408 357680
rect 573509 357576 574408 357594
rect 574500 357576 574508 357680
rect 573509 357564 574508 357576
rect 565760 357540 566070 357542
rect 559732 357510 566070 357540
rect 559732 357450 560728 357510
rect 560788 357450 560928 357510
rect 560988 357450 561128 357510
rect 561188 357450 561328 357510
rect 561388 357450 561528 357510
rect 561588 357450 561728 357510
rect 561788 357450 561928 357510
rect 561988 357450 562128 357510
rect 562188 357450 562328 357510
rect 562388 357450 562528 357510
rect 562588 357450 562728 357510
rect 562788 357450 562928 357510
rect 562988 357450 563128 357510
rect 563188 357450 563328 357510
rect 563388 357450 563528 357510
rect 563588 357450 563728 357510
rect 563788 357450 563928 357510
rect 563988 357450 564128 357510
rect 564188 357450 564328 357510
rect 564388 357450 564528 357510
rect 564588 357450 564728 357510
rect 564788 357450 564928 357510
rect 564988 357450 565128 357510
rect 565188 357450 565328 357510
rect 565388 357450 565528 357510
rect 565588 357450 566070 357510
rect 559732 357422 566070 357450
rect 559732 357420 565856 357422
rect 565950 357230 566070 357422
rect 574644 357440 580030 357470
rect 574644 357380 574702 357440
rect 574762 357380 574902 357440
rect 574962 357380 575102 357440
rect 575162 357380 575302 357440
rect 575362 357380 575502 357440
rect 575562 357380 575702 357440
rect 575762 357380 575902 357440
rect 575962 357380 576102 357440
rect 576162 357380 576302 357440
rect 576362 357380 576502 357440
rect 576562 357380 576702 357440
rect 576762 357380 576902 357440
rect 576962 357380 577102 357440
rect 577162 357380 577302 357440
rect 577362 357380 577502 357440
rect 577562 357380 577702 357440
rect 577762 357380 577902 357440
rect 577962 357380 578102 357440
rect 578162 357380 578302 357440
rect 578362 357380 578502 357440
rect 578562 357380 578702 357440
rect 578762 357380 578902 357440
rect 578962 357380 579102 357440
rect 579162 357380 579302 357440
rect 579362 357380 579502 357440
rect 579562 357380 579702 357440
rect 579762 357380 580030 357440
rect 574644 357350 580030 357380
rect 574762 357230 574882 357350
rect 565950 357110 574882 357230
rect 508586 356418 508596 356602
rect 508732 356418 508742 356602
rect 565598 314298 573770 314418
rect 565598 313112 565718 314298
rect 560404 313082 565718 313112
rect 560404 313022 560590 313082
rect 560650 313022 560790 313082
rect 560850 313022 560990 313082
rect 561050 313022 561190 313082
rect 561250 313022 561390 313082
rect 561450 313022 561590 313082
rect 561650 313022 561790 313082
rect 561850 313022 561990 313082
rect 562050 313022 562190 313082
rect 562250 313022 562390 313082
rect 562450 313022 562590 313082
rect 562650 313022 562790 313082
rect 562850 313022 562990 313082
rect 563050 313022 563190 313082
rect 563250 313022 563390 313082
rect 563450 313022 563590 313082
rect 563650 313022 563790 313082
rect 563850 313022 563990 313082
rect 564050 313022 564190 313082
rect 564250 313022 564390 313082
rect 564450 313022 564590 313082
rect 564650 313022 564790 313082
rect 564850 313022 564990 313082
rect 565050 313022 565190 313082
rect 565250 313022 565390 313082
rect 565450 313022 565718 313082
rect 560404 312992 565718 313022
rect 566116 313610 566126 313804
rect 566346 313794 566356 313804
rect 566346 313610 566362 313794
rect 560409 312660 560455 312672
rect 559642 311536 559652 311744
rect 559860 311714 560240 311744
rect 559860 311564 560094 311714
rect 560226 311564 560240 311714
rect 560409 311684 560415 312660
rect 560449 311684 560455 312660
rect 560409 311672 560455 311684
rect 560667 312660 560713 312672
rect 560667 311684 560673 312660
rect 560707 311684 560713 312660
rect 560667 311672 560713 311684
rect 560925 312660 560971 312672
rect 560925 311684 560931 312660
rect 560965 311684 560971 312660
rect 560925 311672 560971 311684
rect 561183 312660 561229 312672
rect 561183 311684 561189 312660
rect 561223 311684 561229 312660
rect 561183 311672 561229 311684
rect 561441 312660 561487 312672
rect 561441 311684 561447 312660
rect 561481 311684 561487 312660
rect 561441 311672 561487 311684
rect 561699 312660 561745 312672
rect 561699 311684 561705 312660
rect 561739 311684 561745 312660
rect 561699 311672 561745 311684
rect 561957 312660 562003 312672
rect 561957 311684 561963 312660
rect 561997 311684 562003 312660
rect 561957 311672 562003 311684
rect 562215 312660 562261 312672
rect 562215 311684 562221 312660
rect 562255 311684 562261 312660
rect 562215 311672 562261 311684
rect 562473 312660 562519 312672
rect 562473 311684 562479 312660
rect 562513 311684 562519 312660
rect 562473 311672 562519 311684
rect 562731 312660 562777 312672
rect 562731 311684 562737 312660
rect 562771 311684 562777 312660
rect 562731 311672 562777 311684
rect 562989 312660 563035 312672
rect 562989 311684 562995 312660
rect 563029 311684 563035 312660
rect 562989 311672 563035 311684
rect 563247 312660 563293 312672
rect 563247 311684 563253 312660
rect 563287 311684 563293 312660
rect 563247 311672 563293 311684
rect 563505 312660 563551 312672
rect 563505 311684 563511 312660
rect 563545 311684 563551 312660
rect 563505 311672 563551 311684
rect 563763 312660 563809 312672
rect 563763 311684 563769 312660
rect 563803 311684 563809 312660
rect 563763 311672 563809 311684
rect 564021 312660 564067 312672
rect 564021 311684 564027 312660
rect 564061 311684 564067 312660
rect 564021 311672 564067 311684
rect 564279 312660 564325 312672
rect 564279 311684 564285 312660
rect 564319 311684 564325 312660
rect 564279 311672 564325 311684
rect 564537 312660 564583 312672
rect 564537 311684 564543 312660
rect 564577 311684 564583 312660
rect 564537 311672 564583 311684
rect 564795 312660 564841 312672
rect 564795 311684 564801 312660
rect 564835 311684 564841 312660
rect 564795 311672 564841 311684
rect 565053 312660 565099 312672
rect 565053 311684 565059 312660
rect 565093 311684 565099 312660
rect 565053 311672 565099 311684
rect 565311 312660 565357 312672
rect 565311 311684 565317 312660
rect 565351 311684 565357 312660
rect 565311 311672 565357 311684
rect 565569 312660 565615 312672
rect 565569 311684 565575 312660
rect 565609 311684 565615 312660
rect 566116 311684 566362 313610
rect 573546 313182 573770 314298
rect 580844 313778 580948 313782
rect 580756 313770 580948 313778
rect 580748 313602 580758 313770
rect 580944 313602 580954 313770
rect 573546 313152 580478 313182
rect 573546 313092 575150 313152
rect 575210 313092 575350 313152
rect 575410 313092 575550 313152
rect 575610 313092 575750 313152
rect 575810 313092 575950 313152
rect 576010 313092 576150 313152
rect 576210 313092 576350 313152
rect 576410 313092 576550 313152
rect 576610 313092 576750 313152
rect 576810 313092 576950 313152
rect 577010 313092 577150 313152
rect 577210 313092 577350 313152
rect 577410 313092 577550 313152
rect 577610 313092 577750 313152
rect 577810 313092 577950 313152
rect 578010 313092 578150 313152
rect 578210 313092 578350 313152
rect 578410 313092 578550 313152
rect 578610 313092 578750 313152
rect 578810 313092 578950 313152
rect 579010 313092 579150 313152
rect 579210 313092 579350 313152
rect 579410 313092 579550 313152
rect 579610 313092 579750 313152
rect 579810 313092 579950 313152
rect 580010 313092 580150 313152
rect 580210 313092 580478 313152
rect 573546 313062 580478 313092
rect 573546 311742 573800 313062
rect 575133 312730 575179 312742
rect 575133 311754 575139 312730
rect 575173 311754 575179 312730
rect 575133 311742 575179 311754
rect 575391 312730 575437 312742
rect 575391 311754 575397 312730
rect 575431 311754 575437 312730
rect 575391 311742 575437 311754
rect 575649 312730 575695 312742
rect 575649 311754 575655 312730
rect 575689 311754 575695 312730
rect 575649 311742 575695 311754
rect 575907 312730 575953 312742
rect 575907 311754 575913 312730
rect 575947 311754 575953 312730
rect 575907 311742 575953 311754
rect 576165 312730 576211 312742
rect 576165 311754 576171 312730
rect 576205 311754 576211 312730
rect 576165 311742 576211 311754
rect 576423 312730 576469 312742
rect 576423 311754 576429 312730
rect 576463 311754 576469 312730
rect 576423 311742 576469 311754
rect 576681 312730 576727 312742
rect 576681 311754 576687 312730
rect 576721 311754 576727 312730
rect 576681 311742 576727 311754
rect 576939 312730 576985 312742
rect 576939 311754 576945 312730
rect 576979 311754 576985 312730
rect 576939 311742 576985 311754
rect 577197 312730 577243 312742
rect 577197 311754 577203 312730
rect 577237 311754 577243 312730
rect 577197 311742 577243 311754
rect 577455 312730 577501 312742
rect 577455 311754 577461 312730
rect 577495 311754 577501 312730
rect 577455 311742 577501 311754
rect 577713 312730 577759 312742
rect 577713 311754 577719 312730
rect 577753 311754 577759 312730
rect 577713 311742 577759 311754
rect 577971 312730 578017 312742
rect 577971 311754 577977 312730
rect 578011 311754 578017 312730
rect 577971 311742 578017 311754
rect 578229 312730 578275 312742
rect 578229 311754 578235 312730
rect 578269 311754 578275 312730
rect 578229 311742 578275 311754
rect 578487 312730 578533 312742
rect 578487 311754 578493 312730
rect 578527 311754 578533 312730
rect 578487 311742 578533 311754
rect 578745 312730 578791 312742
rect 578745 311754 578751 312730
rect 578785 311754 578791 312730
rect 578745 311742 578791 311754
rect 579003 312730 579049 312742
rect 579003 311754 579009 312730
rect 579043 311754 579049 312730
rect 579003 311742 579049 311754
rect 579261 312730 579307 312742
rect 579261 311754 579267 312730
rect 579301 311754 579307 312730
rect 579261 311742 579307 311754
rect 579519 312730 579565 312742
rect 579519 311754 579525 312730
rect 579559 311754 579565 312730
rect 579519 311742 579565 311754
rect 579777 312730 579823 312742
rect 579777 311754 579783 312730
rect 579817 311754 579823 312730
rect 579777 311742 579823 311754
rect 580035 312730 580081 312742
rect 580035 311754 580041 312730
rect 580075 311754 580081 312730
rect 580035 311742 580081 311754
rect 580293 312730 580339 312742
rect 580293 311754 580299 312730
rect 580333 311754 580339 312730
rect 580293 311742 580339 311754
rect 565569 311672 565615 311684
rect 559860 311536 560240 311564
rect 565812 311660 566362 311684
rect 565812 311552 565828 311660
rect 565988 311552 566362 311660
rect 565812 311536 566362 311552
rect 573432 311700 574046 311742
rect 559648 311232 559880 311536
rect 573432 311420 573492 311700
rect 573834 311590 574046 311700
rect 580756 311658 580948 313602
rect 580452 311646 580948 311658
rect 573834 311524 574952 311590
rect 580452 311558 580464 311646
rect 580554 311558 580948 311646
rect 580452 311554 580948 311558
rect 580452 311552 580566 311554
rect 573834 311512 574956 311524
rect 573834 311420 574856 311512
rect 573432 311408 574856 311420
rect 574948 311408 574956 311512
rect 573432 311396 574956 311408
rect 573432 311392 574952 311396
rect 573432 311382 574050 311392
rect 575092 311272 580478 311302
rect 559648 311202 565718 311232
rect 559648 311142 560590 311202
rect 560650 311142 560790 311202
rect 560850 311142 560990 311202
rect 561050 311142 561190 311202
rect 561250 311142 561390 311202
rect 561450 311142 561590 311202
rect 561650 311142 561790 311202
rect 561850 311142 561990 311202
rect 562050 311142 562190 311202
rect 562250 311142 562390 311202
rect 562450 311142 562590 311202
rect 562650 311142 562790 311202
rect 562850 311142 562990 311202
rect 563050 311142 563190 311202
rect 563250 311142 563390 311202
rect 563450 311142 563590 311202
rect 563650 311142 563790 311202
rect 563850 311142 563990 311202
rect 564050 311142 564190 311202
rect 564250 311142 564390 311202
rect 564450 311142 564590 311202
rect 564650 311142 564790 311202
rect 564850 311142 564990 311202
rect 565050 311142 565190 311202
rect 565250 311142 565390 311202
rect 565450 311172 565718 311202
rect 575092 311212 575150 311272
rect 575210 311212 575350 311272
rect 575410 311212 575550 311272
rect 575610 311212 575750 311272
rect 575810 311212 575950 311272
rect 576010 311212 576150 311272
rect 576210 311212 576350 311272
rect 576410 311212 576550 311272
rect 576610 311212 576750 311272
rect 576810 311212 576950 311272
rect 577010 311212 577150 311272
rect 577210 311212 577350 311272
rect 577410 311212 577550 311272
rect 577610 311212 577750 311272
rect 577810 311212 577950 311272
rect 578010 311212 578150 311272
rect 578210 311212 578350 311272
rect 578410 311212 578550 311272
rect 578610 311212 578750 311272
rect 578810 311212 578950 311272
rect 579010 311212 579150 311272
rect 579210 311212 579350 311272
rect 579410 311212 579550 311272
rect 579610 311212 579750 311272
rect 579810 311212 579950 311272
rect 580010 311212 580150 311272
rect 580210 311212 580478 311272
rect 575092 311182 580478 311212
rect 575092 311172 575350 311182
rect 565450 311142 575350 311172
rect 559648 311052 575350 311142
<< via1 >>
rect 566186 494126 566408 494310
rect 559802 492324 560012 492536
rect 580856 494136 581040 494348
rect 573564 491888 573874 492160
rect 566256 405258 566462 405476
rect 559736 403192 559926 403368
rect 580074 405292 580182 405402
rect 573538 402980 573888 403312
rect 566274 359786 566500 359978
rect 559712 357844 559920 358052
rect 580252 359786 580358 359906
rect 573540 357594 573878 357920
rect 508596 356418 508732 356602
rect 566126 313610 566346 313804
rect 559652 311536 559860 311744
rect 580758 313602 580944 313770
rect 573492 311420 573834 311700
<< metal2 >>
rect 580856 494348 581040 494358
rect 566186 494310 566408 494320
rect 580856 494126 581040 494136
rect 566186 494116 566408 494126
rect 559802 492536 560012 492546
rect 559802 492314 560012 492324
rect 573564 492160 573874 492170
rect 573564 491878 573874 491888
rect 566256 405476 566462 405486
rect 580074 405402 580182 405412
rect 580074 405282 580182 405292
rect 566256 405248 566462 405258
rect 559736 403368 559926 403378
rect 559736 403182 559926 403192
rect 573538 403312 573888 403322
rect 573538 402970 573888 402980
rect 541964 389510 542078 389520
rect 541964 389424 542078 389434
rect 541958 380668 542080 380678
rect 541958 380514 542080 380524
rect 566274 359978 566500 359988
rect 566274 359776 566500 359786
rect 580252 359906 580358 359916
rect 580252 359776 580358 359786
rect 559712 358052 559920 358062
rect 559712 357834 559920 357844
rect 573540 357920 573878 357930
rect 573540 357584 573878 357594
rect 508596 356602 508732 356612
rect 508596 356408 508732 356418
rect 566126 313804 566346 313814
rect 566126 313600 566346 313610
rect 580758 313770 580944 313780
rect 580758 313592 580944 313602
rect 559652 311744 559860 311754
rect 559652 311526 559860 311536
rect 573492 311700 573834 311710
rect 573492 311410 573834 311420
<< via2 >>
rect 566186 494126 566408 494310
rect 580856 494136 581040 494348
rect 559802 492324 560012 492536
rect 573564 491888 573874 492160
rect 566256 405258 566462 405476
rect 580074 405292 580182 405402
rect 559736 403192 559926 403368
rect 573538 402980 573888 403312
rect 541964 389434 542078 389510
rect 541958 380524 542080 380668
rect 566274 359786 566500 359978
rect 580252 359786 580358 359906
rect 559712 357844 559920 358052
rect 573540 357594 573878 357920
rect 508596 356418 508732 356602
rect 566126 313610 566346 313804
rect 580758 313602 580944 313770
rect 559652 311536 559860 311744
rect 573492 311420 573834 311700
<< metal3 >>
rect 413300 698232 418436 703282
rect 465296 698476 470432 703526
rect 510560 701276 515394 703604
rect 510552 701180 515394 701276
rect 510552 700092 515386 701180
rect 510552 699264 515392 700092
rect 510538 697668 515392 699264
rect 510538 697378 515372 697668
rect 510538 696840 510704 697378
rect 510560 689882 510704 696840
rect 515202 689882 515372 697378
rect 510560 689666 515372 689882
rect 520554 697354 525388 703122
rect 566500 698354 571636 703404
rect 520554 689858 520704 697354
rect 525202 689858 525388 697354
rect 520554 689727 525388 689858
rect 577256 677954 582392 683004
rect 567105 644596 581232 644606
rect 567105 644324 582918 644596
rect 567105 640080 567306 644324
rect 573722 640080 582918 644324
rect 567105 639760 582918 640080
rect 567308 634256 583176 634588
rect 567296 630012 567306 634256
rect 573722 630012 583176 634256
rect 567308 629752 583176 630012
rect 580846 494348 581050 494353
rect 566148 494310 566454 494332
rect 566148 494248 566186 494310
rect 501828 494126 566186 494248
rect 566408 494248 566454 494310
rect 580846 494248 580856 494348
rect 566408 494136 580856 494248
rect 581040 494248 581050 494348
rect 581040 494136 583862 494248
rect 566408 494126 583862 494136
rect 501828 494124 583862 494126
rect 501828 414988 501952 494124
rect 566148 494090 566454 494124
rect 559792 492536 560022 492541
rect 559792 492324 559802 492536
rect 560012 492324 560022 492536
rect 559792 492319 560022 492324
rect 573554 492160 573884 492165
rect 573554 491888 573564 492160
rect 573874 491888 573884 492160
rect 573554 491883 573884 491888
rect 501002 414864 501952 414988
rect 501002 414800 501126 414864
rect 566246 405476 566472 405481
rect 566246 405400 566256 405476
rect 542686 405288 566256 405400
rect 542686 389534 542798 405288
rect 566246 405258 566256 405288
rect 566462 405400 566472 405476
rect 580064 405402 580192 405407
rect 580064 405400 580074 405402
rect 566462 405292 580074 405400
rect 580182 405400 580192 405402
rect 580182 405292 583872 405400
rect 566462 405288 583872 405292
rect 566462 405258 566472 405288
rect 580064 405287 580192 405288
rect 566246 405253 566472 405258
rect 559726 403368 559936 403373
rect 559726 403192 559736 403368
rect 559926 403192 559936 403368
rect 559726 403187 559936 403192
rect 573528 403312 573898 403317
rect 573528 402980 573538 403312
rect 573888 402980 573898 403312
rect 573528 402975 573898 402980
rect 541954 389510 542798 389534
rect 541954 389434 541964 389510
rect 542078 389434 542798 389510
rect 541954 389422 542798 389434
rect 541943 380668 545137 380703
rect 541943 380524 541958 380668
rect 542080 380615 545137 380668
rect 542080 380524 545141 380615
rect 541943 380497 545141 380524
rect 545023 359903 545141 380497
rect 566264 359978 566510 359983
rect 566264 359903 566274 359978
rect 545023 359786 566274 359903
rect 566500 359903 566510 359978
rect 580242 359906 580368 359911
rect 580242 359903 580252 359906
rect 566500 359786 580252 359903
rect 580358 359903 580368 359906
rect 580358 359786 580941 359903
rect 545023 359785 580941 359786
rect 566264 359781 566510 359785
rect 580242 359781 580368 359785
rect 580823 358984 580941 359785
rect 580823 358866 583840 358984
rect 580823 358859 580941 358866
rect 559702 358052 559930 358057
rect 559702 357844 559712 358052
rect 559920 357844 559930 358052
rect 559702 357839 559930 357844
rect 573530 357920 573888 357925
rect 573530 357594 573540 357920
rect 573878 357594 573888 357920
rect 573530 357589 573888 357594
rect 508585 356602 509603 356611
rect 508585 356418 508596 356602
rect 508732 356418 509603 356602
rect 508585 356401 509603 356418
rect 509393 313770 509603 356401
rect 566116 313804 566356 313809
rect 566116 313770 566126 313804
rect 509393 313610 566126 313770
rect 566346 313770 566356 313804
rect 580748 313770 580954 313775
rect 566346 313610 580758 313770
rect 509393 313602 580758 313610
rect 580944 313727 583738 313770
rect 580944 313602 583873 313727
rect 509393 313593 583873 313602
rect 559642 311744 559870 311749
rect 559642 311536 559652 311744
rect 559860 311536 559870 311744
rect 559642 311531 559870 311536
rect 573482 311700 573844 311705
rect 573482 311420 573492 311700
rect 573834 311420 573844 311700
rect 573482 311415 573844 311420
<< via3 >>
rect 510704 689882 515202 697378
rect 520704 689858 525202 697354
rect 567306 640080 573722 644324
rect 567306 630012 573722 634256
rect 559802 492324 560012 492536
rect 573564 491888 573874 492160
rect 559736 403192 559926 403368
rect 573538 402980 573888 403312
rect 559712 357844 559920 358052
rect 573540 357594 573878 357920
rect 559652 311536 559860 311744
rect 573492 311420 573834 311700
<< metal4 >>
rect 502376 697378 560022 697790
rect 502376 689882 510704 697378
rect 515202 697354 560022 697378
rect 515202 689882 520704 697354
rect 502376 689858 520704 689882
rect 525202 689858 560022 697354
rect 502376 689742 560022 689858
rect 551974 492536 560022 689742
rect 567305 644324 573723 644325
rect 567305 640080 567306 644324
rect 573722 640080 573723 644324
rect 567305 640079 573723 640080
rect 567305 634256 573723 634257
rect 567305 630012 567306 634256
rect 573722 630012 573723 634256
rect 567305 630011 573723 630012
rect 551974 492324 559802 492536
rect 560012 492324 560022 492536
rect 551974 414054 560022 492324
rect 573563 492160 573875 492161
rect 573563 491888 573564 492160
rect 573874 491888 573875 492160
rect 573563 491887 573875 491888
rect 540412 412422 560022 414054
rect 551974 403368 560022 412422
rect 551974 403192 559736 403368
rect 559926 403192 560022 403368
rect 551974 359050 560022 403192
rect 573537 403312 573889 403313
rect 573537 402980 573538 403312
rect 573888 402980 573889 403312
rect 573537 402979 573889 402980
rect 534818 358052 560022 359050
rect 534818 357844 559712 358052
rect 559920 357844 560022 358052
rect 534818 357418 560022 357844
rect 573539 357920 573879 357921
rect 573539 357594 573540 357920
rect 573878 357594 573879 357920
rect 573539 357593 573879 357594
rect 551974 311744 560022 357418
rect 551974 311536 559652 311744
rect 559860 311536 560022 311744
rect 551974 154934 560022 311536
rect 573491 311700 573835 311701
rect 573491 311420 573492 311700
rect 573834 311420 573835 311700
rect 573491 311419 573835 311420
<< via4 >>
rect 567306 640080 573722 644324
rect 567306 630012 573722 634256
rect 573564 491888 573874 492160
rect 573538 402980 573888 403312
rect 573540 357594 573878 357920
rect 573492 311420 573834 311700
<< metal5 >>
rect 567158 644324 573920 649062
rect 567158 640080 567306 644324
rect 573722 640080 573920 644324
rect 567158 634256 573920 640080
rect 567158 630012 567306 634256
rect 573722 630012 573920 634256
rect 567158 627314 573920 630012
rect 567156 621952 573942 627314
rect 567158 492160 573920 621952
rect 567158 491888 573564 492160
rect 573874 491888 573920 492160
rect 488780 422974 490412 423442
rect 567158 422974 573920 491888
rect 488780 421342 573920 422974
rect 488780 411206 490412 421342
rect 536984 420968 573920 421342
rect 537164 413148 538796 420968
rect 567158 403312 573920 420968
rect 567158 402980 573538 403312
rect 573888 402980 573920 403312
rect 488780 348924 490412 358644
rect 537164 348924 538796 359482
rect 567158 357920 573920 402980
rect 567158 357594 573540 357920
rect 573878 357594 573920 357920
rect 567158 348924 573920 357594
rect 488668 347292 573920 348924
rect 567158 311700 573920 347292
rect 567158 311420 573492 311700
rect 573834 311420 573920 311700
rect 567158 147385 573920 311420
use bgr_final  bgr_final_0
timestamp 1654904630
transform 0 -1 542076 -1 0 414984
box 0 0 58512 56576
<< labels >>
flabel metal3 510596 697782 515352 701406 1 FreeSans 8000 0 0 0 VSSA1
flabel metal3 574704 639800 581232 644606 1 FreeSans 8000 0 0 0 VCCD1
flabel metal1 565560 313022 565620 313082 1 FreeSans 800 0 0 0 nmos_flat_3/VPWR
flabel metal1 565560 311142 565620 311202 1 FreeSans 800 0 0 0 nmos_flat_3/VGND
flabel locali 560404 312862 560464 312922 1 FreeSans 800 0 0 0 nmos_flat_3/SOURCE
flabel locali 560404 311542 560464 311602 1 FreeSans 800 0 0 0 nmos_flat_3/DRAIN
flabel locali 560404 311376 560464 311436 1 FreeSans 800 0 0 0 nmos_flat_3/GATE
flabel nwell 580418 313092 580478 313152 1 FreeSans 800 0 0 0 pmos_flat_2/VPWR
flabel metal1 580320 311212 580478 311272 1 FreeSans 800 0 0 0 pmos_flat_2/VGND
flabel locali 575092 312932 575152 312972 1 FreeSans 800 0 0 0 pmos_flat_2/SOURCE
flabel locali 575092 311552 575152 311612 1 FreeSans 800 0 0 0 pmos_flat_2/DRAIN
flabel locali 575092 311390 575152 311450 1 FreeSans 800 0 0 0 pmos_flat_2/GATE
flabel metal1 565806 493790 565866 493850 1 FreeSans 800 0 0 0 nmos_flat_0/VPWR
flabel metal1 565806 491910 565866 491970 1 FreeSans 800 0 0 0 nmos_flat_0/VGND
flabel locali 560650 493630 560710 493690 1 FreeSans 800 0 0 0 nmos_flat_0/SOURCE
flabel locali 560650 492310 560710 492370 1 FreeSans 800 0 0 0 nmos_flat_0/DRAIN
flabel locali 560650 492144 560710 492204 1 FreeSans 800 0 0 0 nmos_flat_0/GATE
flabel metal1 565742 404648 565802 404708 1 FreeSans 800 0 0 0 nmos_flat_1/VPWR
flabel metal1 565742 402768 565802 402828 1 FreeSans 800 0 0 0 nmos_flat_1/VGND
flabel locali 560586 404488 560646 404548 1 FreeSans 800 0 0 0 nmos_flat_1/SOURCE
flabel locali 560586 403168 560646 403228 1 FreeSans 800 0 0 0 nmos_flat_1/DRAIN
flabel locali 560586 403002 560646 403062 1 FreeSans 800 0 0 0 nmos_flat_1/GATE
flabel metal1 565698 359330 565758 359390 1 FreeSans 800 0 0 0 nmos_flat_2/VPWR
flabel metal1 565698 357450 565758 357510 1 FreeSans 800 0 0 0 nmos_flat_2/VGND
flabel locali 560542 359170 560602 359230 1 FreeSans 800 0 0 0 nmos_flat_2/SOURCE
flabel locali 560542 357850 560602 357910 1 FreeSans 800 0 0 0 nmos_flat_2/DRAIN
flabel locali 560542 357684 560602 357744 1 FreeSans 800 0 0 0 nmos_flat_2/GATE
flabel nwell 579774 404688 579834 404748 1 FreeSans 800 0 0 0 pmos_flat_0/VPWR
flabel metal1 579676 402808 579834 402868 1 FreeSans 800 0 0 0 pmos_flat_0/VGND
flabel locali 574448 404528 574508 404568 1 FreeSans 800 0 0 0 pmos_flat_0/SOURCE
flabel locali 574448 403148 574508 403208 1 FreeSans 800 0 0 0 pmos_flat_0/DRAIN
flabel locali 574448 402986 574508 403046 1 FreeSans 800 0 0 0 pmos_flat_0/GATE
flabel nwell 579970 359260 580030 359320 1 FreeSans 800 0 0 0 pmos_flat_1/VPWR
flabel metal1 579872 357380 580030 357440 1 FreeSans 800 0 0 0 pmos_flat_1/VGND
flabel locali 574644 359100 574704 359140 1 FreeSans 800 0 0 0 pmos_flat_1/SOURCE
flabel locali 574644 357720 574704 357780 1 FreeSans 800 0 0 0 pmos_flat_1/DRAIN
flabel locali 574644 357558 574704 357618 1 FreeSans 800 0 0 0 pmos_flat_1/GATE
flabel nwell 580496 493564 580556 493624 1 FreeSans 800 0 0 0 pmos_flat_3/VPWR
flabel metal1 580398 491684 580556 491744 1 FreeSans 800 0 0 0 pmos_flat_3/VGND
flabel locali 575170 493404 575230 493444 1 FreeSans 800 0 0 0 pmos_flat_3/SOURCE
flabel locali 575170 492024 575230 492084 1 FreeSans 800 0 0 0 pmos_flat_3/DRAIN
flabel locali 575170 491862 575230 491922 1 FreeSans 800 0 0 0 pmos_flat_3/GATE
<< end >>
