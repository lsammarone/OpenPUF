magic
tech sky130A
magscale 1 2
timestamp 1656715967
<< error_p >>
rect -309 142 309 178
<< metal4 >>
rect -309 118 309 142
rect -309 -118 -278 118
rect -42 -118 42 118
rect 278 -118 309 118
rect -309 -142 309 -118
<< via4 >>
rect -278 -118 -42 118
rect 42 -118 278 118
<< metal5 >>
rect -309 118 309 142
rect -309 -118 -278 118
rect -42 -118 42 118
rect 278 -118 309 118
rect -309 -142 309 -118
<< properties >>
string GDS_END 9319710
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/design_merged.gds
string GDS_START 9319450
<< end >>
