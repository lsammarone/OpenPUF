magic
tech sky130A
magscale 1 2
timestamp 1654736712
<< nwell >>
rect 2282 4742 3458 4844
rect 4170 4722 5346 4824
rect 17380 4740 18556 4842
rect 19268 4740 20444 4842
<< locali >>
rect 4626 5009 4668 5012
rect 2742 5005 2784 5008
rect 2742 4971 2746 5005
rect 2780 4971 2784 5005
rect 2742 4968 2784 4971
rect 4626 4975 4630 5009
rect 4664 4975 4668 5009
rect 19724 5009 19766 5012
rect 4626 4972 4668 4975
rect 17840 5005 17882 5008
rect 17840 4971 17844 5005
rect 17878 4971 17882 5005
rect 19724 4975 19728 5009
rect 19762 4975 19766 5009
rect 19724 4972 19766 4975
rect 17840 4968 17882 4971
<< viali >>
rect 2552 5144 2586 5178
rect 2700 5144 2734 5178
rect 2848 5144 2882 5178
rect 2996 5144 3030 5178
rect 4222 5142 4256 5176
rect 4370 5142 4404 5176
rect 4518 5142 4552 5176
rect 4666 5142 4700 5176
rect 17606 5144 17640 5178
rect 17738 5144 17772 5178
rect 17870 5144 17904 5178
rect 18002 5144 18036 5178
rect 19232 5142 19266 5176
rect 19364 5142 19398 5176
rect 19496 5142 19530 5176
rect 19628 5142 19662 5176
rect 2245 4973 2279 5007
rect 2411 4971 2445 5005
rect 2575 4969 2609 5003
rect 2746 4971 2780 5005
rect 2915 4967 2949 5001
rect 3084 4966 3118 5000
rect 3250 4972 3284 5006
rect 3420 4974 3454 5008
rect 4134 4971 4168 5005
rect 4294 4971 4328 5005
rect 4461 4965 4495 4999
rect 4630 4975 4664 5009
rect 4794 4962 4828 4996
rect 4964 4968 4998 5002
rect 5134 4970 5168 5004
rect 5293 4972 5327 5006
rect 17678 4970 17712 5004
rect 17844 4971 17878 5005
rect 18014 4972 18048 5006
rect 18180 4974 18214 5008
rect 19564 4972 19598 5006
rect 19728 4975 19762 5009
rect 19898 4970 19932 5004
rect 20060 4972 20094 5006
<< metal1 >>
rect 3494 5350 4022 5448
rect 18642 5350 19124 5448
rect 2482 5178 4934 5194
rect 2482 5144 2552 5178
rect 2586 5144 2700 5178
rect 2734 5144 2848 5178
rect 2882 5144 2996 5178
rect 3030 5176 4934 5178
rect 3030 5144 4222 5176
rect 2482 5142 4222 5144
rect 4256 5142 4370 5176
rect 4404 5142 4518 5176
rect 4552 5142 4666 5176
rect 4700 5142 4934 5176
rect 2482 5126 4934 5142
rect 17530 5178 19912 5190
rect 17530 5144 17606 5178
rect 17640 5144 17738 5178
rect 17772 5144 17870 5178
rect 17904 5144 18002 5178
rect 18036 5176 19912 5178
rect 18036 5144 19232 5176
rect 17530 5142 19232 5144
rect 19266 5142 19364 5176
rect 19398 5142 19496 5176
rect 19530 5142 19628 5176
rect 19662 5142 19912 5176
rect 17530 5128 19912 5142
rect 2230 5008 3467 5020
rect 17520 5018 18342 5038
rect 2230 5007 3420 5008
rect 2230 4973 2245 5007
rect 2279 5006 3420 5007
rect 2279 5005 3250 5006
rect 2279 5002 2411 5005
rect 2445 5004 2746 5005
rect 2780 5004 3250 5005
rect 2445 5003 2740 5004
rect 2445 5002 2575 5003
rect 2279 4973 2282 5002
rect 2230 4950 2282 4973
rect 2334 4950 2389 5002
rect 2445 4971 2495 5002
rect 2441 4950 2495 4971
rect 2547 4969 2575 5002
rect 2609 5002 2740 5003
rect 2609 4969 2611 5002
rect 2547 4950 2611 4969
rect 2663 4952 2740 5002
rect 2792 5003 3250 5004
rect 3284 5003 3420 5006
rect 2792 4952 2874 5003
rect 2926 5001 2991 5003
rect 2949 4967 2991 5001
rect 2663 4951 2874 4952
rect 2926 4951 2991 4967
rect 3043 5000 3096 5003
rect 3043 4966 3084 5000
rect 3043 4951 3096 4966
rect 3148 4951 3202 5003
rect 3284 4972 3299 5003
rect 3254 4951 3299 4972
rect 3351 4951 3396 5003
rect 3454 4974 3467 5008
rect 3448 4951 3467 4974
rect 2663 4950 3467 4951
rect 2230 4936 3467 4950
rect 4120 5009 5346 5018
rect 4120 5005 4630 5009
rect 4120 4971 4134 5005
rect 4168 4999 4294 5005
rect 4328 4999 4630 5005
rect 4168 4971 4171 4999
rect 4120 4947 4171 4971
rect 4223 4947 4278 4999
rect 4330 4947 4384 4999
rect 4436 4965 4461 4999
rect 4495 4965 4500 4999
rect 4436 4947 4500 4965
rect 4552 4975 4630 4999
rect 4664 5006 5346 5009
rect 4664 5004 5293 5006
rect 4664 5002 5134 5004
rect 4664 5000 4964 5002
rect 4998 5000 5134 5002
rect 5168 5000 5293 5004
rect 5327 5000 5346 5006
rect 4664 4975 4763 5000
rect 4815 4996 4880 5000
rect 4552 4948 4763 4975
rect 4828 4962 4880 4996
rect 4815 4948 4880 4962
rect 4932 4968 4964 5000
rect 4932 4948 4985 4968
rect 5037 4948 5091 5000
rect 5168 4970 5188 5000
rect 5143 4948 5188 4970
rect 5240 4948 5285 5000
rect 5337 4948 5346 5000
rect 4552 4947 5346 4948
rect 4120 4934 5346 4947
rect 17520 5016 18160 5018
rect 17520 4964 17668 5016
rect 17720 5005 18006 5016
rect 17720 5004 17844 5005
rect 17878 5004 18006 5005
rect 17720 4964 17838 5004
rect 17520 4952 17838 4964
rect 17890 4964 18006 5004
rect 18058 4966 18160 5016
rect 18212 5008 18342 5018
rect 18214 4974 18342 5008
rect 18212 4966 18342 4974
rect 18058 4964 18342 4966
rect 17890 4952 18342 4964
rect 17520 4936 18342 4952
rect 19522 5009 20140 5022
rect 19522 5006 19728 5009
rect 19522 4972 19564 5006
rect 19598 5002 19728 5006
rect 19762 5006 20140 5009
rect 19762 5004 20060 5006
rect 19762 5002 19898 5004
rect 19932 5002 20060 5004
rect 19522 4950 19570 4972
rect 19622 4950 19720 5002
rect 19772 4950 19850 5002
rect 19932 4970 19996 5002
rect 19902 4950 19996 4970
rect 20048 4972 20060 5002
rect 20094 4972 20140 5006
rect 20048 4950 20140 4972
rect 19522 4932 20140 4950
<< via1 >>
rect 2282 4950 2334 5002
rect 2389 4971 2411 5002
rect 2411 4971 2441 5002
rect 2389 4950 2441 4971
rect 2495 4950 2547 5002
rect 2611 4950 2663 5002
rect 2740 4971 2746 5004
rect 2746 4971 2780 5004
rect 2780 4971 2792 5004
rect 2740 4952 2792 4971
rect 2874 5001 2926 5003
rect 2874 4967 2915 5001
rect 2915 4967 2926 5001
rect 2874 4951 2926 4967
rect 2991 4951 3043 5003
rect 3096 5000 3148 5003
rect 3096 4966 3118 5000
rect 3118 4966 3148 5000
rect 3096 4951 3148 4966
rect 3202 4972 3250 5003
rect 3250 4972 3254 5003
rect 3202 4951 3254 4972
rect 3299 4951 3351 5003
rect 3396 4974 3420 5003
rect 3420 4974 3448 5003
rect 3396 4951 3448 4974
rect 4171 4947 4223 4999
rect 4278 4971 4294 4999
rect 4294 4971 4328 4999
rect 4328 4971 4330 4999
rect 4278 4947 4330 4971
rect 4384 4947 4436 4999
rect 4500 4947 4552 4999
rect 4763 4996 4815 5000
rect 4763 4962 4794 4996
rect 4794 4962 4815 4996
rect 4763 4948 4815 4962
rect 4880 4948 4932 5000
rect 4985 4968 4998 5000
rect 4998 4968 5037 5000
rect 4985 4948 5037 4968
rect 5091 4970 5134 5000
rect 5134 4970 5143 5000
rect 5091 4948 5143 4970
rect 5188 4948 5240 5000
rect 5285 4972 5293 5000
rect 5293 4972 5327 5000
rect 5327 4972 5337 5000
rect 5285 4948 5337 4972
rect 17668 5004 17720 5016
rect 18006 5006 18058 5016
rect 17668 4970 17678 5004
rect 17678 4970 17712 5004
rect 17712 4970 17720 5004
rect 17668 4964 17720 4970
rect 17838 4971 17844 5004
rect 17844 4971 17878 5004
rect 17878 4971 17890 5004
rect 17838 4952 17890 4971
rect 18006 4972 18014 5006
rect 18014 4972 18048 5006
rect 18048 4972 18058 5006
rect 18006 4964 18058 4972
rect 18160 5008 18212 5018
rect 18160 4974 18180 5008
rect 18180 4974 18212 5008
rect 18160 4966 18212 4974
rect 19570 4972 19598 5002
rect 19598 4972 19622 5002
rect 19570 4950 19622 4972
rect 19720 4975 19728 5002
rect 19728 4975 19762 5002
rect 19762 4975 19772 5002
rect 19720 4950 19772 4975
rect 19850 4970 19898 5002
rect 19898 4970 19902 5002
rect 19850 4950 19902 4970
rect 19996 4950 20048 5002
<< metal2 >>
rect -1439 5082 -413 5083
rect 446 5082 1472 5084
rect 13643 5082 14669 5084
rect 15544 5082 16570 5083
rect 21211 5082 22237 5086
rect 23115 5082 24141 5083
rect -1666 5004 11208 5082
rect 11562 5020 26308 5082
rect -1666 5002 2740 5004
rect -1666 4950 2282 5002
rect 2334 4950 2389 5002
rect 2441 4950 2495 5002
rect 2547 4950 2611 5002
rect 2663 4952 2740 5002
rect 2792 5003 11208 5004
rect 2792 4952 2874 5003
rect 2663 4951 2874 4952
rect 2926 4951 2991 5003
rect 3043 4951 3096 5003
rect 3148 4951 3202 5003
rect 3254 4951 3299 5003
rect 3351 4951 3396 5003
rect 3448 5000 11208 5003
rect 3448 4999 4763 5000
rect 3448 4951 4171 4999
rect 2663 4950 4171 4951
rect -1666 4947 4171 4950
rect 4223 4947 4278 4999
rect 4330 4947 4384 4999
rect 4436 4947 4500 4999
rect 4552 4948 4763 4999
rect 4815 4948 4880 5000
rect 4932 4948 4985 5000
rect 5037 4948 5091 5000
rect 5143 4948 5188 5000
rect 5240 4948 5285 5000
rect 5337 4948 11208 5000
rect 11563 5018 26308 5020
rect 11563 5016 18160 5018
rect 11563 4964 17668 5016
rect 17720 5004 18006 5016
rect 17720 4964 17838 5004
rect 11563 4956 17838 4964
rect 4552 4947 11208 4948
rect -1666 4894 11208 4947
rect 11562 4952 17838 4956
rect 17890 4964 18006 5004
rect 18058 4966 18160 5016
rect 18212 5002 26308 5018
rect 18212 4966 19570 5002
rect 18058 4964 19570 4966
rect 17890 4952 19570 4964
rect 11562 4950 19570 4952
rect 19622 4950 19720 5002
rect 19772 4950 19850 5002
rect 19902 4950 19996 5002
rect 20048 4950 26308 5002
rect 11562 4894 26308 4950
rect -1439 4637 -413 4894
rect 446 4637 1472 4894
rect 2150 4886 5358 4894
rect 2150 4637 3470 4886
rect -1666 4590 3470 4637
rect 4034 4633 5358 4886
rect 6115 4633 7141 4894
rect 8010 4633 9036 4894
rect 9879 4633 10905 4894
rect 11756 4637 12782 4894
rect 13643 4637 14669 4894
rect 15544 4637 16570 4894
rect 17248 4886 20456 4894
rect 17248 4637 18568 4886
rect 19132 4637 20456 4886
rect 21211 4637 22237 4894
rect 23115 4637 24141 4894
rect 24991 4637 26017 4894
rect 4034 4590 11208 4633
rect -1666 4528 11208 4590
rect 11562 4590 26307 4637
rect 11562 4528 26306 4590
rect 2150 4524 3470 4528
rect 4034 4524 11208 4528
rect 17248 4524 18568 4528
rect 19132 4524 20456 4528
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0
timestamp 1654736712
transform 1 0 19092 0 -1 5398
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1654736712
transform 1 0 17210 0 -1 5400
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_2
timestamp 1654736712
transform 1 0 3994 0 -1 5398
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_3
timestamp 1654736712
transform 1 0 2112 0 -1 5400
box -38 -48 1510 592
use unitcell2buf_32  unitcell2buf_32_0
timestamp 1654736712
transform 1 0 23448 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf_32  unitcell2buf_32_1
timestamp 1654736712
transform 1 0 21560 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf_32  unitcell2buf_32_2
timestamp 1654736712
transform 1 0 19672 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf_32  unitcell2buf_32_3
timestamp 1654736712
transform 1 0 17784 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf_32  unitcell2buf_32_4
timestamp 1654736712
transform 1 0 15896 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf_32  unitcell2buf_32_5
timestamp 1654736712
transform 1 0 14008 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf_32  unitcell2buf_32_6
timestamp 1654736712
transform 1 0 12120 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf_32  unitcell2buf_32_7
timestamp 1654736712
transform 1 0 8350 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf_32  unitcell2buf_32_8
timestamp 1654736712
transform 1 0 6462 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf_32  unitcell2buf_32_9
timestamp 1654736712
transform 1 0 4574 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf_32  unitcell2buf_32_10
timestamp 1654736712
transform 1 0 2686 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf_32  unitcell2buf_32_11
timestamp 1654736712
transform 1 0 -1090 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf_32  unitcell2buf_32_12
timestamp 1654736712
transform 1 0 798 0 1 3712
box -574 -1185 1322 1192
use unitcell2bufcut_32  unitcell2bufcut_32_0
timestamp 1654736712
transform 1 0 25336 0 1 3712
box -574 -1185 1322 1192
use unitcell2bufcut_32  unitcell2bufcut_32_1
timestamp 1654736712
transform 1 0 10238 0 1 3712
box -574 -1185 1322 1192
<< end >>
