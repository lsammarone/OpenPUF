magic
tech sky130A
timestamp 1654736712
<< metal2 >>
rect -109 14 109 24
rect -109 -14 -94 14
rect -66 -14 -54 14
rect -26 -14 -14 14
rect 14 -14 26 14
rect 54 -14 66 14
rect 94 -14 109 14
rect -109 -24 109 -14
<< via2 >>
rect -94 -14 -66 14
rect -54 -14 -26 14
rect -14 -14 14 14
rect 26 -14 54 14
rect 66 -14 94 14
<< metal3 >>
rect -109 14 109 24
rect -109 -14 -94 14
rect -66 -14 -54 14
rect -26 -14 -14 14
rect 14 -14 26 14
rect 54 -14 66 14
rect 94 -14 109 14
rect -109 -24 109 -14
<< end >>
