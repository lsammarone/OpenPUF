magic
tech sky130A
magscale 1 2
timestamp 1656715967
<< metal1 >>
rect 33068 17224 39642 17354
rect 33068 16746 33440 17224
rect 33818 16746 39642 17224
rect 33068 16634 39642 16746
rect 40740 17264 132484 17370
rect 40740 16750 131206 17264
rect 131660 16750 132484 17264
rect 40740 16650 132484 16750
rect 36596 10800 43067 10858
rect 36596 10086 36762 10800
rect 37016 10086 43067 10800
rect 36596 10036 43067 10086
rect 44147 10758 128739 10874
rect 44147 10114 127624 10758
rect 128126 10114 128739 10758
rect 44147 10052 128739 10114
<< via1 >>
rect 33440 16746 33818 17224
rect 131206 16750 131660 17264
rect 36762 10086 37016 10800
rect 127624 10114 128126 10758
<< metal2 >>
rect 3305 382079 3759 382237
rect 3305 381971 3427 382079
rect 3649 381971 3759 382079
rect 3305 379301 3759 381971
rect 3305 379165 3481 379301
rect 3597 379165 3759 379301
rect 3305 379121 3759 379165
rect 43661 344377 44243 344460
rect 43661 344307 43703 344377
rect 43767 344307 43841 344377
rect 43905 344307 43979 344377
rect 44043 344307 44117 344377
rect 44181 344307 44243 344377
rect 43661 336159 44243 344307
rect 43661 336041 43739 336159
rect 43871 336041 43991 336159
rect 44123 336041 44243 336159
rect 43661 335969 44243 336041
rect 43661 335851 43739 335969
rect 43871 335851 43991 335969
rect 44123 335851 44243 335969
rect 43661 335753 44243 335851
rect 43363 306697 43967 306767
rect 43363 306585 43393 306697
rect 43453 306585 43525 306697
rect 43585 306585 43657 306697
rect 43717 306585 43789 306697
rect 43849 306585 43967 306697
rect 43363 292947 43967 306585
rect 43363 292707 43447 292947
rect 43619 292707 43725 292947
rect 43897 292707 43967 292947
rect 43363 292543 43967 292707
rect 42575 268903 43475 269281
rect 42575 268749 42645 268903
rect 42711 268749 42811 268903
rect 42877 268749 42977 268903
rect 43043 268749 43143 268903
rect 43209 268749 43309 268903
rect 43375 268749 43475 268903
rect 42575 250345 43475 268749
rect 42575 249932 43691 250345
rect 42575 249654 42662 249932
rect 43608 249654 43691 249932
rect 42575 249445 43691 249654
rect 26048 231191 26774 231576
rect 26048 231043 26105 231191
rect 26199 231043 26271 231191
rect 26365 231043 26437 231191
rect 26531 231043 26603 231191
rect 26697 231043 26774 231191
rect 26048 122707 26774 231043
rect 27939 193395 28791 193697
rect 27939 193181 28009 193395
rect 28117 193181 28213 193395
rect 28321 193181 28417 193395
rect 28525 193181 28621 193395
rect 28729 193181 28791 193395
rect 25805 122391 26907 122707
rect 25805 122085 25899 122391
rect 26121 122085 26405 122391
rect 26627 122085 26907 122391
rect 25805 121981 26907 122085
rect 27939 79147 28791 193181
rect 27939 78783 28021 79147
rect 28185 78783 28307 79147
rect 28471 78783 28593 79147
rect 28757 78783 28791 79147
rect 27939 78703 28791 78783
rect 30243 155645 31045 155996
rect 30243 155563 30311 155645
rect 30399 155563 30513 155645
rect 30601 155563 30715 155645
rect 30803 155563 30917 155645
rect 31005 155563 31045 155645
rect 6147 42407 6895 42465
rect 6147 42341 6279 42407
rect 6363 42341 6459 42407
rect 6543 42341 6639 42407
rect 6723 42341 6895 42407
rect 6147 42229 6895 42341
rect 6365 5125 6601 42229
rect 30243 35831 31045 155563
rect 30243 35593 30329 35831
rect 30469 35593 30585 35831
rect 30725 35593 30841 35831
rect 30981 35593 31045 35831
rect 30243 35273 31045 35593
rect 33371 117822 33899 118389
rect 33371 117754 33424 117822
rect 33860 117754 33899 117822
rect 33371 17224 33899 117754
rect 33371 16746 33440 17224
rect 33818 16746 33899 17224
rect 33371 13415 33899 16746
rect 32801 13189 33899 13415
rect 32801 13057 32959 13189
rect 33105 13057 33293 13189
rect 33439 13057 33627 13189
rect 33773 13057 33899 13189
rect 32801 12887 33899 13057
rect 36721 80134 37057 80259
rect 36721 80062 36748 80134
rect 37010 80062 37057 80134
rect 36721 10800 37057 80062
rect 131110 17264 131760 17513
rect 131110 16750 131206 17264
rect 131660 16750 131760 17264
rect 36721 10086 36762 10800
rect 37016 10086 37057 10800
rect 36721 8547 37057 10086
rect 127554 10758 128204 10997
rect 127554 10114 127624 10758
rect 128126 10114 128204 10758
rect 36355 8445 37449 8547
rect 36355 8339 36469 8445
rect 36599 8339 36727 8445
rect 36857 8339 36985 8445
rect 37115 8339 37449 8445
rect 36355 8211 37449 8339
rect 6331 4872 6953 5125
rect 6331 4790 6376 4872
rect 6934 4790 6953 4872
rect 6331 4683 6953 4790
rect 127554 1188 128204 10114
rect 131110 1202 131760 16750
<< via2 >>
rect 3427 381971 3649 382079
rect 3481 379165 3597 379301
rect 43703 344307 43767 344377
rect 43841 344307 43905 344377
rect 43979 344307 44043 344377
rect 44117 344307 44181 344377
rect 43739 336041 43871 336159
rect 43991 336041 44123 336159
rect 43739 335851 43871 335969
rect 43991 335851 44123 335969
rect 43393 306585 43453 306697
rect 43525 306585 43585 306697
rect 43657 306585 43717 306697
rect 43789 306585 43849 306697
rect 43447 292707 43619 292947
rect 43725 292707 43897 292947
rect 42645 268749 42711 268903
rect 42811 268749 42877 268903
rect 42977 268749 43043 268903
rect 43143 268749 43209 268903
rect 43309 268749 43375 268903
rect 42662 249654 43608 249932
rect 26105 231043 26199 231191
rect 26271 231043 26365 231191
rect 26437 231043 26531 231191
rect 26603 231043 26697 231191
rect 28009 193181 28117 193395
rect 28213 193181 28321 193395
rect 28417 193181 28525 193395
rect 28621 193181 28729 193395
rect 25899 122085 26121 122391
rect 26405 122085 26627 122391
rect 28021 78783 28185 79147
rect 28307 78783 28471 79147
rect 28593 78783 28757 79147
rect 30311 155563 30399 155645
rect 30513 155563 30601 155645
rect 30715 155563 30803 155645
rect 30917 155563 31005 155645
rect 6279 42341 6363 42407
rect 6459 42341 6543 42407
rect 6639 42341 6723 42407
rect 30329 35593 30469 35831
rect 30585 35593 30725 35831
rect 30841 35593 30981 35831
rect 33424 117754 33860 117822
rect 32959 13057 33105 13189
rect 33293 13057 33439 13189
rect 33627 13057 33773 13189
rect 36748 80062 37010 80134
rect 36469 8339 36599 8445
rect 36727 8339 36857 8445
rect 36985 8339 37115 8445
rect 6376 4790 6934 4872
<< metal3 >>
rect 2485 649507 2785 649511
rect 2485 642919 9209 649507
rect 2485 642638 167671 642919
rect 2485 642596 83900 642638
rect 2485 636672 64252 642596
rect 71226 636672 83900 642596
rect 2485 636536 83900 636672
rect 91262 642612 167671 642638
rect 91262 636536 104358 642612
rect 2485 636510 104358 636536
rect 111720 642596 167671 642612
rect 111720 642580 144760 642596
rect 111720 636510 125348 642580
rect 2485 636478 125348 636510
rect 132710 636494 144760 642580
rect 152122 636494 167671 642596
rect 132710 636478 167671 636494
rect 2485 636195 167671 636478
rect 2485 634711 9209 636195
rect 3059 382079 44891 382157
rect 3059 381971 3427 382079
rect 3649 382071 44891 382079
rect 3649 382011 58864 382071
rect 3649 381971 44891 382011
rect 3059 381893 44891 381971
rect 3289 379301 3795 379357
rect 3289 379299 3481 379301
rect 1147 379187 3481 379299
rect 3289 379165 3481 379187
rect 3597 379299 3795 379301
rect 3597 379187 3925 379299
rect 3597 379165 3795 379187
rect 3289 379089 3795 379165
rect 43667 344388 44241 344409
rect 43667 344377 45554 344388
rect 43667 344373 43703 344377
rect 43637 344313 43703 344373
rect 43667 344307 43703 344313
rect 43767 344307 43841 344377
rect 43905 344307 43979 344377
rect 44043 344307 44117 344377
rect 44181 344307 45554 344377
rect 43667 344300 45554 344307
rect 43667 344277 44241 344300
rect 1883 336159 44308 336253
rect 1883 336079 43739 336159
rect 1267 336041 43739 336079
rect 43871 336041 43991 336159
rect 44123 336041 44308 336159
rect 1267 335969 44308 336041
rect 1267 335967 43739 335969
rect 1883 335851 43739 335967
rect 43871 335851 43991 335969
rect 44123 335851 44308 335969
rect 1883 335799 44308 335851
rect 43365 306697 43967 306735
rect 43365 306675 43393 306697
rect 43287 306615 43393 306675
rect 43365 306585 43393 306615
rect 43453 306585 43525 306697
rect 43585 306585 43657 306697
rect 43717 306585 43789 306697
rect 43849 306675 43967 306697
rect 43849 306615 53344 306675
rect 43849 306585 43967 306615
rect 43365 306539 43967 306585
rect 2061 292947 44090 293027
rect 2061 292855 43447 292947
rect 1293 292743 43447 292855
rect 2061 292707 43447 292743
rect 43619 292707 43725 292947
rect 43897 292707 44090 292947
rect 2061 292641 44090 292707
rect 42545 268903 43585 268955
rect 42545 268749 42645 268903
rect 42711 268749 42811 268903
rect 42877 268749 42977 268903
rect 43043 268749 43143 268903
rect 43209 268749 43309 268903
rect 43375 268855 43585 268903
rect 43375 268795 50032 268855
rect 43375 268749 43585 268795
rect 42545 268691 43585 268749
rect 1745 249932 43911 249985
rect 1745 249833 42662 249932
rect 1269 249721 42662 249833
rect 1745 249654 42662 249721
rect 43608 249654 43911 249932
rect 1745 249601 43911 249654
rect 25876 231191 45241 231223
rect 25876 231043 26105 231191
rect 26199 231043 26271 231191
rect 26365 231043 26437 231191
rect 26531 231043 26603 231191
rect 26697 231157 45241 231191
rect 26697 231097 60428 231157
rect 26697 231043 45241 231097
rect 25876 231013 45241 231043
rect 27720 193395 44835 193461
rect 27720 193181 28009 193395
rect 28117 193181 28213 193395
rect 28321 193181 28417 193395
rect 28525 193181 28621 193395
rect 28729 193337 44835 193395
rect 28729 193277 45340 193337
rect 28729 193181 44835 193277
rect 27720 193131 44835 193181
rect 2409 178001 3357 178557
rect 2409 177583 2553 178001
rect 2981 177583 3357 178001
rect 2409 177187 3357 177583
rect 2409 176769 2553 177187
rect 2981 176769 3357 177187
rect 2409 176373 3357 176769
rect 2409 175955 2553 176373
rect 2981 175955 3357 176373
rect 2409 175559 3357 175955
rect 2409 175141 2553 175559
rect 2981 175141 3357 175559
rect 2409 174745 3357 175141
rect 2409 174327 2553 174745
rect 2981 174327 3357 174745
rect 2409 168033 3357 174327
rect 2409 167615 2647 168033
rect 3075 167615 3357 168033
rect 2409 167219 3357 167615
rect 2409 166801 2647 167219
rect 3075 166801 3357 167219
rect 2409 166405 3357 166801
rect 2409 165987 2647 166405
rect 3075 165987 3357 166405
rect 2409 165591 3357 165987
rect 2409 165173 2647 165591
rect 3075 165173 3357 165591
rect 2409 164777 3357 165173
rect 2409 164359 2647 164777
rect 3075 164359 3357 164777
rect 2409 163757 3357 164359
rect 30058 155645 44623 155683
rect 30058 155563 30311 155645
rect 30399 155563 30513 155645
rect 30601 155563 30715 155645
rect 30803 155563 30917 155645
rect 31005 155639 44623 155645
rect 31005 155579 45340 155639
rect 31005 155563 44623 155579
rect 30058 155537 44623 155563
rect 25589 122391 27015 122505
rect 25589 122295 25899 122391
rect 1941 122211 25899 122295
rect 1233 122099 25899 122211
rect 1941 122085 25899 122099
rect 26121 122085 26405 122391
rect 26627 122295 27015 122391
rect 26627 122085 27413 122295
rect 1941 122035 27413 122085
rect 25589 121911 27015 122035
rect 33407 117822 33865 117845
rect 33407 117819 33424 117822
rect 33313 117759 33424 117819
rect 33407 117754 33424 117759
rect 33860 117819 33865 117822
rect 33860 117759 61716 117819
rect 33860 117754 33865 117759
rect 33407 117741 33865 117754
rect 36729 80134 37045 80161
rect 36729 80121 36748 80134
rect 36655 80062 36748 80121
rect 37010 80121 37045 80134
rect 37010 80062 51320 80121
rect 36655 80061 51320 80062
rect 36729 80031 37045 80061
rect 27849 79147 28963 79339
rect 27849 79107 28021 79147
rect 1667 78989 28021 79107
rect 1239 78877 28021 78989
rect 1667 78813 28021 78877
rect 27849 78783 28021 78813
rect 28185 78783 28307 79147
rect 28471 78783 28593 79147
rect 28757 78783 28963 79147
rect 27849 78661 28963 78783
rect 6201 42423 6859 42483
rect 6109 42407 47916 42423
rect 6109 42363 6279 42407
rect 6201 42341 6279 42363
rect 6363 42341 6459 42407
rect 6543 42341 6639 42407
rect 6723 42363 47916 42407
rect 6723 42341 6859 42363
rect 6201 42275 6859 42341
rect 2177 35831 31469 35973
rect 2177 35767 30329 35831
rect 1255 35655 30329 35767
rect 2177 35593 30329 35655
rect 30469 35593 30585 35831
rect 30725 35593 30841 35831
rect 30981 35593 31469 35831
rect 2177 35469 31469 35593
rect 32869 13189 33823 13281
rect 32869 13163 32959 13189
rect 1257 13057 32959 13163
rect 33105 13057 33293 13189
rect 33439 13057 33627 13189
rect 33773 13163 33823 13189
rect 33773 13057 34114 13163
rect 1257 13051 34114 13057
rect 32869 12973 33823 13051
rect 36385 8445 37403 8507
rect 36385 8435 36469 8445
rect 1281 8339 36469 8435
rect 36599 8339 36727 8445
rect 36857 8339 36985 8445
rect 37115 8435 37403 8445
rect 37115 8339 37990 8435
rect 1281 8323 37990 8339
rect 36385 8277 37403 8323
rect 6635 4889 6981 4905
rect 1201 4872 6981 4889
rect 1201 4790 6376 4872
rect 6934 4790 6981 4872
rect 1201 4777 6981 4790
rect 6635 4753 6981 4777
<< via3 >>
rect 64252 636672 71226 642596
rect 83900 636536 91262 642638
rect 104358 636510 111720 642612
rect 125348 636478 132710 642580
rect 144760 636494 152122 642596
rect 2553 177583 2981 178001
rect 2553 176769 2981 177187
rect 2553 175955 2981 176373
rect 2553 175141 2981 175559
rect 2553 174327 2981 174745
rect 2647 167615 3075 168033
rect 2647 166801 3075 167219
rect 2647 165987 3075 166405
rect 2647 165173 3075 165591
rect 2647 164359 3075 164777
<< metal4 >>
rect 63746 642596 71808 642951
rect 63746 636672 64252 642596
rect 71226 636672 71808 642596
rect 36623 352158 42195 353748
rect 36623 347340 36820 352158
rect 41964 347340 42195 352158
rect 36623 316462 42195 347340
rect 36623 311548 36802 316462
rect 41984 311548 42195 316462
rect 36623 280262 42195 311548
rect 36623 275486 36858 280262
rect 41958 275486 42195 280262
rect 36623 244230 42195 275486
rect 36623 239404 36882 244230
rect 42004 239404 42195 244230
rect 36623 207867 42195 239404
rect 36623 207179 37079 207867
rect 37965 207179 38705 207867
rect 39591 207179 40331 207867
rect 41217 207179 42195 207867
rect 36623 206541 42195 207179
rect 36623 205853 37079 206541
rect 37965 205853 38705 206541
rect 39591 205853 40331 206541
rect 41217 205853 42195 206541
rect 36623 205215 42195 205853
rect 36623 204527 37079 205215
rect 37965 204527 38705 205215
rect 39591 204527 40331 205215
rect 41217 204527 42195 205215
rect 2381 178001 3331 178263
rect 2381 177583 2553 178001
rect 2981 177723 3331 178001
rect 2381 177313 2703 177583
rect 3107 177313 3331 177723
rect 2381 177187 3331 177313
rect 2381 176769 2553 177187
rect 2981 177003 3331 177187
rect 2381 176593 2703 176769
rect 3107 176593 3331 177003
rect 2381 176373 3331 176593
rect 2381 175955 2553 176373
rect 2981 176283 3331 176373
rect 2381 175873 2703 175955
rect 3107 175873 3331 176283
rect 2381 175563 3331 175873
rect 2381 175559 2703 175563
rect 2381 175141 2553 175559
rect 3107 175153 3331 175563
rect 2981 175141 3331 175153
rect 2381 174843 3331 175141
rect 2381 174745 2703 174843
rect 2381 174327 2553 174745
rect 3107 174433 3331 174843
rect 2981 174327 3331 174433
rect 2381 174085 3331 174327
rect 36623 177819 42195 204527
rect 36623 177079 37179 177819
rect 37997 177079 38581 177819
rect 39399 177079 39983 177819
rect 40801 177079 42195 177819
rect 36623 176515 42195 177079
rect 36623 175775 37179 176515
rect 37997 175775 38581 176515
rect 39399 175775 39983 176515
rect 40801 175775 42195 176515
rect 36623 175211 42195 175775
rect 36623 174471 37179 175211
rect 37997 174471 38581 175211
rect 39399 174471 39983 175211
rect 40801 174471 42195 175211
rect 2521 168033 3471 168383
rect 2521 167615 2647 168033
rect 3075 167771 3471 168033
rect 2521 167361 2803 167615
rect 3207 167361 3471 167771
rect 2521 167219 3471 167361
rect 2521 166801 2647 167219
rect 3075 167051 3471 167219
rect 2521 166641 2803 166801
rect 3207 166641 3471 167051
rect 2521 166405 3471 166641
rect 2521 165987 2647 166405
rect 3075 166331 3471 166405
rect 2521 165921 2803 165987
rect 3207 165921 3471 166331
rect 2521 165611 3471 165921
rect 2521 165591 2803 165611
rect 2521 165173 2647 165591
rect 3207 165201 3471 165611
rect 3075 165173 3471 165201
rect 2521 164891 3471 165173
rect 2521 164777 2803 164891
rect 2521 164359 2647 164777
rect 3207 164481 3471 164891
rect 3075 164359 3471 164481
rect 2521 164205 3471 164359
rect 36623 167894 42195 174471
rect 36623 164574 36962 167894
rect 41870 164574 42195 167894
rect 36623 136222 42195 164574
rect 36623 131844 36764 136222
rect 42008 131844 42195 136222
rect 36623 100046 42195 131844
rect 36623 95716 36812 100046
rect 41874 95716 42195 100046
rect 36623 66520 42195 95716
rect 36623 62184 36804 66520
rect 41998 62184 42195 66520
rect 36623 60418 42195 62184
rect 48921 350098 49541 382259
rect 48921 347242 49010 350098
rect 49452 347242 49541 350098
rect 48921 314162 49541 347242
rect 48921 311486 49004 314162
rect 49442 311486 49541 314162
rect 48921 278126 49541 311486
rect 48921 275388 49016 278126
rect 49446 275388 49541 278126
rect 48921 242178 49541 275388
rect 48921 239268 48998 242178
rect 49456 239268 49541 242178
rect 48921 207699 49541 239268
rect 48921 207359 49047 207699
rect 49395 207359 49541 207699
rect 48921 206951 49541 207359
rect 48921 206611 49047 206951
rect 49395 206611 49541 206951
rect 48921 206203 49541 206611
rect 48921 205863 49047 206203
rect 49395 205863 49541 206203
rect 48921 205455 49541 205863
rect 48921 205115 49047 205455
rect 49395 205115 49541 205455
rect 48921 204707 49541 205115
rect 48921 204367 49047 204707
rect 49395 204367 49541 204707
rect 48921 177697 49541 204367
rect 48921 177343 49043 177697
rect 49419 177343 49541 177697
rect 48921 176953 49541 177343
rect 48921 176599 49043 176953
rect 49419 176599 49541 176953
rect 48921 176209 49541 176599
rect 48921 175855 49043 176209
rect 49419 175855 49541 176209
rect 48921 175465 49541 175855
rect 48921 175111 49043 175465
rect 49419 175111 49541 175465
rect 48921 174721 49541 175111
rect 48921 174367 49043 174721
rect 49419 174367 49541 174721
rect 48921 167855 49541 174367
rect 48921 167501 49073 167855
rect 49449 167501 49541 167855
rect 48921 167111 49541 167501
rect 48921 166757 49073 167111
rect 49449 166757 49541 167111
rect 48921 166367 49541 166757
rect 48921 166013 49073 166367
rect 49449 166013 49541 166367
rect 48921 165623 49541 166013
rect 48921 165269 49073 165623
rect 49449 165269 49541 165623
rect 48921 164879 49541 165269
rect 48921 164525 49073 164879
rect 49449 164525 49541 164879
rect 48921 134146 49541 164525
rect 48921 131760 49012 134146
rect 49450 131760 49541 134146
rect 48921 98136 49541 131760
rect 48921 95596 49030 98136
rect 49448 95596 49541 98136
rect 48921 66604 49541 95596
rect 48921 64408 49028 66604
rect 49408 64408 49541 66604
rect 48921 42259 49541 64408
rect 50161 42259 50781 382259
rect 63746 377104 71808 636672
rect 63746 376654 64162 377104
rect 68782 376654 71808 377104
rect 63746 376554 71808 376654
rect 83512 642638 91574 643159
rect 83512 636536 83900 642638
rect 91262 636536 91574 642638
rect 83512 377076 91574 636536
rect 83512 376604 83716 377076
rect 88746 376604 91574 377076
rect 83512 376470 91574 376604
rect 104050 642612 112112 643095
rect 104050 636510 104358 642612
rect 111720 636510 112112 642612
rect 104050 377080 112112 636510
rect 104050 376604 104244 377080
rect 108940 376604 112112 377080
rect 104050 376518 112112 376604
rect 124996 642580 133058 643095
rect 124996 636478 125348 642580
rect 132710 636478 133058 642580
rect 124996 377672 133058 636478
rect 144402 642596 152464 643095
rect 144402 636494 144760 642596
rect 152122 636494 152464 642596
rect 124996 377084 133062 377672
rect 144402 377480 152464 636494
rect 124996 376638 125230 377084
rect 128792 376638 133062 377084
rect 124996 376432 133062 376638
rect 144400 377132 152466 377480
rect 144400 376576 144642 377132
rect 148844 376576 152466 377132
rect 144400 376420 152466 376576
<< via4 >>
rect 36820 347340 41964 352158
rect 36802 311548 41984 316462
rect 36858 275486 41958 280262
rect 36882 239404 42004 244230
rect 37079 207179 37965 207867
rect 38705 207179 39591 207867
rect 40331 207179 41217 207867
rect 37079 205853 37965 206541
rect 38705 205853 39591 206541
rect 40331 205853 41217 206541
rect 37079 204527 37965 205215
rect 38705 204527 39591 205215
rect 40331 204527 41217 205215
rect 2703 177583 2981 177723
rect 2981 177583 3107 177723
rect 2703 177313 3107 177583
rect 2703 176769 2981 177003
rect 2981 176769 3107 177003
rect 2703 176593 3107 176769
rect 2703 175955 2981 176283
rect 2981 175955 3107 176283
rect 2703 175873 3107 175955
rect 2703 175559 3107 175563
rect 2703 175153 2981 175559
rect 2981 175153 3107 175559
rect 2703 174745 3107 174843
rect 2703 174433 2981 174745
rect 2981 174433 3107 174745
rect 37179 177079 37997 177819
rect 38581 177079 39399 177819
rect 39983 177079 40801 177819
rect 37179 175775 37997 176515
rect 38581 175775 39399 176515
rect 39983 175775 40801 176515
rect 37179 174471 37997 175211
rect 38581 174471 39399 175211
rect 39983 174471 40801 175211
rect 2803 167615 3075 167771
rect 3075 167615 3207 167771
rect 2803 167361 3207 167615
rect 2803 166801 3075 167051
rect 3075 166801 3207 167051
rect 2803 166641 3207 166801
rect 2803 165987 3075 166331
rect 3075 165987 3207 166331
rect 2803 165921 3207 165987
rect 2803 165591 3207 165611
rect 2803 165201 3075 165591
rect 3075 165201 3207 165591
rect 2803 164777 3207 164891
rect 2803 164481 3075 164777
rect 3075 164481 3207 164777
rect 36962 164574 41870 167894
rect 36764 131844 42008 136222
rect 36812 95716 41874 100046
rect 36804 62184 41998 66520
rect 49010 347242 49452 350098
rect 49004 311486 49442 314162
rect 49016 275388 49446 278126
rect 48998 239268 49456 242178
rect 49047 205863 49395 206203
rect 49047 205115 49395 205455
rect 49047 204367 49395 204707
rect 49043 177343 49419 177697
rect 49043 176599 49419 176953
rect 49043 175855 49419 176209
rect 49043 175111 49419 175465
rect 49043 174367 49419 174721
rect 49073 167501 49449 167855
rect 49073 166757 49449 167111
rect 49073 166013 49449 166367
rect 49073 165269 49449 165623
rect 49073 164525 49449 164879
rect 49012 131760 49450 134146
rect 49030 95596 49448 98136
rect 49028 64408 49408 66604
rect 64162 376654 68782 377104
rect 83716 376604 88746 377076
rect 104244 376604 108940 377080
rect 125230 376638 128792 377084
rect 144642 376576 148844 377132
<< metal5 >>
rect 45077 377787 165045 378407
rect 45077 377132 165045 377167
rect 45077 377104 144642 377132
rect 45077 376654 64162 377104
rect 68782 377084 144642 377104
rect 68782 377080 125230 377084
rect 68782 377076 104244 377080
rect 68782 376654 83716 377076
rect 45077 376604 83716 376654
rect 88746 376604 104244 377076
rect 108940 376638 125230 377080
rect 128792 376638 144642 377084
rect 108940 376604 144642 376638
rect 45077 376576 144642 376604
rect 148844 376576 165045 377132
rect 45077 376547 165045 376576
rect 36320 352158 49689 352400
rect 36320 347340 36820 352158
rect 41964 350098 49689 352158
rect 41964 347340 49010 350098
rect 36320 347242 49010 347340
rect 49452 347242 49689 350098
rect 36320 347122 49689 347242
rect 36426 316462 49795 316640
rect 36426 311548 36802 316462
rect 41984 314162 49795 316462
rect 41984 311548 49004 314162
rect 36426 311486 49004 311548
rect 49442 311486 49795 314162
rect 36426 311362 49795 311486
rect 36327 280262 49696 280556
rect 36327 275486 36858 280262
rect 41958 278126 49696 280262
rect 41958 275486 49016 278126
rect 36327 275388 49016 275486
rect 49446 275388 49696 278126
rect 36327 275278 49696 275388
rect 36432 244230 49660 244456
rect 36432 239404 36882 244230
rect 42004 242178 49660 244230
rect 42004 239404 48998 242178
rect 36432 239268 48998 239404
rect 49456 239268 49660 242178
rect 36432 239178 49660 239268
rect 36525 207867 49559 208537
rect 36525 207179 37079 207867
rect 37965 207179 38705 207867
rect 39591 207179 40331 207867
rect 41217 207179 49559 207867
rect 36525 206541 49559 207179
rect 36525 205853 37079 206541
rect 37965 205853 38705 206541
rect 39591 205853 40331 206541
rect 41217 206203 49559 206541
rect 41217 205863 49047 206203
rect 49395 205863 49559 206203
rect 41217 205853 49559 205863
rect 36525 205455 49559 205853
rect 36525 205215 49047 205455
rect 36525 204527 37079 205215
rect 37965 204527 38705 205215
rect 39591 204527 40331 205215
rect 41217 205115 49047 205215
rect 49395 205115 49559 205455
rect 41217 204707 49559 205115
rect 41217 204527 49047 204707
rect 36525 204367 49047 204527
rect 49395 204367 49559 204707
rect 36525 204165 49559 204367
rect 2523 177819 49694 178147
rect 2523 177723 37179 177819
rect 2523 177313 2703 177723
rect 3107 177313 37179 177723
rect 2523 177079 37179 177313
rect 37997 177079 38581 177819
rect 39399 177079 39983 177819
rect 40801 177697 49694 177819
rect 40801 177343 49043 177697
rect 49419 177343 49694 177697
rect 40801 177079 49694 177343
rect 2523 177003 49694 177079
rect 2523 176593 2703 177003
rect 3107 176953 49694 177003
rect 3107 176599 49043 176953
rect 49419 176599 49694 176953
rect 3107 176593 49694 176599
rect 2523 176515 49694 176593
rect 2523 176283 37179 176515
rect 2523 175873 2703 176283
rect 3107 175873 37179 176283
rect 2523 175775 37179 175873
rect 37997 175775 38581 176515
rect 39399 175775 39983 176515
rect 40801 176209 49694 176515
rect 40801 175855 49043 176209
rect 49419 175855 49694 176209
rect 40801 175775 49694 175855
rect 2523 175563 49694 175775
rect 2523 175153 2703 175563
rect 3107 175465 49694 175563
rect 3107 175211 49043 175465
rect 3107 175153 37179 175211
rect 2523 174843 37179 175153
rect 2523 174433 2703 174843
rect 3107 174471 37179 174843
rect 37997 174471 38581 175211
rect 39399 174471 39983 175211
rect 40801 175111 49043 175211
rect 49419 175111 49694 175465
rect 40801 174721 49694 175111
rect 40801 174471 49043 174721
rect 3107 174433 49043 174471
rect 2523 174367 49043 174433
rect 49419 174367 49694 174721
rect 2523 174217 49694 174367
rect 2613 167894 49836 168229
rect 2613 167771 36962 167894
rect 2613 167361 2803 167771
rect 3207 167361 36962 167771
rect 2613 167051 36962 167361
rect 2613 166641 2803 167051
rect 3207 166641 36962 167051
rect 2613 166331 36962 166641
rect 2613 165921 2803 166331
rect 3207 165921 36962 166331
rect 2613 165611 36962 165921
rect 2613 165201 2803 165611
rect 3207 165201 36962 165611
rect 2613 164891 36962 165201
rect 2613 164481 2803 164891
rect 3207 164574 36962 164891
rect 41870 167855 49836 167894
rect 41870 167501 49073 167855
rect 49449 167501 49836 167855
rect 41870 167111 49836 167501
rect 41870 166757 49073 167111
rect 49449 166757 49836 167111
rect 41870 166367 49836 166757
rect 41870 166013 49073 166367
rect 49449 166013 49836 166367
rect 41870 165623 49836 166013
rect 41870 165269 49073 165623
rect 49449 165269 49836 165623
rect 41870 164879 49836 165269
rect 41870 164574 49073 164879
rect 3207 164525 49073 164574
rect 49449 164525 49836 164879
rect 3207 164481 49836 164525
rect 2613 164299 49836 164481
rect 36614 136222 49642 136476
rect 36614 131844 36764 136222
rect 42008 134146 49642 136222
rect 42008 131844 49012 134146
rect 36614 131760 49012 131844
rect 49450 131760 49642 134146
rect 36614 131642 49642 131760
rect 36626 100046 49654 100310
rect 36626 95716 36812 100046
rect 41874 98136 49654 100046
rect 41874 95716 49030 98136
rect 36626 95596 49030 95716
rect 49448 95596 49654 98136
rect 36626 95476 49654 95596
rect 36588 66604 49616 66768
rect 36588 66520 49028 66604
rect 36588 62184 36804 66520
rect 41998 64408 49028 66520
rect 49408 64408 49616 66604
rect 41998 62184 49616 64408
rect 36588 61934 49616 62184
use puf_super  puf_super_0
timestamp 1656715967
transform 1 0 45077 0 1 42259
box 0 0 119968 340000
use sky130_fd_pr__res_generic_m1_DBNWX4  sky130_fd_pr__res_generic_m1_DBNWX4_0
timestamp 1656715967
transform 0 1 40193 -1 0 16982
box -500 -557 500 557
use sky130_fd_pr__res_generic_m1_DBNWX4  sky130_fd_pr__res_generic_m1_DBNWX4_1
timestamp 1656715967
transform 0 1 43603 -1 0 10422
box -500 -557 500 557
<< end >>
