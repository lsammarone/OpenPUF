magic
tech sky130A
magscale 1 2
timestamp 1483428465
<< checkpaint >>
rect -1411 -1413 1411 1413
<< pwell >>
rect -151 -91 151 91
<< nmos >>
rect -63 -65 -33 65
rect 33 -65 63 65
<< ndiff >>
rect -125 51 -63 65
rect -125 17 -113 51
rect -79 17 -63 51
rect -125 -17 -63 17
rect -125 -51 -113 -17
rect -79 -51 -63 -17
rect -125 -65 -63 -51
rect -33 51 33 65
rect -33 17 -17 51
rect 17 17 33 51
rect -33 -17 33 17
rect -33 -51 -17 -17
rect 17 -51 33 -17
rect -33 -65 33 -51
rect 63 51 125 65
rect 63 17 79 51
rect 113 17 125 51
rect 63 -17 125 17
rect 63 -51 79 -17
rect 113 -51 125 -17
rect 63 -65 125 -51
<< ndiffc >>
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -17 17 17 51
rect -17 -51 17 -17
rect 79 17 113 51
rect 79 -51 113 -17
<< poly >>
rect 15 137 81 153
rect 15 103 31 137
rect 65 103 81 137
rect -63 65 -33 91
rect 15 87 81 103
rect 33 65 63 87
rect -63 -87 -33 -65
rect -81 -103 -15 -87
rect 33 -91 63 -65
rect -81 -137 -65 -103
rect -31 -137 -15 -103
rect -81 -153 -15 -137
<< polycont >>
rect 31 103 65 137
rect -65 -137 -31 -103
<< locali >>
rect 15 103 31 137
rect 65 103 81 137
rect -113 53 -79 69
rect -113 -17 -79 17
rect -113 -69 -79 -53
rect -17 53 17 69
rect -17 -17 17 17
rect -17 -69 17 -53
rect 79 53 113 69
rect 79 -17 113 17
rect 79 -69 113 -53
rect -81 -137 -65 -103
rect -31 -137 -15 -103
<< viali >>
rect 31 103 65 137
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect -65 -137 -31 -103
<< metal1 >>
rect 19 137 77 143
rect 19 103 31 137
rect 65 103 77 137
rect 19 97 77 103
rect -119 53 -73 65
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -65 -73 -53
rect -23 53 23 65
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -65 23 -53
rect 73 53 119 65
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -65 119 -53
rect -77 -103 -19 -97
rect -77 -137 -65 -103
rect -31 -137 -19 -103
rect -77 -143 -19 -137
<< end >>
