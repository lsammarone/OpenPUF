magic
tech sky130A
magscale 1 2
timestamp 1655322987
<< metal4 >>
rect -309 918 309 981
rect -309 -918 -278 918
rect 278 -918 309 918
rect -309 -981 309 -918
<< via4 >>
rect -278 -918 278 918
<< metal5 >>
rect -309 918 309 981
rect -309 -918 -278 918
rect 278 -918 309 918
rect -309 -981 309 -918
<< end >>
