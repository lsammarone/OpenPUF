magic
tech sky130A
magscale 1 2
timestamp 1483428465
<< checkpaint >>
rect -1478 -1293 1478 1293
<< metal3 >>
rect -218 32 218 33
rect -218 -32 -192 32
rect -128 -32 -112 32
rect -48 -32 -32 32
rect 32 -32 48 32
rect 112 -32 128 32
rect 192 -32 218 32
rect -218 -33 218 -32
<< via3 >>
rect -192 -32 -128 32
rect -112 -32 -48 32
rect -32 -32 32 32
rect 48 -32 112 32
rect 128 -32 192 32
<< metal4 >>
rect -218 32 218 33
rect -218 -32 -192 32
rect -128 -32 -112 32
rect -48 -32 -32 32
rect 32 -32 48 32
rect 112 -32 128 32
rect 192 -32 218 32
rect -218 -33 218 -32
<< end >>
