magic
tech sky130A
magscale 1 2
timestamp 1656729169
<< metal2 >>
rect -662 28 662 33
rect -662 -28 -628 28
rect -572 -28 -548 28
rect -492 -28 -468 28
rect -412 -28 -388 28
rect -332 -28 -308 28
rect -252 -28 -228 28
rect -172 -28 -148 28
rect -92 -28 -68 28
rect -12 -28 12 28
rect 68 -28 92 28
rect 148 -28 172 28
rect 228 -28 252 28
rect 308 -28 332 28
rect 388 -28 412 28
rect 468 -28 492 28
rect 548 -28 572 28
rect 628 -28 662 28
rect -662 -33 662 -28
<< via2 >>
rect -628 -28 -572 28
rect -548 -28 -492 28
rect -468 -28 -412 28
rect -388 -28 -332 28
rect -308 -28 -252 28
rect -228 -28 -172 28
rect -148 -28 -92 28
rect -68 -28 -12 28
rect 12 -28 68 28
rect 92 -28 148 28
rect 172 -28 228 28
rect 252 -28 308 28
rect 332 -28 388 28
rect 412 -28 468 28
rect 492 -28 548 28
rect 572 -28 628 28
<< metal3 >>
rect -662 28 662 33
rect -662 -28 -628 28
rect -572 -28 -548 28
rect -492 -28 -468 28
rect -412 -28 -388 28
rect -332 -28 -308 28
rect -252 -28 -228 28
rect -172 -28 -148 28
rect -92 -28 -68 28
rect -12 -28 12 28
rect 68 -28 92 28
rect 148 -28 172 28
rect 228 -28 252 28
rect 308 -28 332 28
rect 388 -28 412 28
rect 468 -28 492 28
rect 548 -28 572 28
rect 628 -28 662 28
rect -662 -33 662 -28
<< properties >>
string GDS_END 9359802
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/merge/design_merged.gds
string GDS_START 9358646
<< end >>
