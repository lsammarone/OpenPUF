magic
tech sky130A
timestamp 1656715967
<< metal1 >>
rect -500 13 500 24
rect -500 -13 -493 13
rect -467 -13 -461 13
rect -435 -13 -429 13
rect -403 -13 -397 13
rect -371 -13 -365 13
rect -339 -13 -333 13
rect -307 -13 -301 13
rect -275 -13 -269 13
rect -243 -13 -237 13
rect -211 -13 -205 13
rect -179 -13 -173 13
rect -147 -13 -141 13
rect -115 -13 -109 13
rect -83 -13 -77 13
rect -51 -13 -45 13
rect -19 -13 -13 13
rect 13 -13 19 13
rect 45 -13 51 13
rect 77 -13 83 13
rect 109 -13 115 13
rect 141 -13 147 13
rect 173 -13 179 13
rect 205 -13 211 13
rect 237 -13 243 13
rect 269 -13 275 13
rect 301 -13 307 13
rect 333 -13 339 13
rect 365 -13 371 13
rect 397 -13 403 13
rect 429 -13 435 13
rect 461 -13 467 13
rect 493 -13 500 13
rect -500 -24 500 -13
<< via1 >>
rect -493 -13 -467 13
rect -461 -13 -435 13
rect -429 -13 -403 13
rect -397 -13 -371 13
rect -365 -13 -339 13
rect -333 -13 -307 13
rect -301 -13 -275 13
rect -269 -13 -243 13
rect -237 -13 -211 13
rect -205 -13 -179 13
rect -173 -13 -147 13
rect -141 -13 -115 13
rect -109 -13 -83 13
rect -77 -13 -51 13
rect -45 -13 -19 13
rect -13 -13 13 13
rect 19 -13 45 13
rect 51 -13 77 13
rect 83 -13 109 13
rect 115 -13 141 13
rect 147 -13 173 13
rect 179 -13 205 13
rect 211 -13 237 13
rect 243 -13 269 13
rect 275 -13 301 13
rect 307 -13 333 13
rect 339 -13 365 13
rect 371 -13 397 13
rect 403 -13 429 13
rect 435 -13 461 13
rect 467 -13 493 13
<< metal2 >>
rect -500 13 500 24
rect -500 -13 -493 13
rect -467 -13 -461 13
rect -435 -13 -429 13
rect -403 -13 -397 13
rect -371 -13 -365 13
rect -339 -13 -333 13
rect -307 -13 -301 13
rect -275 -13 -269 13
rect -243 -13 -237 13
rect -211 -13 -205 13
rect -179 -13 -173 13
rect -147 -13 -141 13
rect -115 -13 -109 13
rect -83 -13 -77 13
rect -51 -13 -45 13
rect -19 -13 -13 13
rect 13 -13 19 13
rect 45 -13 51 13
rect 77 -13 83 13
rect 109 -13 115 13
rect 141 -13 147 13
rect 173 -13 179 13
rect 205 -13 211 13
rect 237 -13 243 13
rect 269 -13 275 13
rect 301 -13 307 13
rect 333 -13 339 13
rect 365 -13 371 13
rect 397 -13 403 13
rect 429 -13 435 13
rect 461 -13 467 13
rect 493 -13 500 13
rect -500 -24 500 -13
<< properties >>
string GDS_END 9312454
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/design_merged.gds
string GDS_START 9310338
<< end >>
