magic
tech sky130A
magscale 1 2
timestamp 1483428465
<< checkpaint >>
rect -1663 -1440 1663 1440
<< metal3 >>
rect -403 152 403 180
rect -403 -152 -392 152
rect 392 -152 403 152
rect -403 -180 403 -152
<< via3 >>
rect -392 -152 392 152
<< metal4 >>
rect -403 152 403 180
rect -403 -152 -392 152
rect 392 -152 403 152
rect -403 -180 403 -152
<< end >>
