magic
tech sky130A
timestamp 1654736712
<< metal2 >>
rect -500 14 500 24
rect -500 -14 -494 14
rect -466 -14 -454 14
rect -426 -14 -414 14
rect -386 -14 -374 14
rect -346 -14 -334 14
rect -306 -14 -294 14
rect -266 -14 -254 14
rect -226 -14 -214 14
rect -186 -14 -174 14
rect -146 -14 -134 14
rect -106 -14 -94 14
rect -66 -14 -54 14
rect -26 -14 -14 14
rect 14 -14 26 14
rect 54 -14 66 14
rect 94 -14 106 14
rect 134 -14 146 14
rect 174 -14 186 14
rect 214 -14 226 14
rect 254 -14 266 14
rect 294 -14 306 14
rect 334 -14 346 14
rect 374 -14 386 14
rect 414 -14 426 14
rect 454 -14 466 14
rect 494 -14 500 14
rect -500 -24 500 -14
<< via2 >>
rect -494 -14 -466 14
rect -454 -14 -426 14
rect -414 -14 -386 14
rect -374 -14 -346 14
rect -334 -14 -306 14
rect -294 -14 -266 14
rect -254 -14 -226 14
rect -214 -14 -186 14
rect -174 -14 -146 14
rect -134 -14 -106 14
rect -94 -14 -66 14
rect -54 -14 -26 14
rect -14 -14 14 14
rect 26 -14 54 14
rect 66 -14 94 14
rect 106 -14 134 14
rect 146 -14 174 14
rect 186 -14 214 14
rect 226 -14 254 14
rect 266 -14 294 14
rect 306 -14 334 14
rect 346 -14 374 14
rect 386 -14 414 14
rect 426 -14 454 14
rect 466 -14 494 14
<< metal3 >>
rect -500 14 500 24
rect -500 -14 -494 14
rect -466 -14 -454 14
rect -426 -14 -414 14
rect -386 -14 -374 14
rect -346 -14 -334 14
rect -306 -14 -294 14
rect -266 -14 -254 14
rect -226 -14 -214 14
rect -186 -14 -174 14
rect -146 -14 -134 14
rect -106 -14 -94 14
rect -66 -14 -54 14
rect -26 -14 -14 14
rect 14 -14 26 14
rect 54 -14 66 14
rect 94 -14 106 14
rect 134 -14 146 14
rect 174 -14 186 14
rect 214 -14 226 14
rect 254 -14 266 14
rect 294 -14 306 14
rect 334 -14 346 14
rect 374 -14 386 14
rect 414 -14 426 14
rect 454 -14 466 14
rect 494 -14 500 14
rect -500 -24 500 -14
<< end >>
