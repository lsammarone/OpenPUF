magic
tech sky130A
magscale 1 2
timestamp 1483428465
<< checkpaint >>
rect -1283 -1289 1283 1289
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -23 17 23 29
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -29 23 -17
<< end >>
