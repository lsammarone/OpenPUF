magic
tech sky130A
timestamp 1654736712
<< metal4 >>
rect -500 129 500 184
rect -500 -149 -425 129
rect 333 -149 500 129
rect -500 -184 500 -149
<< via4 >>
rect -425 -149 333 129
<< metal5 >>
rect -500 129 500 184
rect -500 -149 -425 129
rect 333 -149 500 129
rect -500 -184 500 -149
<< end >>
