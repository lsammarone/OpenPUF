magic
tech sky130A
magscale 1 2
timestamp 1656729169
<< nwell >>
rect 31039 9642 31151 9963
rect 31318 9642 31407 9963
<< viali >>
rect 28312 9722 28346 9756
rect 29829 9735 29863 9769
rect 29997 9735 30031 9769
rect 30165 9735 30199 9769
rect 30333 9735 30367 9769
rect 30501 9735 30535 9769
rect 30669 9735 30703 9769
rect 30837 9735 30871 9769
rect 31577 9734 31611 9768
rect 31745 9734 31779 9768
rect 31913 9734 31947 9768
rect 32081 9734 32115 9768
rect 32249 9734 32283 9768
rect 32417 9734 32451 9768
rect 32585 9734 32619 9768
rect 28126 9596 28160 9630
rect 28801 9602 28835 9636
rect 28883 9602 28917 9636
rect 28974 9602 29008 9636
rect 29068 9602 29102 9636
rect 29388 9595 29422 9629
rect 29589 9600 29623 9634
rect 29708 9600 29742 9634
rect 29827 9600 29861 9634
rect 29946 9600 29980 9634
rect 30065 9600 30099 9634
rect 30184 9600 30218 9634
rect 30303 9600 30337 9634
rect 31513 9602 31547 9636
rect 31632 9602 31666 9636
rect 31751 9602 31785 9636
rect 31870 9602 31904 9636
rect 31989 9602 32023 9636
rect 32108 9602 32142 9636
rect 32227 9602 32261 9636
<< metal1 >>
rect 338 13891 1233 13911
rect 338 13887 1175 13891
rect 338 13835 357 13887
rect 409 13839 1175 13887
rect 1227 13839 1233 13891
rect 409 13835 1233 13839
rect 338 13814 1233 13835
rect 266 13418 1240 13435
rect 198 13412 1240 13418
rect 198 13398 1172 13412
rect 198 13346 214 13398
rect 266 13360 1172 13398
rect 1224 13360 1240 13412
rect 266 13346 1240 13360
rect 198 13338 1240 13346
rect 63486 13150 64108 13226
rect 0 12219 29658 12224
rect 62092 12221 64102 12222
rect 0 12167 29568 12219
rect 29620 12167 29658 12219
rect 0 12163 29658 12167
rect 31417 12216 64102 12221
rect 31417 12164 31455 12216
rect 31507 12164 64102 12216
rect 0 12162 490 12163
rect 31417 12160 64102 12164
rect 0 12077 27750 12082
rect 62092 12079 64102 12080
rect 0 12025 27680 12077
rect 27732 12025 27750 12077
rect 0 12021 27750 12025
rect 33325 12074 64102 12079
rect 33325 12022 33343 12074
rect 33395 12022 64102 12074
rect 0 12020 490 12021
rect 33325 12018 64102 12022
rect 0 11936 25892 11940
rect 62092 11937 64102 11938
rect 0 11884 25793 11936
rect 25845 11884 25892 11936
rect 0 11879 25892 11884
rect 35183 11933 64102 11937
rect 35183 11881 35230 11933
rect 35282 11881 64102 11933
rect 0 11878 490 11879
rect 35183 11876 64102 11881
rect 0 11795 23968 11798
rect 62092 11795 64102 11796
rect 0 11743 23904 11795
rect 23956 11743 23968 11795
rect 0 11737 23968 11743
rect 37107 11792 64102 11795
rect 37107 11740 37119 11792
rect 37171 11740 64102 11792
rect 0 11736 490 11737
rect 37107 11734 64102 11740
rect 0 11652 22092 11656
rect 62092 11653 64102 11654
rect 0 11600 22016 11652
rect 22068 11600 22092 11652
rect 0 11595 22092 11600
rect 38983 11649 64102 11653
rect 38983 11597 39007 11649
rect 39059 11597 64102 11649
rect 0 11594 490 11595
rect 38983 11592 64102 11597
rect 0 11509 20210 11514
rect 62092 11511 64102 11512
rect 0 11457 20126 11509
rect 20178 11457 20210 11509
rect 0 11453 20210 11457
rect 40865 11506 64102 11511
rect 40865 11454 40897 11506
rect 40949 11454 64102 11506
rect 0 11452 490 11453
rect 40865 11450 64102 11454
rect 0 11368 18302 11372
rect 62092 11369 64102 11370
rect 0 11316 18240 11368
rect 18292 11316 18302 11368
rect 0 11311 18302 11316
rect 42773 11365 64102 11369
rect 42773 11313 42783 11365
rect 42835 11313 64102 11365
rect 0 11310 490 11311
rect 42773 11308 64102 11313
rect 0 11225 16426 11230
rect 62092 11227 64102 11228
rect 0 11173 16352 11225
rect 16404 11173 16426 11225
rect 0 11169 16426 11173
rect 44649 11222 64102 11227
rect 44649 11170 44671 11222
rect 44723 11170 64102 11222
rect 0 11168 490 11169
rect 44649 11166 64102 11170
rect 0 11083 14556 11088
rect 62092 11085 64102 11086
rect 0 11031 14471 11083
rect 14523 11031 14556 11083
rect 0 11027 14556 11031
rect 46519 11080 64102 11085
rect 46519 11028 46552 11080
rect 46604 11028 64102 11080
rect 0 11026 490 11027
rect 46519 11024 64102 11028
rect 0 10940 12684 10946
rect 62092 10943 64102 10944
rect 0 10888 12583 10940
rect 12635 10888 12684 10940
rect 0 10885 12684 10888
rect 48391 10937 64102 10943
rect 48391 10885 48440 10937
rect 48492 10885 64102 10937
rect 0 10884 490 10885
rect 48391 10882 64102 10885
rect 0 10798 10798 10804
rect 62092 10801 64102 10802
rect 0 10746 10695 10798
rect 10747 10746 10798 10798
rect 0 10743 10798 10746
rect 50277 10800 60256 10801
rect 61624 10800 64102 10801
rect 50277 10795 64102 10800
rect 50277 10743 50328 10795
rect 50380 10743 64102 10795
rect 0 10742 490 10743
rect 50277 10740 64102 10743
rect 60159 10739 62096 10740
rect 0 10656 8887 10662
rect 62092 10659 64102 10660
rect 0 10604 8808 10656
rect 8860 10604 8887 10656
rect 0 10601 8887 10604
rect 52188 10653 64102 10659
rect 52188 10601 52215 10653
rect 52267 10601 64102 10653
rect 0 10600 490 10601
rect 52188 10598 64102 10601
rect 0 10515 7011 10520
rect 62092 10517 64102 10518
rect 0 10463 6918 10515
rect 6970 10463 7011 10515
rect 0 10459 7011 10463
rect 54064 10512 64102 10517
rect 54064 10460 54105 10512
rect 54157 10460 64102 10512
rect 0 10458 490 10459
rect 54064 10456 64102 10460
rect 0 10373 5114 10378
rect 62092 10375 64102 10376
rect 0 10321 5031 10373
rect 5083 10321 5114 10373
rect 0 10317 5114 10321
rect 55961 10370 64102 10375
rect 55961 10318 55992 10370
rect 56044 10318 64102 10370
rect 0 10316 490 10317
rect 55961 10314 64102 10318
rect 0 10230 3242 10236
rect 62092 10233 64102 10234
rect 0 10178 3142 10230
rect 3194 10178 3242 10230
rect 0 10175 3242 10178
rect 57833 10227 64102 10233
rect 57833 10175 57881 10227
rect 57933 10175 64102 10227
rect 0 10174 490 10175
rect 57833 10172 64102 10175
rect 0 10089 1383 10094
rect 62092 10091 64102 10092
rect 0 10037 1254 10089
rect 1306 10037 1383 10089
rect 0 10033 1383 10037
rect 59692 10086 64102 10091
rect 59692 10034 59769 10086
rect 59821 10034 64102 10086
rect 0 10032 490 10033
rect 59692 10030 64102 10034
rect 28549 9877 28625 9973
rect 29453 9877 29529 9973
rect 31001 9877 31188 9973
rect 31280 9877 31467 9973
rect 62092 9949 64102 9950
rect 59927 9944 64102 9949
rect 59927 9892 59999 9944
rect 60051 9892 64102 9944
rect 59927 9888 64102 9892
rect 0 9808 3464 9810
rect 0 9756 3368 9808
rect 3420 9756 3464 9808
rect 62092 9807 64102 9808
rect 58068 9805 64102 9807
rect 0 9749 3464 9756
rect 28302 9756 28355 9773
rect 0 9748 490 9749
rect 28302 9722 28312 9756
rect 28346 9722 28355 9756
rect 0 9663 5375 9668
rect 0 9611 5257 9663
rect 5309 9611 5375 9663
rect 0 9607 5375 9611
rect 7610 9652 7957 9674
rect 7610 9640 28178 9652
rect 0 9606 490 9607
rect 7610 9588 7699 9640
rect 7751 9588 7797 9640
rect 7849 9630 28178 9640
rect 7849 9596 28126 9630
rect 28160 9596 28178 9630
rect 7849 9588 28178 9596
rect 28302 9651 28355 9722
rect 29817 9769 32634 9794
rect 29817 9735 29829 9769
rect 29863 9735 29997 9769
rect 30031 9735 30165 9769
rect 30199 9735 30333 9769
rect 30367 9735 30501 9769
rect 30535 9735 30669 9769
rect 30703 9735 30837 9769
rect 30871 9768 32634 9769
rect 30871 9760 31577 9768
rect 30871 9735 31049 9760
rect 29817 9708 31049 9735
rect 31101 9708 31152 9760
rect 31204 9708 31255 9760
rect 31307 9708 31358 9760
rect 31410 9734 31577 9760
rect 31611 9734 31745 9768
rect 31779 9734 31913 9768
rect 31947 9734 32081 9768
rect 32115 9734 32249 9768
rect 32283 9734 32417 9768
rect 32451 9734 32585 9768
rect 32619 9734 32634 9768
rect 58068 9753 58112 9805
rect 58164 9753 64102 9805
rect 58068 9746 64102 9753
rect 31410 9708 32634 9734
rect 29817 9686 32634 9708
rect 62092 9665 64102 9666
rect 56157 9660 64102 9665
rect 28302 9636 29147 9651
rect 28302 9602 28801 9636
rect 28835 9602 28883 9636
rect 28917 9602 28974 9636
rect 29008 9602 29068 9636
rect 29102 9602 29147 9636
rect 28302 9590 29147 9602
rect 29366 9636 32557 9645
rect 29366 9634 31513 9636
rect 29366 9629 29589 9634
rect 29366 9595 29388 9629
rect 29422 9600 29589 9629
rect 29623 9600 29708 9634
rect 29742 9600 29827 9634
rect 29861 9600 29946 9634
rect 29980 9600 30065 9634
rect 30099 9600 30184 9634
rect 30218 9600 30303 9634
rect 30337 9602 31513 9634
rect 31547 9602 31632 9636
rect 31666 9602 31751 9636
rect 31785 9602 31870 9636
rect 31904 9602 31989 9636
rect 32023 9602 32108 9636
rect 32142 9602 32227 9636
rect 32261 9602 32557 9636
rect 56157 9608 56223 9660
rect 56275 9608 64102 9660
rect 56157 9604 64102 9608
rect 30337 9600 32557 9602
rect 29422 9595 32557 9600
rect 29366 9588 32557 9595
rect 7610 9578 28178 9588
rect 7610 9550 7957 9578
rect 0 9522 7221 9526
rect 62092 9523 64102 9524
rect 0 9470 7146 9522
rect 7198 9470 7221 9522
rect 0 9465 7221 9470
rect 54311 9519 64102 9523
rect 54311 9467 54334 9519
rect 54386 9467 64102 9519
rect 0 9464 490 9465
rect 54311 9462 64102 9467
rect 0 9378 9112 9384
rect 0 9326 9033 9378
rect 9085 9326 9112 9378
rect 28549 9333 28625 9429
rect 29453 9332 29529 9428
rect 31001 9333 31188 9429
rect 31280 9333 31467 9429
rect 62092 9381 64102 9382
rect 52420 9375 64102 9381
rect 0 9323 9112 9326
rect 52420 9323 52447 9375
rect 52499 9323 64102 9375
rect 0 9322 490 9323
rect 52420 9320 64102 9323
rect 0 9237 11000 9242
rect 62092 9239 64102 9240
rect 0 9185 10921 9237
rect 10973 9185 11000 9237
rect 0 9181 11000 9185
rect 50532 9234 64102 9239
rect 50532 9182 50559 9234
rect 50611 9182 64102 9234
rect 0 9180 490 9181
rect 50532 9178 64102 9182
rect 0 9095 12901 9100
rect 62092 9097 64102 9098
rect 0 9043 12810 9095
rect 12862 9043 12901 9095
rect 0 9039 12901 9043
rect 48631 9092 64102 9097
rect 48631 9040 48670 9092
rect 48722 9040 64102 9092
rect 0 9038 490 9039
rect 48631 9036 64102 9040
rect 0 8950 14776 8958
rect 62092 8955 64102 8956
rect 0 8898 14698 8950
rect 14750 8898 14776 8950
rect 0 8897 14776 8898
rect 46756 8947 64102 8955
rect 0 8896 490 8897
rect 46756 8895 46782 8947
rect 46834 8895 64102 8947
rect 46756 8894 64102 8895
rect 0 8811 16687 8816
rect 62092 8813 64102 8814
rect 0 8759 16576 8811
rect 16628 8759 16687 8811
rect 0 8755 16687 8759
rect 44845 8808 64102 8813
rect 44845 8756 44904 8808
rect 44956 8756 64102 8808
rect 0 8754 490 8755
rect 44845 8752 64102 8756
rect 0 8670 18585 8674
rect 62092 8671 64102 8672
rect 0 8618 18467 8670
rect 18519 8618 18585 8670
rect 0 8613 18585 8618
rect 42947 8667 64102 8671
rect 42947 8615 43013 8667
rect 43065 8615 64102 8667
rect 0 8612 490 8613
rect 42947 8610 64102 8615
rect 0 8529 20492 8532
rect 62092 8529 64102 8530
rect 0 8477 20352 8529
rect 20404 8477 20492 8529
rect 0 8471 20492 8477
rect 41040 8526 64102 8529
rect 41040 8474 41128 8526
rect 41180 8474 64102 8526
rect 0 8470 490 8471
rect 41040 8468 64102 8474
rect 0 8386 22342 8390
rect 62092 8387 64102 8388
rect 0 8334 22243 8386
rect 22295 8334 22342 8386
rect 0 8329 22342 8334
rect 39190 8383 64102 8387
rect 39190 8331 39237 8383
rect 39289 8331 64102 8383
rect 0 8328 490 8329
rect 39190 8326 64102 8331
rect 0 8243 24217 8248
rect 62092 8245 64102 8246
rect 0 8191 24133 8243
rect 24185 8191 24217 8243
rect 0 8187 24217 8191
rect 37315 8240 64102 8245
rect 37315 8188 37347 8240
rect 37399 8188 64102 8240
rect 0 8186 490 8187
rect 37315 8184 64102 8188
rect 0 8099 26114 8106
rect 62092 8103 64102 8104
rect 0 8047 26016 8099
rect 26068 8047 26114 8099
rect 0 8045 26114 8047
rect 35418 8096 64102 8103
rect 0 8044 490 8045
rect 35418 8044 35464 8096
rect 35516 8044 64102 8096
rect 35418 8042 64102 8044
rect 0 7957 28044 7964
rect 62092 7961 64102 7962
rect 0 7905 27906 7957
rect 27958 7905 28044 7957
rect 0 7903 28044 7905
rect 33488 7954 64102 7961
rect 0 7902 490 7903
rect 33488 7902 33574 7954
rect 33626 7902 64102 7954
rect 33488 7900 64102 7902
rect 0 7817 29894 7822
rect 62092 7819 64102 7820
rect 0 7765 29798 7817
rect 29850 7765 29894 7817
rect 0 7761 29894 7765
rect 31638 7814 64102 7819
rect 31638 7762 31682 7814
rect 31734 7762 64102 7814
rect 0 7760 490 7761
rect 31638 7758 64102 7762
rect 478 6588 1396 6609
rect 478 6536 492 6588
rect 544 6536 1334 6588
rect 1386 6536 1396 6588
rect 478 6516 1396 6536
rect 622 6112 1403 6127
rect 622 6104 1344 6112
rect 622 6052 639 6104
rect 691 6060 1344 6104
rect 1396 6060 1403 6112
rect 691 6052 1403 6060
rect 622 6034 1403 6052
<< via1 >>
rect 31085 15452 31137 15504
rect 31202 15452 31254 15504
rect 31319 15452 31371 15504
rect 357 13835 409 13887
rect 1175 13839 1227 13891
rect 214 13346 266 13398
rect 1172 13360 1224 13412
rect 29568 12167 29620 12219
rect 31455 12164 31507 12216
rect 27680 12025 27732 12077
rect 33343 12022 33395 12074
rect 25793 11884 25845 11936
rect 35230 11881 35282 11933
rect 23904 11743 23956 11795
rect 37119 11740 37171 11792
rect 22016 11600 22068 11652
rect 39007 11597 39059 11649
rect 20126 11457 20178 11509
rect 40897 11454 40949 11506
rect 18240 11316 18292 11368
rect 42783 11313 42835 11365
rect 16352 11173 16404 11225
rect 44671 11170 44723 11222
rect 14471 11031 14523 11083
rect 46552 11028 46604 11080
rect 12583 10888 12635 10940
rect 48440 10885 48492 10937
rect 10695 10746 10747 10798
rect 50328 10743 50380 10795
rect 8808 10604 8860 10656
rect 52215 10601 52267 10653
rect 6918 10463 6970 10515
rect 54105 10460 54157 10512
rect 5031 10321 5083 10373
rect 55992 10318 56044 10370
rect 3142 10178 3194 10230
rect 57881 10175 57933 10227
rect 1254 10037 1306 10089
rect 59769 10034 59821 10086
rect 32152 9891 32204 9943
rect 32282 9891 32334 9943
rect 32412 9891 32464 9943
rect 59999 9892 60051 9944
rect 3368 9756 3420 9808
rect 5257 9611 5309 9663
rect 7699 9588 7751 9640
rect 7797 9588 7849 9640
rect 31049 9708 31101 9760
rect 31152 9708 31204 9760
rect 31255 9708 31307 9760
rect 31358 9708 31410 9760
rect 58112 9753 58164 9805
rect 56223 9608 56275 9660
rect 7146 9470 7198 9522
rect 54334 9467 54386 9519
rect 9033 9326 9085 9378
rect 32142 9361 32194 9413
rect 32255 9361 32307 9413
rect 32368 9361 32420 9413
rect 32481 9361 32533 9413
rect 32594 9361 32646 9413
rect 52447 9323 52499 9375
rect 10921 9185 10973 9237
rect 50559 9182 50611 9234
rect 12810 9043 12862 9095
rect 48670 9040 48722 9092
rect 14698 8898 14750 8950
rect 46782 8895 46834 8947
rect 16576 8759 16628 8811
rect 44904 8756 44956 8808
rect 18467 8618 18519 8670
rect 43013 8615 43065 8667
rect 20352 8477 20404 8529
rect 41128 8474 41180 8526
rect 22243 8334 22295 8386
rect 39237 8331 39289 8383
rect 24133 8191 24185 8243
rect 37347 8188 37399 8240
rect 26016 8047 26068 8099
rect 35464 8044 35516 8096
rect 27906 7905 27958 7957
rect 33574 7902 33626 7954
rect 29798 7765 29850 7817
rect 31682 7762 31734 7814
rect 32142 7472 32194 7524
rect 32255 7472 32307 7524
rect 32368 7472 32420 7524
rect 32481 7472 32533 7524
rect 32594 7472 32646 7524
rect 32142 7367 32194 7419
rect 32255 7367 32307 7419
rect 32368 7367 32420 7419
rect 32481 7367 32533 7419
rect 32594 7367 32646 7419
rect 492 6536 544 6588
rect 1334 6536 1386 6588
rect 639 6052 691 6104
rect 1344 6060 1396 6112
rect 31074 3223 31126 3275
rect 31157 3223 31209 3275
rect 31240 3223 31292 3275
rect 31323 3223 31375 3275
<< metal2 >>
rect 2628 19017 2672 20184
rect 4516 19017 4560 19992
rect 6404 19017 6448 19992
rect 8292 19017 8336 19992
rect 10180 19017 10224 19992
rect 12068 19017 12112 19992
rect 13956 19017 14000 19992
rect 15844 19017 15888 19992
rect 17732 19017 17776 19992
rect 19620 19017 19664 19992
rect 21508 19017 21552 19992
rect 23396 19017 23440 19992
rect 25284 19017 25328 19992
rect 27172 19017 27216 19992
rect 29060 19017 29104 19992
rect 30948 19017 30992 19992
rect 32836 19017 32880 19992
rect 34724 19017 34768 19992
rect 36612 19017 36656 19992
rect 38500 19017 38544 19992
rect 40388 19017 40432 19992
rect 42276 19017 42320 19992
rect 44164 19017 44208 19992
rect 46052 19017 46096 19992
rect 47940 19017 47984 19992
rect 49828 19017 49872 20151
rect 51716 19017 51760 19992
rect 53604 19017 53648 19992
rect 55492 19017 55536 19992
rect 57380 19017 57424 19992
rect 59268 19017 59312 19992
rect 61156 19017 61200 19992
rect 63982 18814 64095 18836
rect 488 18772 896 18804
rect 61100 18778 64095 18814
rect 326 13887 448 13916
rect 326 13835 357 13887
rect 409 13835 448 13887
rect 326 13807 448 13835
rect 198 13398 284 13418
rect 198 13346 214 13398
rect 266 13346 284 13398
rect 198 13338 284 13346
rect 219 1170 257 13338
rect 373 1650 409 13807
rect 488 6606 520 18772
rect 63730 18335 63843 18364
rect 630 18294 866 18326
rect 61020 18299 63843 18335
rect 478 6588 572 6606
rect 478 6536 492 6588
rect 544 6536 572 6588
rect 478 6512 572 6536
rect 630 6127 666 18294
rect 31021 15559 31417 15588
rect 31021 15503 31052 15559
rect 31108 15504 31161 15559
rect 31217 15504 31270 15559
rect 31326 15504 31417 15559
rect 31137 15503 31161 15504
rect 31254 15503 31270 15504
rect 31021 15457 31085 15503
rect 31137 15457 31202 15503
rect 31254 15457 31319 15503
rect 31021 15401 31052 15457
rect 31137 15452 31161 15457
rect 31254 15452 31270 15457
rect 31371 15452 31417 15504
rect 31108 15401 31161 15452
rect 31217 15401 31270 15452
rect 31326 15401 31417 15452
rect 31021 15380 31417 15401
rect 61286 14735 62528 14923
rect 61818 14478 62528 14735
rect 61295 14463 62528 14478
rect 61295 14369 62527 14463
rect 1162 13891 1266 13914
rect 1162 13839 1175 13891
rect 1227 13879 1266 13891
rect 63730 13879 63843 18299
rect 1227 13843 1438 13879
rect 61114 13843 61731 13879
rect 63465 13843 63843 13879
rect 1227 13839 1266 13843
rect 1162 13814 1266 13839
rect 1142 13412 1246 13440
rect 1142 13360 1172 13412
rect 1224 13405 1246 13412
rect 1224 13360 1327 13405
rect 63982 13396 64095 18778
rect 63504 13360 64095 13396
rect 1142 13343 1327 13360
rect 63982 13358 64095 13360
rect 1142 13336 1246 13343
rect 1258 10099 1302 13161
rect 3146 10242 3190 13161
rect 5034 10382 5078 13161
rect 6922 10526 6966 13161
rect 8810 10666 8854 13161
rect 10698 10808 10742 12753
rect 12586 10950 12630 12773
rect 14474 11092 14518 12763
rect 16356 11233 16400 12770
rect 18244 11374 18288 12823
rect 20132 11519 20176 12763
rect 22020 11662 22064 12743
rect 23908 11804 23952 12743
rect 25796 11945 25840 12703
rect 27684 12088 27728 12747
rect 29572 12234 29616 12757
rect 29549 12219 29643 12234
rect 31459 12231 31503 12596
rect 29549 12167 29568 12219
rect 29620 12167 29643 12219
rect 29549 12153 29643 12167
rect 31432 12216 31526 12231
rect 31432 12164 31455 12216
rect 31507 12164 31526 12216
rect 29572 12109 29616 12153
rect 31432 12150 31526 12164
rect 31459 12106 31503 12150
rect 27669 12077 27746 12088
rect 33347 12085 33391 12617
rect 27669 12025 27680 12077
rect 27732 12025 27746 12077
rect 27669 12015 27746 12025
rect 33329 12074 33406 12085
rect 33329 12022 33343 12074
rect 33395 12022 33406 12074
rect 27684 11972 27728 12015
rect 33329 12012 33406 12022
rect 33347 11969 33391 12012
rect 25780 11936 25857 11945
rect 35235 11942 35279 12673
rect 25780 11884 25793 11936
rect 25845 11884 25857 11936
rect 25780 11872 25857 11884
rect 35218 11933 35295 11942
rect 35218 11881 35230 11933
rect 35282 11881 35295 11933
rect 25796 11842 25840 11872
rect 35218 11869 35295 11881
rect 35235 11839 35279 11869
rect 23893 11795 23970 11804
rect 37123 11801 37167 12598
rect 23893 11743 23904 11795
rect 23956 11743 23970 11795
rect 23893 11731 23970 11743
rect 37105 11792 37182 11801
rect 37105 11740 37119 11792
rect 37171 11740 37182 11792
rect 23908 11695 23952 11731
rect 37105 11728 37182 11740
rect 37123 11692 37167 11728
rect 22004 11652 22081 11662
rect 39011 11659 39055 12608
rect 22004 11600 22016 11652
rect 22068 11600 22081 11652
rect 22004 11589 22081 11600
rect 38994 11649 39071 11659
rect 38994 11597 39007 11649
rect 39059 11597 39071 11649
rect 22020 11555 22064 11589
rect 38994 11586 39071 11597
rect 39011 11552 39055 11586
rect 20118 11509 20195 11519
rect 40899 11516 40943 12636
rect 20118 11457 20126 11509
rect 20178 11457 20195 11509
rect 20118 11446 20195 11457
rect 40880 11506 40957 11516
rect 40880 11454 40897 11506
rect 40949 11454 40957 11506
rect 20132 11404 20176 11446
rect 40880 11443 40957 11454
rect 40899 11401 40943 11443
rect 18227 11368 18304 11374
rect 42787 11371 42831 12629
rect 18227 11316 18240 11368
rect 18292 11316 18304 11368
rect 18227 11301 18304 11316
rect 42771 11365 42848 11371
rect 42771 11313 42783 11365
rect 42835 11313 42848 11365
rect 18244 11258 18288 11301
rect 42771 11298 42848 11313
rect 42787 11255 42831 11298
rect 16340 11225 16417 11233
rect 44675 11230 44719 12627
rect 16340 11173 16352 11225
rect 16404 11173 16417 11225
rect 16340 11160 16417 11173
rect 44658 11222 44735 11230
rect 44658 11170 44671 11222
rect 44723 11170 44735 11222
rect 16356 11131 16400 11160
rect 44658 11157 44735 11170
rect 44675 11128 44719 11157
rect 14459 11083 14536 11092
rect 46557 11089 46601 12595
rect 14459 11031 14471 11083
rect 14523 11031 14536 11083
rect 14459 11019 14536 11031
rect 46539 11080 46616 11089
rect 46539 11028 46552 11080
rect 46604 11028 46616 11080
rect 14474 10991 14518 11019
rect 46539 11016 46616 11028
rect 46557 10988 46601 11016
rect 12571 10940 12648 10950
rect 48445 10947 48489 12633
rect 12571 10888 12583 10940
rect 12635 10888 12648 10940
rect 12571 10877 12648 10888
rect 48427 10937 48504 10947
rect 48427 10885 48440 10937
rect 48492 10885 48504 10937
rect 12586 10854 12630 10877
rect 48427 10874 48504 10885
rect 48445 10851 48489 10874
rect 10682 10798 10759 10808
rect 50333 10805 50377 12618
rect 10682 10746 10695 10798
rect 10747 10746 10759 10798
rect 10682 10735 10759 10746
rect 50316 10795 50393 10805
rect 50316 10743 50328 10795
rect 50380 10743 50393 10795
rect 10698 10697 10742 10735
rect 50316 10732 50393 10743
rect 50333 10694 50377 10732
rect 8796 10656 8873 10666
rect 52221 10663 52265 12618
rect 8796 10604 8808 10656
rect 8860 10604 8873 10656
rect 8796 10593 8873 10604
rect 52202 10653 52279 10663
rect 52202 10601 52215 10653
rect 52267 10601 52279 10653
rect 8810 10560 8854 10593
rect 52202 10590 52279 10601
rect 52221 10557 52265 10590
rect 6908 10515 6985 10526
rect 54109 10523 54153 12631
rect 6908 10463 6918 10515
rect 6970 10463 6985 10515
rect 6908 10453 6985 10463
rect 54090 10512 54167 10523
rect 54090 10460 54105 10512
rect 54157 10460 54167 10512
rect 6922 10417 6966 10453
rect 54090 10450 54167 10460
rect 5018 10373 5095 10382
rect 5018 10321 5031 10373
rect 5083 10321 5095 10373
rect 5018 10309 5095 10321
rect 31022 10377 31419 10416
rect 54109 10414 54153 10450
rect 55997 10379 56041 12648
rect 31022 10321 31045 10377
rect 31101 10321 31149 10377
rect 31205 10321 31253 10377
rect 31309 10321 31357 10377
rect 31413 10321 31419 10377
rect 5034 10270 5078 10309
rect 31022 10278 31419 10321
rect 55980 10370 56057 10379
rect 55980 10318 55992 10370
rect 56044 10318 56057 10370
rect 55980 10306 56057 10318
rect 3134 10230 3211 10242
rect 3134 10178 3142 10230
rect 3194 10178 3211 10230
rect 3134 10169 3211 10178
rect 31022 10222 31045 10278
rect 31101 10222 31149 10278
rect 31205 10222 31253 10278
rect 31309 10222 31357 10278
rect 31413 10222 31419 10278
rect 55997 10267 56041 10306
rect 57885 10239 57929 12646
rect 3146 10133 3190 10169
rect 1241 10089 1318 10099
rect 1241 10037 1254 10089
rect 1306 10037 1318 10089
rect 1241 10026 1318 10037
rect 1258 10003 1302 10026
rect 3375 9817 3419 9861
rect 3356 9808 3435 9817
rect 3356 9756 3368 9808
rect 3420 9756 3435 9808
rect 3356 9741 3435 9756
rect 31022 9760 31419 10222
rect 57864 10227 57941 10239
rect 57864 10175 57881 10227
rect 57933 10175 57941 10227
rect 57864 10166 57941 10175
rect 57885 10130 57929 10166
rect 59773 10096 59817 12644
rect 61662 12036 61706 12762
rect 61612 12006 61760 12036
rect 61612 11950 61655 12006
rect 61711 11950 61760 12006
rect 61612 11934 61760 11950
rect 59757 10086 59834 10096
rect 59757 10034 59769 10086
rect 59821 10034 59834 10086
rect 59757 10023 59834 10034
rect 59773 10000 59817 10023
rect 32113 9947 32514 9972
rect 60001 9955 60045 9985
rect 32113 9891 32152 9947
rect 32208 9891 32281 9947
rect 32337 9891 32410 9947
rect 32466 9891 32514 9947
rect 32113 9878 32514 9891
rect 59983 9944 60062 9955
rect 59983 9892 59999 9944
rect 60051 9892 60062 9944
rect 59983 9879 60062 9892
rect 58113 9814 58157 9858
rect 3375 7204 3419 9741
rect 5263 9671 5307 9744
rect 31022 9708 31049 9760
rect 31101 9708 31152 9760
rect 31204 9708 31255 9760
rect 31307 9708 31358 9760
rect 31410 9708 31419 9760
rect 58097 9805 58176 9814
rect 58097 9753 58112 9805
rect 58164 9753 58176 9805
rect 5238 9663 5317 9671
rect 5238 9611 5257 9663
rect 5309 9611 5317 9663
rect 5238 9595 5317 9611
rect 7610 9644 7957 9674
rect 7610 9640 7700 9644
rect 5263 7167 5307 9595
rect 7151 9530 7195 9604
rect 7610 9588 7699 9640
rect 7756 9588 7797 9644
rect 7853 9588 7957 9644
rect 7610 9550 7957 9588
rect 7133 9522 7212 9530
rect 7133 9470 7146 9522
rect 7198 9470 7212 9522
rect 7133 9454 7212 9470
rect 7151 7216 7195 9454
rect 9039 9389 9083 9438
rect 9022 9378 9101 9389
rect 9022 9326 9033 9378
rect 9085 9326 9101 9378
rect 9022 9313 9101 9326
rect 9039 7253 9083 9313
rect 10927 9247 10971 9292
rect 10910 9237 10989 9247
rect 10910 9185 10921 9237
rect 10973 9185 10989 9237
rect 10910 9171 10989 9185
rect 10927 7216 10971 9171
rect 12815 9104 12859 9145
rect 12799 9095 12878 9104
rect 12799 9043 12810 9095
rect 12862 9043 12878 9095
rect 12799 9028 12878 9043
rect 31022 9048 31419 9708
rect 56225 9668 56269 9741
rect 58097 9738 58176 9753
rect 56215 9660 56294 9668
rect 56215 9608 56223 9660
rect 56275 9608 56294 9660
rect 54337 9527 54381 9601
rect 56215 9592 56294 9608
rect 54320 9519 54399 9527
rect 54320 9467 54334 9519
rect 54386 9467 54399 9519
rect 54320 9451 54399 9467
rect 12815 7192 12859 9028
rect 31022 8992 31058 9048
rect 31114 8992 31146 9048
rect 31202 8992 31234 9048
rect 31290 8992 31322 9048
rect 31378 8992 31419 9048
rect 14703 8959 14747 8986
rect 14687 8950 14766 8959
rect 14687 8898 14698 8950
rect 14750 8898 14766 8950
rect 14687 8883 14766 8898
rect 31022 8953 31419 8992
rect 31022 8897 31058 8953
rect 31114 8897 31146 8953
rect 31202 8897 31234 8953
rect 31290 8897 31322 8953
rect 31378 8897 31419 8953
rect 14703 7216 14747 8883
rect 31022 8866 31419 8897
rect 32087 9413 32754 9430
rect 32087 9361 32142 9413
rect 32194 9361 32255 9413
rect 32307 9361 32368 9413
rect 32420 9361 32481 9413
rect 32533 9361 32594 9413
rect 32646 9361 32754 9413
rect 52449 9386 52493 9435
rect 16585 8821 16629 8863
rect 16565 8811 16644 8821
rect 16565 8759 16576 8811
rect 16628 8759 16644 8811
rect 16565 8745 16644 8759
rect 16585 7161 16629 8745
rect 18473 8679 18517 8735
rect 18455 8670 18534 8679
rect 18455 8618 18467 8670
rect 18519 8618 18534 8670
rect 18455 8603 18534 8618
rect 18473 7192 18517 8603
rect 20361 8538 20405 8594
rect 20341 8529 20420 8538
rect 20341 8477 20352 8529
rect 20404 8477 20420 8529
rect 20341 8462 20420 8477
rect 20361 7234 20405 8462
rect 22249 8396 22293 8453
rect 22231 8386 22310 8396
rect 22231 8334 22243 8386
rect 22295 8334 22310 8386
rect 22231 8320 22310 8334
rect 22249 7210 22293 8320
rect 24137 8253 24181 8319
rect 24121 8243 24200 8253
rect 24121 8191 24133 8243
rect 24185 8191 24200 8243
rect 24121 8177 24200 8191
rect 24137 7161 24181 8177
rect 26025 8112 26069 8166
rect 26003 8099 26082 8112
rect 26003 8047 26016 8099
rect 26068 8047 26082 8099
rect 26003 8036 26082 8047
rect 26025 7192 26069 8036
rect 27913 7970 27957 8007
rect 27897 7957 27976 7970
rect 27897 7905 27906 7957
rect 27958 7905 27976 7957
rect 27897 7894 27976 7905
rect 27913 7192 27957 7894
rect 29801 7828 29845 7903
rect 29787 7817 29866 7828
rect 31687 7825 31731 7900
rect 29787 7765 29798 7817
rect 29850 7765 29866 7817
rect 29787 7752 29866 7765
rect 31666 7814 31745 7825
rect 31666 7762 31682 7814
rect 31734 7762 31745 7814
rect 29801 7198 29845 7752
rect 31666 7749 31745 7762
rect 31687 7293 31731 7749
rect 32087 7524 32754 9361
rect 52431 9375 52510 9386
rect 52431 9323 52447 9375
rect 52499 9323 52510 9375
rect 52431 9310 52510 9323
rect 50561 9244 50605 9289
rect 50543 9234 50622 9244
rect 50543 9182 50559 9234
rect 50611 9182 50622 9234
rect 50543 9168 50622 9182
rect 48673 9101 48717 9142
rect 48654 9092 48733 9101
rect 48654 9040 48670 9092
rect 48722 9040 48733 9092
rect 48654 9025 48733 9040
rect 46785 8956 46829 8983
rect 46766 8947 46845 8956
rect 46766 8895 46782 8947
rect 46834 8895 46845 8947
rect 46766 8880 46845 8895
rect 44903 8818 44947 8860
rect 44888 8808 44967 8818
rect 44888 8756 44904 8808
rect 44956 8756 44967 8808
rect 44888 8742 44967 8756
rect 43015 8676 43059 8732
rect 42998 8667 43077 8676
rect 42998 8615 43013 8667
rect 43065 8615 43077 8667
rect 42998 8600 43077 8615
rect 41127 8535 41171 8591
rect 41112 8526 41191 8535
rect 41112 8474 41128 8526
rect 41180 8474 41191 8526
rect 41112 8459 41191 8474
rect 39239 8393 39283 8450
rect 39222 8383 39301 8393
rect 39222 8331 39237 8383
rect 39289 8331 39301 8383
rect 39222 8317 39301 8331
rect 37351 8250 37395 8316
rect 37332 8240 37411 8250
rect 37332 8188 37347 8240
rect 37399 8188 37411 8240
rect 37332 8174 37411 8188
rect 35463 8109 35507 8163
rect 35450 8096 35529 8109
rect 35450 8044 35464 8096
rect 35516 8044 35529 8096
rect 35450 8033 35529 8044
rect 33575 7967 33619 8004
rect 33556 7954 33635 7967
rect 33556 7902 33574 7954
rect 33626 7902 33635 7954
rect 33556 7891 33635 7902
rect 32087 7472 32142 7524
rect 32194 7472 32255 7524
rect 32307 7472 32368 7524
rect 32420 7472 32481 7524
rect 32533 7472 32594 7524
rect 32646 7472 32754 7524
rect 32087 7419 32754 7472
rect 32087 7367 32142 7419
rect 32194 7367 32255 7419
rect 32307 7367 32368 7419
rect 32420 7367 32481 7419
rect 32533 7367 32594 7419
rect 32646 7367 32754 7419
rect 32087 7319 32754 7367
rect 33575 7340 33619 7891
rect 35463 7302 35507 8033
rect 37351 7299 37395 8174
rect 39239 7293 39283 8317
rect 41127 7319 41171 8459
rect 43015 7244 43059 8600
rect 44903 7287 44947 8742
rect 46785 7306 46829 8880
rect 48673 7270 48717 9025
rect 50561 7259 50605 9168
rect 52449 7285 52493 9310
rect 54337 7310 54381 9451
rect 56225 7268 56269 9592
rect 58113 7329 58157 9738
rect 60001 7299 60045 9879
rect 1300 6588 1402 6616
rect 62964 6594 63082 6623
rect 1300 6536 1334 6588
rect 1386 6584 1402 6588
rect 1386 6548 3477 6584
rect 61864 6560 63082 6594
rect 1386 6536 1402 6548
rect 1300 6510 1402 6536
rect 629 6104 740 6127
rect 629 6052 639 6104
rect 691 6052 740 6104
rect 629 6012 740 6052
rect 1337 6112 1407 6133
rect 1337 6060 1344 6112
rect 1396 6104 1407 6112
rect 1396 6068 3436 6104
rect 61848 6068 62762 6102
rect 1396 6060 1407 6068
rect 1337 6029 1407 6060
rect 31022 3324 31419 3357
rect 31022 3268 31063 3324
rect 31119 3275 31155 3324
rect 31211 3275 31247 3324
rect 31303 3275 31339 3324
rect 31126 3268 31155 3275
rect 31211 3268 31240 3275
rect 31303 3268 31323 3275
rect 31395 3268 31419 3324
rect 31022 3233 31074 3268
rect 31126 3233 31157 3268
rect 31209 3233 31240 3268
rect 31292 3233 31323 3268
rect 31375 3233 31419 3268
rect 31022 3177 31063 3233
rect 31126 3223 31155 3233
rect 31211 3223 31240 3233
rect 31303 3223 31323 3233
rect 31119 3177 31155 3223
rect 31211 3177 31247 3223
rect 31303 3177 31339 3223
rect 31395 3177 31419 3233
rect 31022 3151 31419 3177
rect 373 1612 1094 1650
rect 62644 1648 62762 6068
rect 61249 1612 62762 1648
rect 62964 1174 63082 6560
rect 219 1132 1080 1170
rect 61383 1112 63082 1174
rect 62964 1103 63082 1112
rect 2857 0 2913 930
rect 4745 0 4801 930
rect 6633 0 6689 930
rect 8521 0 8577 930
rect 10409 0 10465 930
rect 12297 0 12353 930
rect 14185 0 14241 930
rect 16073 0 16129 930
rect 17961 0 18017 930
rect 19849 0 19905 930
rect 21737 0 21793 930
rect 23625 0 23681 930
rect 25513 0 25569 930
rect 27401 0 27457 930
rect 29289 0 29345 930
rect 31177 0 31233 930
rect 33065 0 33121 930
rect 34953 0 35009 930
rect 36841 0 36897 930
rect 38729 0 38785 930
rect 40617 0 40673 930
rect 42505 0 42561 930
rect 44393 0 44449 930
rect 46281 0 46337 930
rect 48169 0 48225 930
rect 50057 0 50113 930
rect 51945 0 52001 930
rect 53833 0 53889 930
rect 55721 0 55777 930
rect 57609 0 57665 930
rect 59497 0 59553 930
rect 61385 0 61441 930
<< via2 >>
rect 31052 15504 31108 15559
rect 31161 15504 31217 15559
rect 31270 15504 31326 15559
rect 31052 15503 31085 15504
rect 31085 15503 31108 15504
rect 31161 15503 31202 15504
rect 31202 15503 31217 15504
rect 31270 15503 31319 15504
rect 31319 15503 31326 15504
rect 31052 15452 31085 15457
rect 31085 15452 31108 15457
rect 31161 15452 31202 15457
rect 31202 15452 31217 15457
rect 31270 15452 31319 15457
rect 31319 15452 31326 15457
rect 31052 15401 31108 15452
rect 31161 15401 31217 15452
rect 31270 15401 31326 15452
rect 31045 10321 31101 10377
rect 31149 10321 31205 10377
rect 31253 10321 31309 10377
rect 31357 10321 31413 10377
rect 31045 10222 31101 10278
rect 31149 10222 31205 10278
rect 31253 10222 31309 10278
rect 31357 10222 31413 10278
rect 61655 11950 61711 12006
rect 32152 9943 32208 9947
rect 32152 9891 32204 9943
rect 32204 9891 32208 9943
rect 32281 9943 32337 9947
rect 32281 9891 32282 9943
rect 32282 9891 32334 9943
rect 32334 9891 32337 9943
rect 32410 9943 32466 9947
rect 32410 9891 32412 9943
rect 32412 9891 32464 9943
rect 32464 9891 32466 9943
rect 7700 9640 7756 9644
rect 7700 9588 7751 9640
rect 7751 9588 7756 9640
rect 7797 9640 7853 9644
rect 7797 9588 7849 9640
rect 7849 9588 7853 9640
rect 31058 8992 31114 9048
rect 31146 8992 31202 9048
rect 31234 8992 31290 9048
rect 31322 8992 31378 9048
rect 31058 8897 31114 8953
rect 31146 8897 31202 8953
rect 31234 8897 31290 8953
rect 31322 8897 31378 8953
rect 31063 3275 31119 3324
rect 31155 3275 31211 3324
rect 31247 3275 31303 3324
rect 31339 3275 31395 3324
rect 31063 3268 31074 3275
rect 31074 3268 31119 3275
rect 31155 3268 31157 3275
rect 31157 3268 31209 3275
rect 31209 3268 31211 3275
rect 31247 3268 31292 3275
rect 31292 3268 31303 3275
rect 31339 3268 31375 3275
rect 31375 3268 31395 3275
rect 31063 3223 31074 3233
rect 31074 3223 31119 3233
rect 31155 3223 31157 3233
rect 31157 3223 31209 3233
rect 31209 3223 31211 3233
rect 31247 3223 31292 3233
rect 31292 3223 31303 3233
rect 31339 3223 31375 3233
rect 31375 3223 31395 3233
rect 31063 3177 31119 3223
rect 31155 3177 31211 3223
rect 31247 3177 31303 3223
rect 31339 3177 31395 3223
<< metal3 >>
rect 20583 19764 20689 19781
rect 20583 19700 20604 19764
rect 20668 19700 20689 19764
rect 20583 19684 20689 19700
rect 20583 19620 20604 19684
rect 20668 19620 20689 19684
rect 20583 19603 20689 19620
rect 20757 19764 20863 19781
rect 20757 19700 20778 19764
rect 20842 19700 20863 19764
rect 20757 19684 20863 19700
rect 20757 19620 20778 19684
rect 20842 19620 20863 19684
rect 20757 19603 20863 19620
rect 20931 19764 21037 19781
rect 20931 19700 20952 19764
rect 21016 19700 21037 19764
rect 20931 19684 21037 19700
rect 20931 19620 20952 19684
rect 21016 19620 21037 19684
rect 20931 19603 21037 19620
rect 35558 19741 35664 19758
rect 35558 19677 35579 19741
rect 35643 19677 35664 19741
rect 35558 19661 35664 19677
rect 35558 19597 35579 19661
rect 35643 19597 35664 19661
rect 35558 19580 35664 19597
rect 35741 19741 35847 19758
rect 35741 19677 35762 19741
rect 35826 19677 35847 19741
rect 35741 19661 35847 19677
rect 35741 19597 35762 19661
rect 35826 19597 35847 19661
rect 35741 19580 35847 19597
rect 35924 19741 36030 19758
rect 35924 19677 35945 19741
rect 36009 19677 36030 19741
rect 35924 19661 36030 19677
rect 35924 19597 35945 19661
rect 36009 19597 36030 19661
rect 35924 19580 36030 19597
rect 51056 19754 51162 19771
rect 51056 19690 51077 19754
rect 51141 19690 51162 19754
rect 51056 19674 51162 19690
rect 51056 19610 51077 19674
rect 51141 19610 51162 19674
rect 51056 19593 51162 19610
rect 51239 19754 51345 19771
rect 51239 19690 51260 19754
rect 51324 19690 51345 19754
rect 51239 19674 51345 19690
rect 51239 19610 51260 19674
rect 51324 19610 51345 19674
rect 51239 19593 51345 19610
rect 51422 19754 51528 19771
rect 51422 19690 51443 19754
rect 51507 19690 51528 19754
rect 51422 19674 51528 19690
rect 51422 19610 51443 19674
rect 51507 19610 51528 19674
rect 51422 19593 51528 19610
rect 19060 17620 19166 17637
rect 19060 17556 19081 17620
rect 19145 17556 19166 17620
rect 19060 17540 19166 17556
rect 19060 17476 19081 17540
rect 19145 17476 19166 17540
rect 19060 17459 19166 17476
rect 19234 17620 19340 17637
rect 19234 17556 19255 17620
rect 19319 17556 19340 17620
rect 19234 17540 19340 17556
rect 19234 17476 19255 17540
rect 19319 17476 19340 17540
rect 19234 17459 19340 17476
rect 19408 17620 19514 17637
rect 19408 17556 19429 17620
rect 19493 17556 19514 17620
rect 19408 17540 19514 17556
rect 19408 17476 19429 17540
rect 19493 17476 19514 17540
rect 19408 17459 19514 17476
rect 34037 17625 34143 17642
rect 34037 17561 34058 17625
rect 34122 17561 34143 17625
rect 34037 17545 34143 17561
rect 34037 17481 34058 17545
rect 34122 17481 34143 17545
rect 34037 17464 34143 17481
rect 34220 17625 34326 17642
rect 34220 17561 34241 17625
rect 34305 17561 34326 17625
rect 34220 17545 34326 17561
rect 34220 17481 34241 17545
rect 34305 17481 34326 17545
rect 34220 17464 34326 17481
rect 34403 17625 34509 17642
rect 34403 17561 34424 17625
rect 34488 17561 34509 17625
rect 34403 17545 34509 17561
rect 34403 17481 34424 17545
rect 34488 17481 34509 17545
rect 34403 17464 34509 17481
rect 49531 17616 49637 17633
rect 49531 17552 49552 17616
rect 49616 17552 49637 17616
rect 49531 17536 49637 17552
rect 49531 17472 49552 17536
rect 49616 17472 49637 17536
rect 49531 17455 49637 17472
rect 49714 17616 49820 17633
rect 49714 17552 49735 17616
rect 49799 17552 49820 17616
rect 49714 17536 49820 17552
rect 49714 17472 49735 17536
rect 49799 17472 49820 17536
rect 49714 17455 49820 17472
rect 49897 17616 50003 17633
rect 49897 17552 49918 17616
rect 49982 17552 50003 17616
rect 49897 17536 50003 17552
rect 49897 17472 49918 17536
rect 49982 17472 50003 17536
rect 49897 17455 50003 17472
rect 31021 15559 31416 15588
rect 31021 15503 31052 15559
rect 31108 15514 31161 15559
rect 31108 15503 31111 15514
rect 31217 15503 31270 15559
rect 31326 15503 31416 15559
rect 31021 15457 31111 15503
rect 31175 15457 31416 15503
rect 31021 15401 31052 15457
rect 31108 15450 31111 15457
rect 31108 15401 31161 15450
rect 31217 15401 31270 15457
rect 31326 15401 31416 15457
rect 31021 15380 31416 15401
rect 19073 14692 19179 14709
rect 19073 14628 19094 14692
rect 19158 14628 19179 14692
rect 19073 14612 19179 14628
rect 19073 14548 19094 14612
rect 19158 14548 19179 14612
rect 19073 14531 19179 14548
rect 19247 14692 19353 14709
rect 19247 14628 19268 14692
rect 19332 14628 19353 14692
rect 19247 14612 19353 14628
rect 19247 14548 19268 14612
rect 19332 14548 19353 14612
rect 19247 14531 19353 14548
rect 19421 14692 19527 14709
rect 19421 14628 19442 14692
rect 19506 14628 19527 14692
rect 19421 14612 19527 14628
rect 19421 14548 19442 14612
rect 19506 14548 19527 14612
rect 19421 14531 19527 14548
rect 32158 14689 32282 14700
rect 32158 14625 32188 14689
rect 32252 14625 32282 14689
rect 32158 14609 32282 14625
rect 32158 14545 32188 14609
rect 32252 14545 32282 14609
rect 32158 14534 32282 14545
rect 32357 14689 32481 14700
rect 32357 14625 32387 14689
rect 32451 14625 32481 14689
rect 32357 14609 32481 14625
rect 32357 14545 32387 14609
rect 32451 14545 32481 14609
rect 32357 14534 32481 14545
rect 34023 14690 34129 14707
rect 34023 14626 34044 14690
rect 34108 14626 34129 14690
rect 34023 14610 34129 14626
rect 34023 14546 34044 14610
rect 34108 14546 34129 14610
rect 34023 14529 34129 14546
rect 34206 14690 34312 14707
rect 34206 14626 34227 14690
rect 34291 14626 34312 14690
rect 34206 14610 34312 14626
rect 34206 14546 34227 14610
rect 34291 14546 34312 14610
rect 34206 14529 34312 14546
rect 34389 14690 34495 14707
rect 34389 14626 34410 14690
rect 34474 14626 34495 14690
rect 34389 14610 34495 14626
rect 34389 14546 34410 14610
rect 34474 14546 34495 14610
rect 34389 14529 34495 14546
rect 49562 14687 49668 14704
rect 49562 14623 49583 14687
rect 49647 14623 49668 14687
rect 49562 14607 49668 14623
rect 49562 14543 49583 14607
rect 49647 14543 49668 14607
rect 49562 14526 49668 14543
rect 49745 14687 49851 14704
rect 49745 14623 49766 14687
rect 49830 14623 49851 14687
rect 49745 14607 49851 14623
rect 49745 14543 49766 14607
rect 49830 14543 49851 14607
rect 49745 14526 49851 14543
rect 49928 14687 50034 14704
rect 49928 14623 49949 14687
rect 50013 14623 50034 14687
rect 49928 14607 50034 14623
rect 49928 14543 49949 14607
rect 50013 14543 50034 14607
rect 49928 14526 50034 14543
rect 20583 12556 20689 12573
rect 20583 12492 20604 12556
rect 20668 12492 20689 12556
rect 20583 12476 20689 12492
rect 20583 12412 20604 12476
rect 20668 12412 20689 12476
rect 20583 12395 20689 12412
rect 20757 12556 20863 12573
rect 20757 12492 20778 12556
rect 20842 12492 20863 12556
rect 20757 12476 20863 12492
rect 20757 12412 20778 12476
rect 20842 12412 20863 12476
rect 20757 12395 20863 12412
rect 20931 12556 21037 12573
rect 20931 12492 20952 12556
rect 21016 12492 21037 12556
rect 20931 12476 21037 12492
rect 20931 12412 20952 12476
rect 21016 12412 21037 12476
rect 20931 12395 21037 12412
rect 35573 12567 35679 12584
rect 35573 12503 35594 12567
rect 35658 12503 35679 12567
rect 35573 12487 35679 12503
rect 35573 12423 35594 12487
rect 35658 12423 35679 12487
rect 35573 12406 35679 12423
rect 35756 12567 35862 12584
rect 35756 12503 35777 12567
rect 35841 12503 35862 12567
rect 35756 12487 35862 12503
rect 35756 12423 35777 12487
rect 35841 12423 35862 12487
rect 35756 12406 35862 12423
rect 35939 12567 36045 12584
rect 35939 12503 35960 12567
rect 36024 12503 36045 12567
rect 35939 12487 36045 12503
rect 35939 12423 35960 12487
rect 36024 12423 36045 12487
rect 35939 12406 36045 12423
rect 51031 12558 51137 12575
rect 51031 12494 51052 12558
rect 51116 12494 51137 12558
rect 51031 12478 51137 12494
rect 51031 12414 51052 12478
rect 51116 12414 51137 12478
rect 51031 12397 51137 12414
rect 51214 12558 51320 12575
rect 51214 12494 51235 12558
rect 51299 12494 51320 12558
rect 51214 12478 51320 12494
rect 51214 12414 51235 12478
rect 51299 12414 51320 12478
rect 51214 12397 51320 12414
rect 51397 12558 51503 12575
rect 51397 12494 51418 12558
rect 51482 12494 51503 12558
rect 51397 12478 51503 12494
rect 51397 12414 51418 12478
rect 51482 12414 51503 12478
rect 51397 12397 51503 12414
rect 61612 12006 64105 12036
rect 61612 11950 61655 12006
rect 61711 11950 64105 12006
rect 61612 11938 64105 11950
rect 31021 10377 31418 10419
rect 31021 10321 31045 10377
rect 31101 10330 31149 10377
rect 31101 10321 31102 10330
rect 31205 10321 31253 10377
rect 31309 10330 31357 10377
rect 31348 10321 31357 10330
rect 31413 10321 31418 10377
rect 31021 10278 31102 10321
rect 31166 10278 31284 10321
rect 31348 10278 31418 10321
rect 31021 10222 31045 10278
rect 31101 10266 31102 10278
rect 31101 10222 31149 10266
rect 31205 10222 31253 10278
rect 31348 10266 31357 10278
rect 31309 10222 31357 10266
rect 31413 10222 31418 10278
rect 31021 10195 31418 10222
rect 32113 9961 32514 9972
rect 32113 9947 32249 9961
rect 32313 9947 32329 9961
rect 32393 9947 32514 9961
rect 32113 9891 32152 9947
rect 32208 9897 32249 9947
rect 32393 9897 32410 9947
rect 32208 9891 32281 9897
rect 32337 9891 32410 9897
rect 32466 9891 32514 9947
rect 32113 9878 32514 9891
rect 7610 9660 7957 9674
rect 509 9644 7957 9660
rect 509 9588 7700 9644
rect 7756 9588 7797 9644
rect 7853 9588 7957 9644
rect 509 9570 7957 9588
rect 7610 9550 7957 9570
rect 31022 9048 31419 9106
rect 31022 8992 31058 9048
rect 31114 9007 31146 9048
rect 31202 8992 31234 9048
rect 31290 9007 31322 9048
rect 31378 8992 31419 9048
rect 31022 8953 31094 8992
rect 31158 8953 31284 8992
rect 31348 8953 31419 8992
rect 31022 8897 31058 8953
rect 31114 8897 31146 8943
rect 31202 8897 31234 8953
rect 31290 8897 31322 8943
rect 31378 8897 31419 8953
rect 31022 8866 31419 8897
rect 3781 7515 3887 7532
rect 3781 7451 3802 7515
rect 3866 7451 3887 7515
rect 3781 7435 3887 7451
rect 3781 7371 3802 7435
rect 3866 7371 3887 7435
rect 3781 7354 3887 7371
rect 4032 7515 4138 7532
rect 4032 7451 4053 7515
rect 4117 7451 4138 7515
rect 4032 7435 4138 7451
rect 4032 7371 4053 7435
rect 4117 7371 4138 7435
rect 4032 7354 4138 7371
rect 4283 7515 4389 7532
rect 4283 7451 4304 7515
rect 4368 7451 4389 7515
rect 4283 7435 4389 7451
rect 4283 7371 4304 7435
rect 4368 7371 4389 7435
rect 4283 7354 4389 7371
rect 20561 7518 20667 7535
rect 20561 7454 20582 7518
rect 20646 7454 20667 7518
rect 20561 7438 20667 7454
rect 20561 7374 20582 7438
rect 20646 7374 20667 7438
rect 20561 7357 20667 7374
rect 20735 7518 20841 7535
rect 20735 7454 20756 7518
rect 20820 7454 20841 7518
rect 20735 7438 20841 7454
rect 20735 7374 20756 7438
rect 20820 7374 20841 7438
rect 20735 7357 20841 7374
rect 20909 7518 21015 7535
rect 20909 7454 20930 7518
rect 20994 7454 21015 7518
rect 20909 7438 21015 7454
rect 20909 7374 20930 7438
rect 20994 7374 21015 7438
rect 20909 7357 21015 7374
rect 35528 7525 35634 7542
rect 35528 7461 35549 7525
rect 35613 7461 35634 7525
rect 35528 7445 35634 7461
rect 35528 7381 35549 7445
rect 35613 7381 35634 7445
rect 35528 7364 35634 7381
rect 35711 7525 35817 7542
rect 35711 7461 35732 7525
rect 35796 7461 35817 7525
rect 35711 7445 35817 7461
rect 35711 7381 35732 7445
rect 35796 7381 35817 7445
rect 35711 7364 35817 7381
rect 35894 7525 36000 7542
rect 35894 7461 35915 7525
rect 35979 7461 36000 7525
rect 35894 7445 36000 7461
rect 35894 7381 35915 7445
rect 35979 7381 36000 7445
rect 35894 7364 36000 7381
rect 51033 7517 51139 7534
rect 51033 7453 51054 7517
rect 51118 7453 51139 7517
rect 51033 7437 51139 7453
rect 51033 7373 51054 7437
rect 51118 7373 51139 7437
rect 51033 7356 51139 7373
rect 51216 7517 51322 7534
rect 51216 7453 51237 7517
rect 51301 7453 51322 7517
rect 51216 7437 51322 7453
rect 51216 7373 51237 7437
rect 51301 7373 51322 7437
rect 51216 7356 51322 7373
rect 51399 7517 51505 7534
rect 51399 7453 51420 7517
rect 51484 7453 51505 7517
rect 51399 7437 51505 7453
rect 51399 7373 51420 7437
rect 51484 7373 51505 7437
rect 51399 7356 51505 7373
rect 2488 5386 3490 5456
rect 2488 5322 2577 5386
rect 2641 5322 2753 5386
rect 2817 5322 2929 5386
rect 2993 5322 3490 5386
rect 2488 5306 3490 5322
rect 2488 5242 2577 5306
rect 2641 5242 2753 5306
rect 2817 5242 2929 5306
rect 2993 5242 3490 5306
rect 2488 5202 3490 5242
rect 19059 5392 19165 5409
rect 19059 5328 19080 5392
rect 19144 5328 19165 5392
rect 19059 5312 19165 5328
rect 19059 5248 19080 5312
rect 19144 5248 19165 5312
rect 19059 5231 19165 5248
rect 19233 5392 19339 5409
rect 19233 5328 19254 5392
rect 19318 5328 19339 5392
rect 19233 5312 19339 5328
rect 19233 5248 19254 5312
rect 19318 5248 19339 5312
rect 19233 5231 19339 5248
rect 19407 5392 19513 5409
rect 19407 5328 19428 5392
rect 19492 5328 19513 5392
rect 19407 5312 19513 5328
rect 19407 5248 19428 5312
rect 19492 5248 19513 5312
rect 19407 5231 19513 5248
rect 34035 5393 34141 5410
rect 34035 5329 34056 5393
rect 34120 5329 34141 5393
rect 34035 5313 34141 5329
rect 34035 5249 34056 5313
rect 34120 5249 34141 5313
rect 34035 5232 34141 5249
rect 34218 5393 34324 5410
rect 34218 5329 34239 5393
rect 34303 5329 34324 5393
rect 34218 5313 34324 5329
rect 34218 5249 34239 5313
rect 34303 5249 34324 5313
rect 34218 5232 34324 5249
rect 34401 5393 34507 5410
rect 34401 5329 34422 5393
rect 34486 5329 34507 5393
rect 34401 5313 34507 5329
rect 34401 5249 34422 5313
rect 34486 5249 34507 5313
rect 34401 5232 34507 5249
rect 49530 5389 49636 5406
rect 49530 5325 49551 5389
rect 49615 5325 49636 5389
rect 49530 5309 49636 5325
rect 49530 5245 49551 5309
rect 49615 5245 49636 5309
rect 49530 5228 49636 5245
rect 49713 5389 49819 5406
rect 49713 5325 49734 5389
rect 49798 5325 49819 5389
rect 49713 5309 49819 5325
rect 49713 5245 49734 5309
rect 49798 5245 49819 5309
rect 49713 5228 49819 5245
rect 49896 5389 50002 5406
rect 49896 5325 49917 5389
rect 49981 5325 50002 5389
rect 49896 5309 50002 5325
rect 49896 5245 49917 5309
rect 49981 5245 50002 5309
rect 49896 5228 50002 5245
rect 31022 3324 31419 3357
rect 31022 3268 31063 3324
rect 31119 3278 31155 3324
rect 31211 3268 31247 3324
rect 31303 3279 31339 3324
rect 31395 3268 31419 3324
rect 31022 3233 31106 3268
rect 31170 3233 31280 3268
rect 31344 3233 31419 3268
rect 31022 3177 31063 3233
rect 31119 3177 31155 3214
rect 31211 3177 31247 3233
rect 31303 3177 31339 3215
rect 31395 3177 31419 3233
rect 31022 3151 31419 3177
rect 2552 2453 2658 2470
rect 2552 2389 2573 2453
rect 2637 2389 2658 2453
rect 2552 2373 2658 2389
rect 2552 2309 2573 2373
rect 2637 2309 2658 2373
rect 2552 2292 2658 2309
rect 2728 2453 2834 2470
rect 2728 2389 2749 2453
rect 2813 2389 2834 2453
rect 2728 2373 2834 2389
rect 2728 2309 2749 2373
rect 2813 2309 2834 2373
rect 2728 2292 2834 2309
rect 2904 2453 3010 2470
rect 2904 2389 2925 2453
rect 2989 2389 3010 2453
rect 2904 2373 3010 2389
rect 2904 2309 2925 2373
rect 2989 2309 3010 2373
rect 2904 2292 3010 2309
rect 19056 2456 19162 2473
rect 19056 2392 19077 2456
rect 19141 2392 19162 2456
rect 19056 2376 19162 2392
rect 19056 2312 19077 2376
rect 19141 2312 19162 2376
rect 19056 2295 19162 2312
rect 19230 2456 19336 2473
rect 19230 2392 19251 2456
rect 19315 2392 19336 2456
rect 19230 2376 19336 2392
rect 19230 2312 19251 2376
rect 19315 2312 19336 2376
rect 19230 2295 19336 2312
rect 19404 2456 19510 2473
rect 19404 2392 19425 2456
rect 19489 2392 19510 2456
rect 19404 2376 19510 2392
rect 19404 2312 19425 2376
rect 19489 2312 19510 2376
rect 19404 2295 19510 2312
rect 34047 2452 34153 2469
rect 34047 2388 34068 2452
rect 34132 2388 34153 2452
rect 34047 2372 34153 2388
rect 34047 2308 34068 2372
rect 34132 2308 34153 2372
rect 34047 2291 34153 2308
rect 34230 2452 34336 2469
rect 34230 2388 34251 2452
rect 34315 2388 34336 2452
rect 34230 2372 34336 2388
rect 34230 2308 34251 2372
rect 34315 2308 34336 2372
rect 34230 2291 34336 2308
rect 34413 2452 34519 2469
rect 34413 2388 34434 2452
rect 34498 2388 34519 2452
rect 34413 2372 34519 2388
rect 34413 2308 34434 2372
rect 34498 2308 34519 2372
rect 34413 2291 34519 2308
rect 49538 2456 49644 2473
rect 49538 2392 49559 2456
rect 49623 2392 49644 2456
rect 49538 2376 49644 2392
rect 49538 2312 49559 2376
rect 49623 2312 49644 2376
rect 49538 2295 49644 2312
rect 49721 2456 49827 2473
rect 49721 2392 49742 2456
rect 49806 2392 49827 2456
rect 49721 2376 49827 2392
rect 49721 2312 49742 2376
rect 49806 2312 49827 2376
rect 49721 2295 49827 2312
rect 49904 2456 50010 2473
rect 49904 2392 49925 2456
rect 49989 2392 50010 2456
rect 49904 2376 50010 2392
rect 49904 2312 49925 2376
rect 49989 2312 50010 2376
rect 49904 2295 50010 2312
rect 3815 331 3921 348
rect 3815 267 3836 331
rect 3900 267 3921 331
rect 3815 251 3921 267
rect 3815 187 3836 251
rect 3900 187 3921 251
rect 3815 170 3921 187
rect 4066 331 4172 348
rect 4066 267 4087 331
rect 4151 267 4172 331
rect 4066 251 4172 267
rect 4066 187 4087 251
rect 4151 187 4172 251
rect 4066 170 4172 187
rect 4317 331 4423 348
rect 4317 267 4338 331
rect 4402 267 4423 331
rect 4317 251 4423 267
rect 4317 187 4338 251
rect 4402 187 4423 251
rect 4317 170 4423 187
rect 20565 334 20671 351
rect 20565 270 20586 334
rect 20650 270 20671 334
rect 20565 254 20671 270
rect 20565 190 20586 254
rect 20650 190 20671 254
rect 20565 173 20671 190
rect 20739 334 20845 351
rect 20739 270 20760 334
rect 20824 270 20845 334
rect 20739 254 20845 270
rect 20739 190 20760 254
rect 20824 190 20845 254
rect 20739 173 20845 190
rect 20913 334 21019 351
rect 20913 270 20934 334
rect 20998 270 21019 334
rect 20913 254 21019 270
rect 20913 190 20934 254
rect 20998 190 21019 254
rect 20913 173 21019 190
rect 35574 345 35680 362
rect 35574 281 35595 345
rect 35659 281 35680 345
rect 35574 265 35680 281
rect 35574 201 35595 265
rect 35659 201 35680 265
rect 35574 184 35680 201
rect 35757 345 35863 362
rect 35757 281 35778 345
rect 35842 281 35863 345
rect 35757 265 35863 281
rect 35757 201 35778 265
rect 35842 201 35863 265
rect 35757 184 35863 201
rect 35940 345 36046 362
rect 35940 281 35961 345
rect 36025 281 36046 345
rect 35940 265 36046 281
rect 35940 201 35961 265
rect 36025 201 36046 265
rect 35940 184 36046 201
rect 51074 337 51180 354
rect 51074 273 51095 337
rect 51159 273 51180 337
rect 51074 257 51180 273
rect 51074 193 51095 257
rect 51159 193 51180 257
rect 51074 176 51180 193
rect 51257 337 51363 354
rect 51257 273 51278 337
rect 51342 273 51363 337
rect 51257 257 51363 273
rect 51257 193 51278 257
rect 51342 193 51363 257
rect 51257 176 51363 193
rect 51440 337 51546 354
rect 51440 273 51461 337
rect 51525 273 51546 337
rect 51440 257 51546 273
rect 51440 193 51461 257
rect 51525 193 51546 257
rect 51440 176 51546 193
<< via3 >>
rect 20604 19700 20668 19764
rect 20604 19620 20668 19684
rect 20778 19700 20842 19764
rect 20778 19620 20842 19684
rect 20952 19700 21016 19764
rect 20952 19620 21016 19684
rect 35579 19677 35643 19741
rect 35579 19597 35643 19661
rect 35762 19677 35826 19741
rect 35762 19597 35826 19661
rect 35945 19677 36009 19741
rect 35945 19597 36009 19661
rect 51077 19690 51141 19754
rect 51077 19610 51141 19674
rect 51260 19690 51324 19754
rect 51260 19610 51324 19674
rect 51443 19690 51507 19754
rect 51443 19610 51507 19674
rect 19081 17556 19145 17620
rect 19081 17476 19145 17540
rect 19255 17556 19319 17620
rect 19255 17476 19319 17540
rect 19429 17556 19493 17620
rect 19429 17476 19493 17540
rect 34058 17561 34122 17625
rect 34058 17481 34122 17545
rect 34241 17561 34305 17625
rect 34241 17481 34305 17545
rect 34424 17561 34488 17625
rect 34424 17481 34488 17545
rect 49552 17552 49616 17616
rect 49552 17472 49616 17536
rect 49735 17552 49799 17616
rect 49735 17472 49799 17536
rect 49918 17552 49982 17616
rect 49918 17472 49982 17536
rect 31111 15503 31161 15514
rect 31161 15503 31175 15514
rect 31111 15457 31175 15503
rect 31111 15450 31161 15457
rect 31161 15450 31175 15457
rect 19094 14628 19158 14692
rect 19094 14548 19158 14612
rect 19268 14628 19332 14692
rect 19268 14548 19332 14612
rect 19442 14628 19506 14692
rect 19442 14548 19506 14612
rect 32188 14625 32252 14689
rect 32188 14545 32252 14609
rect 32387 14625 32451 14689
rect 32387 14545 32451 14609
rect 34044 14626 34108 14690
rect 34044 14546 34108 14610
rect 34227 14626 34291 14690
rect 34227 14546 34291 14610
rect 34410 14626 34474 14690
rect 34410 14546 34474 14610
rect 49583 14623 49647 14687
rect 49583 14543 49647 14607
rect 49766 14623 49830 14687
rect 49766 14543 49830 14607
rect 49949 14623 50013 14687
rect 49949 14543 50013 14607
rect 20604 12492 20668 12556
rect 20604 12412 20668 12476
rect 20778 12492 20842 12556
rect 20778 12412 20842 12476
rect 20952 12492 21016 12556
rect 20952 12412 21016 12476
rect 35594 12503 35658 12567
rect 35594 12423 35658 12487
rect 35777 12503 35841 12567
rect 35777 12423 35841 12487
rect 35960 12503 36024 12567
rect 35960 12423 36024 12487
rect 51052 12494 51116 12558
rect 51052 12414 51116 12478
rect 51235 12494 51299 12558
rect 51235 12414 51299 12478
rect 51418 12494 51482 12558
rect 51418 12414 51482 12478
rect 31102 10321 31149 10330
rect 31149 10321 31166 10330
rect 31284 10321 31309 10330
rect 31309 10321 31348 10330
rect 31102 10278 31166 10321
rect 31284 10278 31348 10321
rect 31102 10266 31149 10278
rect 31149 10266 31166 10278
rect 31284 10266 31309 10278
rect 31309 10266 31348 10278
rect 32249 9947 32313 9961
rect 32329 9947 32393 9961
rect 32249 9897 32281 9947
rect 32281 9897 32313 9947
rect 32329 9897 32337 9947
rect 32337 9897 32393 9947
rect 31094 8992 31114 9007
rect 31114 8992 31146 9007
rect 31146 8992 31158 9007
rect 31284 8992 31290 9007
rect 31290 8992 31322 9007
rect 31322 8992 31348 9007
rect 31094 8953 31158 8992
rect 31284 8953 31348 8992
rect 31094 8943 31114 8953
rect 31114 8943 31146 8953
rect 31146 8943 31158 8953
rect 31284 8943 31290 8953
rect 31290 8943 31322 8953
rect 31322 8943 31348 8953
rect 3802 7451 3866 7515
rect 3802 7371 3866 7435
rect 4053 7451 4117 7515
rect 4053 7371 4117 7435
rect 4304 7451 4368 7515
rect 4304 7371 4368 7435
rect 20582 7454 20646 7518
rect 20582 7374 20646 7438
rect 20756 7454 20820 7518
rect 20756 7374 20820 7438
rect 20930 7454 20994 7518
rect 20930 7374 20994 7438
rect 35549 7461 35613 7525
rect 35549 7381 35613 7445
rect 35732 7461 35796 7525
rect 35732 7381 35796 7445
rect 35915 7461 35979 7525
rect 35915 7381 35979 7445
rect 51054 7453 51118 7517
rect 51054 7373 51118 7437
rect 51237 7453 51301 7517
rect 51237 7373 51301 7437
rect 51420 7453 51484 7517
rect 51420 7373 51484 7437
rect 2577 5322 2641 5386
rect 2753 5322 2817 5386
rect 2929 5322 2993 5386
rect 2577 5242 2641 5306
rect 2753 5242 2817 5306
rect 2929 5242 2993 5306
rect 19080 5328 19144 5392
rect 19080 5248 19144 5312
rect 19254 5328 19318 5392
rect 19254 5248 19318 5312
rect 19428 5328 19492 5392
rect 19428 5248 19492 5312
rect 34056 5329 34120 5393
rect 34056 5249 34120 5313
rect 34239 5329 34303 5393
rect 34239 5249 34303 5313
rect 34422 5329 34486 5393
rect 34422 5249 34486 5313
rect 49551 5325 49615 5389
rect 49551 5245 49615 5309
rect 49734 5325 49798 5389
rect 49734 5245 49798 5309
rect 49917 5325 49981 5389
rect 49917 5245 49981 5309
rect 31106 3268 31119 3278
rect 31119 3268 31155 3278
rect 31155 3268 31170 3278
rect 31280 3268 31303 3279
rect 31303 3268 31339 3279
rect 31339 3268 31344 3279
rect 31106 3233 31170 3268
rect 31280 3233 31344 3268
rect 31106 3214 31119 3233
rect 31119 3214 31155 3233
rect 31155 3214 31170 3233
rect 31280 3215 31303 3233
rect 31303 3215 31339 3233
rect 31339 3215 31344 3233
rect 2573 2389 2637 2453
rect 2573 2309 2637 2373
rect 2749 2389 2813 2453
rect 2749 2309 2813 2373
rect 2925 2389 2989 2453
rect 2925 2309 2989 2373
rect 19077 2392 19141 2456
rect 19077 2312 19141 2376
rect 19251 2392 19315 2456
rect 19251 2312 19315 2376
rect 19425 2392 19489 2456
rect 19425 2312 19489 2376
rect 34068 2388 34132 2452
rect 34068 2308 34132 2372
rect 34251 2388 34315 2452
rect 34251 2308 34315 2372
rect 34434 2388 34498 2452
rect 34434 2308 34498 2372
rect 49559 2392 49623 2456
rect 49559 2312 49623 2376
rect 49742 2392 49806 2456
rect 49742 2312 49806 2376
rect 49925 2392 49989 2456
rect 49925 2312 49989 2376
rect 3836 267 3900 331
rect 3836 187 3900 251
rect 4087 267 4151 331
rect 4087 187 4151 251
rect 4338 267 4402 331
rect 4338 187 4402 251
rect 20586 270 20650 334
rect 20586 190 20650 254
rect 20760 270 20824 334
rect 20760 190 20824 254
rect 20934 270 20998 334
rect 20934 190 20998 254
rect 35595 281 35659 345
rect 35595 201 35659 265
rect 35778 281 35842 345
rect 35778 201 35842 265
rect 35961 281 36025 345
rect 35961 201 36025 265
rect 51095 273 51159 337
rect 51095 193 51159 257
rect 51278 273 51342 337
rect 51278 193 51342 257
rect 51461 273 51525 337
rect 51461 193 51525 257
<< metal4 >>
rect 2472 5386 3090 20087
rect 2472 5322 2577 5386
rect 2641 5322 2753 5386
rect 2817 5322 2929 5386
rect 2993 5322 3090 5386
rect 2472 5306 3090 5322
rect 2472 5242 2577 5306
rect 2641 5242 2753 5306
rect 2817 5242 2929 5306
rect 2993 5242 3090 5306
rect 2472 2453 3090 5242
rect 2472 2389 2573 2453
rect 2637 2389 2749 2453
rect 2813 2389 2925 2453
rect 2989 2389 3090 2453
rect 2472 2373 3090 2389
rect 2472 2309 2573 2373
rect 2637 2309 2749 2373
rect 2813 2309 2925 2373
rect 2989 2309 3090 2373
rect 2472 38 3090 2309
rect 3705 7515 4489 20087
rect 3705 7451 3802 7515
rect 3866 7451 4053 7515
rect 4117 7451 4304 7515
rect 4368 7451 4489 7515
rect 3705 7435 4489 7451
rect 3705 7371 3802 7435
rect 3866 7371 4053 7435
rect 4117 7371 4304 7435
rect 4368 7371 4489 7435
rect 3705 331 4489 7371
rect 3705 267 3836 331
rect 3900 267 4087 331
rect 4151 267 4338 331
rect 4402 267 4489 331
rect 3705 251 4489 267
rect 3705 187 3836 251
rect 3900 187 4087 251
rect 4151 187 4338 251
rect 4402 187 4489 251
rect 3705 74 4489 187
rect 18972 17620 19590 20087
rect 18972 17556 19081 17620
rect 19145 17556 19255 17620
rect 19319 17556 19429 17620
rect 19493 17556 19590 17620
rect 18972 17540 19590 17556
rect 18972 17476 19081 17540
rect 19145 17476 19255 17540
rect 19319 17476 19429 17540
rect 19493 17476 19590 17540
rect 18972 14692 19590 17476
rect 18972 14628 19094 14692
rect 19158 14628 19268 14692
rect 19332 14628 19442 14692
rect 19506 14628 19590 14692
rect 18972 14612 19590 14628
rect 18972 14548 19094 14612
rect 19158 14548 19268 14612
rect 19332 14548 19442 14612
rect 19506 14548 19590 14612
rect 18972 5392 19590 14548
rect 18972 5328 19080 5392
rect 19144 5328 19254 5392
rect 19318 5328 19428 5392
rect 19492 5328 19590 5392
rect 18972 5312 19590 5328
rect 18972 5248 19080 5312
rect 19144 5248 19254 5312
rect 19318 5248 19428 5312
rect 19492 5248 19590 5312
rect 18972 2456 19590 5248
rect 18972 2392 19077 2456
rect 19141 2392 19251 2456
rect 19315 2392 19425 2456
rect 19489 2392 19590 2456
rect 18972 2376 19590 2392
rect 18972 2312 19077 2376
rect 19141 2312 19251 2376
rect 19315 2312 19425 2376
rect 19489 2312 19590 2376
rect 18972 38 19590 2312
rect 20472 19764 21090 20087
rect 20472 19700 20604 19764
rect 20668 19700 20778 19764
rect 20842 19700 20952 19764
rect 21016 19700 21090 19764
rect 20472 19684 21090 19700
rect 20472 19620 20604 19684
rect 20668 19620 20778 19684
rect 20842 19620 20952 19684
rect 21016 19620 21090 19684
rect 20472 12556 21090 19620
rect 33972 17625 34590 20087
rect 33972 17561 34058 17625
rect 34122 17561 34241 17625
rect 34305 17561 34424 17625
rect 34488 17561 34590 17625
rect 33972 17545 34590 17561
rect 33972 17481 34058 17545
rect 34122 17481 34241 17545
rect 34305 17481 34424 17545
rect 34488 17481 34590 17545
rect 20472 12492 20604 12556
rect 20668 12492 20778 12556
rect 20842 12492 20952 12556
rect 21016 12492 21090 12556
rect 20472 12476 21090 12492
rect 20472 12412 20604 12476
rect 20668 12412 20778 12476
rect 20842 12412 20952 12476
rect 21016 12412 21090 12476
rect 20472 7518 21090 12412
rect 31021 15514 31418 15648
rect 31021 15450 31111 15514
rect 31175 15450 31418 15514
rect 31021 10856 31418 15450
rect 31020 10495 31418 10856
rect 31021 10330 31418 10495
rect 31021 10266 31102 10330
rect 31166 10266 31284 10330
rect 31348 10266 31418 10330
rect 31021 10195 31418 10266
rect 32106 14689 32510 14819
rect 32106 14625 32188 14689
rect 32252 14625 32387 14689
rect 32451 14625 32510 14689
rect 32106 14609 32510 14625
rect 32106 14545 32188 14609
rect 32252 14545 32387 14609
rect 32451 14545 32510 14609
rect 32106 9989 32510 14545
rect 33972 14690 34590 17481
rect 33972 14626 34044 14690
rect 34108 14626 34227 14690
rect 34291 14626 34410 14690
rect 34474 14626 34590 14690
rect 33972 14610 34590 14626
rect 33972 14546 34044 14610
rect 34108 14546 34227 14610
rect 34291 14546 34410 14610
rect 34474 14546 34590 14610
rect 32106 9967 32514 9989
rect 32113 9961 32514 9967
rect 32113 9897 32249 9961
rect 32313 9897 32329 9961
rect 32393 9897 32514 9961
rect 32113 9878 32514 9897
rect 20472 7454 20582 7518
rect 20646 7454 20756 7518
rect 20820 7454 20930 7518
rect 20994 7454 21090 7518
rect 20472 7438 21090 7454
rect 20472 7374 20582 7438
rect 20646 7374 20756 7438
rect 20820 7374 20930 7438
rect 20994 7374 21090 7438
rect 20472 334 21090 7374
rect 31023 9007 31419 9105
rect 31023 8943 31094 9007
rect 31158 8943 31284 9007
rect 31348 8943 31419 9007
rect 31023 3279 31419 8943
rect 31023 3278 31280 3279
rect 31023 3214 31106 3278
rect 31170 3215 31280 3278
rect 31344 3215 31419 3279
rect 31170 3214 31419 3215
rect 31023 3089 31419 3214
rect 33972 5393 34590 14546
rect 33972 5329 34056 5393
rect 34120 5329 34239 5393
rect 34303 5329 34422 5393
rect 34486 5329 34590 5393
rect 33972 5313 34590 5329
rect 33972 5249 34056 5313
rect 34120 5249 34239 5313
rect 34303 5249 34422 5313
rect 34486 5249 34590 5313
rect 20472 270 20586 334
rect 20650 270 20760 334
rect 20824 270 20934 334
rect 20998 270 21090 334
rect 20472 254 21090 270
rect 20472 190 20586 254
rect 20650 190 20760 254
rect 20824 190 20934 254
rect 20998 190 21090 254
rect 20472 38 21090 190
rect 33972 2452 34590 5249
rect 33972 2388 34068 2452
rect 34132 2388 34251 2452
rect 34315 2388 34434 2452
rect 34498 2388 34590 2452
rect 33972 2372 34590 2388
rect 33972 2308 34068 2372
rect 34132 2308 34251 2372
rect 34315 2308 34434 2372
rect 34498 2308 34590 2372
rect 33972 38 34590 2308
rect 35472 19741 36090 20087
rect 35472 19677 35579 19741
rect 35643 19677 35762 19741
rect 35826 19677 35945 19741
rect 36009 19677 36090 19741
rect 35472 19661 36090 19677
rect 35472 19597 35579 19661
rect 35643 19597 35762 19661
rect 35826 19597 35945 19661
rect 36009 19597 36090 19661
rect 35472 12567 36090 19597
rect 35472 12503 35594 12567
rect 35658 12503 35777 12567
rect 35841 12503 35960 12567
rect 36024 12503 36090 12567
rect 35472 12487 36090 12503
rect 35472 12423 35594 12487
rect 35658 12423 35777 12487
rect 35841 12423 35960 12487
rect 36024 12423 36090 12487
rect 35472 7525 36090 12423
rect 35472 7461 35549 7525
rect 35613 7461 35732 7525
rect 35796 7461 35915 7525
rect 35979 7461 36090 7525
rect 35472 7445 36090 7461
rect 35472 7381 35549 7445
rect 35613 7381 35732 7445
rect 35796 7381 35915 7445
rect 35979 7381 36090 7445
rect 35472 345 36090 7381
rect 35472 281 35595 345
rect 35659 281 35778 345
rect 35842 281 35961 345
rect 36025 281 36090 345
rect 35472 265 36090 281
rect 35472 201 35595 265
rect 35659 201 35778 265
rect 35842 201 35961 265
rect 36025 201 36090 265
rect 35472 38 36090 201
rect 49472 17616 50090 20087
rect 49472 17552 49552 17616
rect 49616 17552 49735 17616
rect 49799 17552 49918 17616
rect 49982 17552 50090 17616
rect 49472 17536 50090 17552
rect 49472 17472 49552 17536
rect 49616 17472 49735 17536
rect 49799 17472 49918 17536
rect 49982 17472 50090 17536
rect 49472 14687 50090 17472
rect 49472 14623 49583 14687
rect 49647 14623 49766 14687
rect 49830 14623 49949 14687
rect 50013 14623 50090 14687
rect 49472 14607 50090 14623
rect 49472 14543 49583 14607
rect 49647 14543 49766 14607
rect 49830 14543 49949 14607
rect 50013 14543 50090 14607
rect 49472 5389 50090 14543
rect 49472 5325 49551 5389
rect 49615 5325 49734 5389
rect 49798 5325 49917 5389
rect 49981 5325 50090 5389
rect 49472 5309 50090 5325
rect 49472 5245 49551 5309
rect 49615 5245 49734 5309
rect 49798 5245 49917 5309
rect 49981 5245 50090 5309
rect 49472 2456 50090 5245
rect 49472 2392 49559 2456
rect 49623 2392 49742 2456
rect 49806 2392 49925 2456
rect 49989 2392 50090 2456
rect 49472 2376 50090 2392
rect 49472 2312 49559 2376
rect 49623 2312 49742 2376
rect 49806 2312 49925 2376
rect 49989 2312 50090 2376
rect 49472 38 50090 2312
rect 50972 19754 51590 20087
rect 50972 19690 51077 19754
rect 51141 19690 51260 19754
rect 51324 19690 51443 19754
rect 51507 19690 51590 19754
rect 50972 19674 51590 19690
rect 50972 19610 51077 19674
rect 51141 19610 51260 19674
rect 51324 19610 51443 19674
rect 51507 19610 51590 19674
rect 50972 12558 51590 19610
rect 50972 12494 51052 12558
rect 51116 12494 51235 12558
rect 51299 12494 51418 12558
rect 51482 12494 51590 12558
rect 50972 12478 51590 12494
rect 50972 12414 51052 12478
rect 51116 12414 51235 12478
rect 51299 12414 51418 12478
rect 51482 12414 51590 12478
rect 50972 7517 51590 12414
rect 50972 7453 51054 7517
rect 51118 7453 51237 7517
rect 51301 7453 51420 7517
rect 51484 7453 51590 7517
rect 50972 7437 51590 7453
rect 50972 7373 51054 7437
rect 51118 7373 51237 7437
rect 51301 7373 51420 7437
rect 51484 7373 51590 7437
rect 50972 337 51590 7373
rect 50972 273 51095 337
rect 51159 273 51278 337
rect 51342 273 51461 337
rect 51525 273 51590 337
rect 50972 257 51590 273
rect 50972 193 51095 257
rect 51159 193 51278 257
rect 51342 193 51461 257
rect 51525 193 51590 257
rect 50972 38 51590 193
use NBR128half  NBR128half_0
timestamp 1656729169
transform 1 0 1238 0 1 12369
box -430 -58 60412 7443
use NBR128half_bottom  NBR128half_bottom_0
timestamp 1656729169
transform -1 0 61449 0 1 138
box -430 -58 60604 7443
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0
timestamp 1656729169
transform 1 0 28089 0 1 9381
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0
timestamp 1656729169
transform 1 0 28625 0 1 9381
box -38 -48 866 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0
timestamp 1656729169
transform 1 0 31445 0 1 9381
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1656729169
transform 1 0 29529 0 1 9381
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1656729169
transform 1 0 28457 0 1 9381
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1656729169
transform 1 0 31188 0 1 9381
box -38 -48 130 592
use unitcell_nbr  unitcell_nbr_0
timestamp 1656729169
transform 1 0 62216 0 1 13553
box -574 -1185 1322 1192
<< labels >>
flabel metal3 s 509 9570 755 9660 1 FreeSans 500 0 0 0 RESET
port 1 nsew
flabel metal4 s 2472 38 3090 20087 1 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal4 s 18972 38 19590 20087 1 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal4 s 33972 38 34590 20087 1 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal4 s 49472 38 50090 20087 1 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal4 s 3705 74 4489 20087 1 FreeSans 2000 0 0 0 VSS
port 3 nsew
flabel metal4 s 20472 38 21090 20087 1 FreeSans 2000 0 0 0 VSS
port 3 nsew
flabel metal4 s 35472 38 36090 20087 1 FreeSans 2000 0 0 0 VSS
port 3 nsew
flabel metal4 s 50972 38 51590 20087 1 FreeSans 2000 0 0 0 VSS
port 3 nsew
flabel metal2 s 61156 19017 61200 19992 1 FreeSans 2000 0 0 0 C[0]
port 4 nsew
flabel metal2 s 59268 19017 59312 19992 1 FreeSans 2000 0 0 0 C[1]
port 5 nsew
flabel metal2 s 57380 19017 57424 19992 1 FreeSans 2000 0 0 0 C[2]
port 6 nsew
flabel metal2 s 55492 19017 55536 19992 1 FreeSans 2000 0 0 0 C[3]
port 7 nsew
flabel metal2 s 53604 19017 53648 19992 1 FreeSans 2000 0 0 0 C[4]
port 8 nsew
flabel metal2 s 51716 19017 51760 19992 1 FreeSans 2000 0 0 0 C[5]
port 9 nsew
flabel metal2 s 47940 19017 47984 19992 1 FreeSans 2000 0 0 0 C[7]
port 10 nsew
flabel metal2 s 46052 19017 46096 19992 1 FreeSans 2000 0 0 0 C[8]
port 11 nsew
flabel metal2 s 44164 19017 44208 19992 1 FreeSans 2000 0 0 0 C[9]
port 12 nsew
flabel metal2 s 42276 19017 42320 19992 1 FreeSans 2000 0 0 0 C[10]
port 13 nsew
flabel metal2 s 40388 19017 40432 19992 1 FreeSans 2000 0 0 0 C[11]
port 14 nsew
flabel metal2 s 38500 19017 38544 19992 1 FreeSans 2000 0 0 0 C[12]
port 15 nsew
flabel metal2 s 36612 19017 36656 19992 1 FreeSans 2000 0 0 0 C[13]
port 16 nsew
flabel metal2 s 34724 19017 34768 19992 1 FreeSans 2000 0 0 0 C[14]
port 17 nsew
flabel metal2 s 32836 19017 32880 19992 1 FreeSans 2000 0 0 0 C[15]
port 18 nsew
flabel metal2 s 30948 19017 30992 19992 1 FreeSans 2000 0 0 0 C[16]
port 19 nsew
flabel metal2 s 29060 19017 29104 19992 1 FreeSans 2000 0 0 0 C[17]
port 20 nsew
flabel metal2 s 27172 19017 27216 19992 1 FreeSans 2000 0 0 0 C[18]
port 21 nsew
flabel metal2 s 25284 19017 25328 19992 1 FreeSans 2000 0 0 0 C[19]
port 22 nsew
flabel metal2 s 23396 19017 23440 19992 1 FreeSans 2000 0 0 0 C[20]
port 23 nsew
flabel metal2 s 21508 19017 21552 19992 1 FreeSans 2000 0 0 0 C[21]
port 24 nsew
flabel metal2 s 19620 19017 19664 19992 1 FreeSans 2000 0 0 0 C[22]
port 25 nsew
flabel metal2 s 17732 19017 17776 19992 1 FreeSans 2000 0 0 0 C[23]
port 26 nsew
flabel metal2 s 15844 19017 15888 19992 1 FreeSans 2000 0 0 0 C[24]
port 27 nsew
flabel metal2 s 13956 19017 14000 19992 1 FreeSans 2000 0 0 0 C[25]
port 28 nsew
flabel metal2 s 12068 19017 12112 19992 1 FreeSans 2000 0 0 0 C[26]
port 29 nsew
flabel metal2 s 10180 19017 10224 19992 1 FreeSans 2000 0 0 0 C[27]
port 30 nsew
flabel metal2 s 8292 19017 8336 19992 1 FreeSans 2000 0 0 0 C[28]
port 31 nsew
flabel metal2 s 6404 19017 6448 19992 1 FreeSans 2000 0 0 0 C[29]
port 32 nsew
flabel metal2 s 4516 19017 4560 19992 1 FreeSans 2000 0 0 0 C[30]
port 33 nsew
flabel metal2 s 49828 19017 49872 20151 1 FreeSans 1000 0 0 0 C[6]
port 34 nsew
flabel metal2 s 2628 19017 2672 20184 1 FreeSans 2000 0 0 0 C[31]
port 35 nsew
flabel metal1 s 0 9748 490 9810 1 FreeSans 1000 0 0 0 C[32]
port 36 nsew
flabel metal1 s 0 9606 490 9668 1 FreeSans 1000 0 0 0 C[33]
port 37 nsew
flabel metal1 s 0 9464 490 9526 1 FreeSans 1000 0 0 0 C[34]
port 38 nsew
flabel metal1 s 0 9322 490 9384 1 FreeSans 1000 0 0 0 C[35]
port 39 nsew
flabel metal1 s 0 9180 490 9242 1 FreeSans 1000 0 0 0 C[36]
port 40 nsew
flabel metal1 s 0 9038 490 9100 1 FreeSans 1000 0 0 0 C[37]
port 41 nsew
flabel metal1 s 0 8896 490 8958 1 FreeSans 1000 0 0 0 C[38]
port 42 nsew
flabel metal1 s 0 8754 490 8816 1 FreeSans 1000 0 0 0 C[39]
port 43 nsew
flabel metal1 s 0 8612 490 8674 1 FreeSans 1000 0 0 0 C[40]
port 44 nsew
flabel metal1 s 0 8470 490 8532 1 FreeSans 1000 0 0 0 C[41]
port 45 nsew
flabel metal1 s 0 8328 490 8390 1 FreeSans 1000 0 0 0 C[42]
port 46 nsew
flabel metal1 s 0 8186 490 8248 1 FreeSans 1000 0 0 0 C[43]
port 47 nsew
flabel metal1 s 0 8044 490 8106 1 FreeSans 1000 0 0 0 C[44]
port 48 nsew
flabel metal1 s 0 7902 490 7964 1 FreeSans 1000 0 0 0 C[45]
port 49 nsew
flabel metal1 s 0 7760 490 7822 1 FreeSans 1000 0 0 0 C[46]
port 50 nsew
flabel metal1 s 62092 7758 64102 7820 1 FreeSans 1000 0 0 0 C[47]
port 51 nsew
flabel metal1 s 62092 7900 64102 7962 1 FreeSans 1000 0 0 0 C[48]
port 52 nsew
flabel metal1 s 62092 8042 64102 8104 1 FreeSans 1000 0 0 0 C[49]
port 53 nsew
flabel metal1 s 62092 8184 64102 8246 1 FreeSans 1000 0 0 0 C[50]
port 54 nsew
flabel metal1 s 62092 8326 64102 8388 1 FreeSans 1000 0 0 0 C[51]
port 55 nsew
flabel metal1 s 62092 8468 64102 8530 1 FreeSans 1000 0 0 0 C[52]
port 56 nsew
flabel metal1 s 62092 8610 64102 8672 1 FreeSans 1000 0 0 0 C[53]
port 57 nsew
flabel metal1 s 62092 8752 64102 8814 1 FreeSans 1000 0 0 0 C[54]
port 58 nsew
flabel metal1 s 62092 8894 64102 8956 1 FreeSans 1000 0 0 0 C[55]
port 59 nsew
flabel metal1 s 62092 9036 64102 9098 1 FreeSans 1000 0 0 0 C[56]
port 60 nsew
flabel metal1 s 62092 9178 64102 9240 1 FreeSans 1000 0 0 0 C[57]
port 61 nsew
flabel metal1 s 62092 9320 64102 9382 1 FreeSans 1000 0 0 0 C[58]
port 62 nsew
flabel metal1 s 62092 9462 64102 9524 1 FreeSans 1000 0 0 0 C[59]
port 63 nsew
flabel metal1 s 62092 9604 64102 9666 1 FreeSans 1000 0 0 0 C[60]
port 64 nsew
flabel metal1 s 62092 9746 64102 9808 1 FreeSans 1000 0 0 0 C[61]
port 65 nsew
flabel metal1 s 62092 9888 64102 9950 1 FreeSans 1000 0 0 0 C[62]
port 66 nsew
flabel metal1 s 0 10032 490 10094 1 FreeSans 1000 0 0 0 C[95]
port 67 nsew
flabel metal1 s 0 10174 490 10236 1 FreeSans 1000 0 0 0 C[96]
port 68 nsew
flabel metal1 s 0 10316 490 10378 1 FreeSans 1000 0 0 0 C[97]
port 69 nsew
flabel metal1 s 0 10458 490 10520 1 FreeSans 1000 0 0 0 C[98]
port 70 nsew
flabel metal1 s 0 10600 490 10662 1 FreeSans 1000 0 0 0 C[99]
port 71 nsew
flabel metal1 s 0 10742 490 10804 1 FreeSans 1000 0 0 0 C[100]
port 72 nsew
flabel metal1 s 0 10884 490 10946 1 FreeSans 1000 0 0 0 C[101]
port 73 nsew
flabel metal1 s 0 11026 490 11088 1 FreeSans 1000 0 0 0 C[102]
port 74 nsew
flabel metal1 s 0 11168 490 11230 1 FreeSans 1000 0 0 0 C[103]
port 75 nsew
flabel metal1 s 0 11310 490 11372 1 FreeSans 1000 0 0 0 C[104]
port 76 nsew
flabel metal1 s 0 11452 490 11514 1 FreeSans 1000 0 0 0 C[105]
port 77 nsew
flabel metal1 s 0 11594 490 11656 1 FreeSans 1000 0 0 0 C[106]
port 78 nsew
flabel metal1 s 0 11736 490 11798 1 FreeSans 1000 0 0 0 C[107]
port 79 nsew
flabel metal1 s 0 11878 490 11940 1 FreeSans 1000 0 0 0 C[108]
port 80 nsew
flabel metal1 s 0 12020 490 12082 1 FreeSans 1000 0 0 0 C[109]
port 81 nsew
flabel metal1 s 0 12162 490 12224 1 FreeSans 1000 0 0 0 C[110]
port 82 nsew
flabel metal1 s 62092 12160 64102 12222 1 FreeSans 1000 0 0 0 C[111]
port 83 nsew
flabel metal1 s 62092 12018 64102 12080 1 FreeSans 1000 0 0 0 C[112]
port 84 nsew
flabel metal1 s 62092 11876 64102 11938 1 FreeSans 1000 0 0 0 C[113]
port 85 nsew
flabel metal1 s 62092 11734 64102 11796 1 FreeSans 1000 0 0 0 C[114]
port 86 nsew
flabel metal1 s 62092 11592 64102 11654 1 FreeSans 1000 0 0 0 C[115]
port 87 nsew
flabel metal1 s 62092 11450 64102 11512 1 FreeSans 1000 0 0 0 C[116]
port 88 nsew
flabel metal1 s 62092 11308 64102 11370 1 FreeSans 1000 0 0 0 C[117]
port 89 nsew
flabel metal1 s 62092 11166 64102 11228 1 FreeSans 1000 0 0 0 C[118]
port 90 nsew
flabel metal1 s 62092 11024 64102 11086 1 FreeSans 1000 0 0 0 C[119]
port 91 nsew
flabel metal1 s 62092 10882 64102 10944 1 FreeSans 1000 0 0 0 C[120]
port 92 nsew
flabel metal1 s 62092 10740 64102 10802 1 FreeSans 1000 0 0 0 C[121]
port 93 nsew
flabel metal1 s 62092 10598 64102 10660 1 FreeSans 1000 0 0 0 C[122]
port 94 nsew
flabel metal1 s 62092 10456 64102 10518 1 FreeSans 1000 0 0 0 C[123]
port 95 nsew
flabel metal1 s 62092 10314 64102 10376 1 FreeSans 1000 0 0 0 C[124]
port 96 nsew
flabel metal1 s 62092 10172 64102 10234 1 FreeSans 1000 0 0 0 C[125]
port 97 nsew
flabel metal1 s 62092 10030 64102 10092 1 FreeSans 1000 0 0 0 C[126]
port 98 nsew
flabel metal3 s 61722 11938 64105 12036 1 FreeSans 1000 0 0 0 C[127]
port 99 nsew
flabel metal2 s 61385 0 61441 930 1 FreeSans 2000 0 0 0 C[63]
port 100 nsew
flabel metal2 s 59497 0 59553 930 1 FreeSans 2000 0 0 0 C[64]
port 101 nsew
flabel metal2 s 57609 0 57665 930 1 FreeSans 2000 0 0 0 C[65]
port 102 nsew
flabel metal2 s 55721 0 55777 930 1 FreeSans 2000 0 0 0 C[66]
port 103 nsew
flabel metal2 s 53833 0 53889 930 1 FreeSans 2000 0 0 0 C[67]
port 104 nsew
flabel metal2 s 51945 0 52001 930 1 FreeSans 2000 0 0 0 C[68]
port 105 nsew
flabel metal2 s 50057 0 50113 930 1 FreeSans 2000 0 0 0 C[69]
port 106 nsew
flabel metal2 s 48169 0 48225 930 1 FreeSans 2000 0 0 0 C[70]
port 107 nsew
flabel metal2 s 46281 0 46337 930 1 FreeSans 2000 0 0 0 C[71]
port 108 nsew
flabel metal2 s 44393 0 44449 930 1 FreeSans 2000 0 0 0 C[72]
port 109 nsew
flabel metal2 s 42505 0 42561 930 1 FreeSans 2000 0 0 0 C[73]
port 110 nsew
flabel metal2 s 40617 0 40673 930 1 FreeSans 2000 0 0 0 C[74]
port 111 nsew
flabel metal2 s 38729 0 38785 930 1 FreeSans 2000 0 0 0 C[75]
port 112 nsew
flabel metal2 s 36841 0 36897 930 1 FreeSans 2000 0 0 0 C[76]
port 113 nsew
flabel metal2 s 34953 0 35009 930 1 FreeSans 2000 0 0 0 C[77]
port 114 nsew
flabel metal2 s 33065 0 33121 930 1 FreeSans 2000 0 0 0 C[78]
port 115 nsew
flabel metal2 s 31177 0 31233 930 1 FreeSans 2000 0 0 0 C[79]
port 116 nsew
flabel metal2 s 29289 0 29345 930 1 FreeSans 2000 0 0 0 C[80]
port 117 nsew
flabel metal2 s 27401 0 27457 930 1 FreeSans 2000 0 0 0 C[81]
port 118 nsew
flabel metal2 s 25513 0 25569 930 1 FreeSans 2000 0 0 0 C[82]
port 119 nsew
flabel metal2 s 23625 0 23681 930 1 FreeSans 2000 0 0 0 C[83]
port 120 nsew
flabel metal2 s 21737 0 21793 930 1 FreeSans 2000 0 0 0 C[84]
port 121 nsew
flabel metal2 s 19849 0 19905 930 1 FreeSans 2000 0 0 0 C[85]
port 122 nsew
flabel metal2 s 17961 0 18017 930 1 FreeSans 2000 0 0 0 C[86]
port 123 nsew
flabel metal2 s 16073 0 16129 930 1 FreeSans 2000 0 0 0 C[87]
port 124 nsew
flabel metal2 s 14185 0 14241 930 1 FreeSans 2000 0 0 0 C[88]
port 125 nsew
flabel metal2 s 12297 0 12353 930 1 FreeSans 2000 0 0 0 C[89]
port 126 nsew
flabel metal2 s 10409 0 10465 930 1 FreeSans 2000 0 0 0 C[90]
port 127 nsew
flabel metal2 s 8521 0 8577 930 1 FreeSans 2000 0 0 0 C[91]
port 128 nsew
flabel metal2 s 6633 0 6689 930 1 FreeSans 2000 0 0 0 C[92]
port 129 nsew
flabel metal2 s 4745 0 4801 930 1 FreeSans 2000 0 0 0 C[93]
port 130 nsew
flabel metal2 s 2857 0 2913 930 1 FreeSans 2000 0 0 0 C[94]
port 131 nsew
flabel metal1 s 63486 13150 64108 13226 1 FreeSans 4000 0 0 0 OUT
port 132 nsew
<< properties >>
string GDS_END 9253134
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/merge/design_merged.gds
string GDS_START 9171970
<< end >>
