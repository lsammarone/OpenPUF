magic
tech sky130A
timestamp 1483428465
<< checkpaint >>
rect -1130 -720 1130 720
<< metal3 >>
rect -500 76 500 90
rect -500 -76 -496 76
rect 496 -76 500 76
rect -500 -90 500 -76
<< via3 >>
rect -496 -76 496 76
<< metal4 >>
rect -500 76 500 90
rect -500 -76 -496 76
rect 496 -76 500 76
rect -500 -90 500 -76
<< end >>
