magic
tech sky130A
timestamp 1483428465
<< checkpaint >>
rect -739 -654 739 654
<< metal1 >>
rect -109 13 109 24
rect -83 -13 -77 13
rect -51 -13 -45 13
rect -19 -13 -13 13
rect 13 -13 19 13
rect 45 -13 51 13
rect 77 -13 83 13
rect -109 -24 109 -13
<< via1 >>
rect -109 -13 -83 13
rect -77 -13 -51 13
rect -45 -13 -19 13
rect -13 -13 13 13
rect 19 -13 45 13
rect 51 -13 77 13
rect 83 -13 109 13
<< metal2 >>
rect -109 13 109 24
rect -83 -13 -77 13
rect -51 -13 -45 13
rect -19 -13 -13 13
rect 13 -13 19 13
rect 45 -13 51 13
rect 77 -13 83 13
rect -109 -24 109 -13
<< end >>
