magic
tech sky130A
magscale 1 2
timestamp 1483428465
<< checkpaint >>
rect -2312 -1440 2311 1440
<< metal3 >>
rect -1052 152 1051 180
rect -1052 -152 -1032 152
rect 1032 -152 1051 152
rect -1052 -180 1051 -152
<< via3 >>
rect -1032 -152 1032 152
<< metal4 >>
rect -1052 152 1051 180
rect -1052 -152 -1032 152
rect 1032 -152 1051 152
rect -1052 -180 1051 -152
<< end >>
