magic
tech sky130A
magscale 1 2
timestamp 1655348380
<< nwell >>
rect -404 1022 772 1034
rect -396 704 772 1022
rect -404 700 772 704
rect 258 -422 630 -22
<< poly >>
rect 194 218 224 220
rect 194 188 328 218
rect 298 20 328 188
rect 24 -10 506 20
rect 24 -168 54 -10
rect 474 -92 506 -10
rect 24 -198 110 -168
rect 80 -272 110 -198
<< locali >>
rect -398 970 -336 1004
rect -114 998 68 1003
rect 180 1002 458 1004
rect 346 998 460 1002
rect -109 969 78 998
rect 342 969 487 998
rect 160 818 226 856
rect -322 666 -321 700
rect -287 666 -286 700
rect -150 662 -148 696
rect -114 662 -112 696
rect 256 690 258 692
rect 490 690 491 698
rect 224 658 258 690
rect 480 664 491 690
rect 525 690 526 698
rect 525 664 544 690
rect 664 664 665 698
rect 699 664 700 698
rect 480 658 544 664
rect -240 580 -204 582
rect -240 546 -239 580
rect -205 546 -204 580
rect -240 544 -204 546
rect 578 575 614 576
rect 578 541 579 575
rect 613 541 614 575
rect 578 540 614 541
rect -356 425 -330 458
rect -356 214 -322 425
rect -125 122 -91 457
rect 240 240 622 280
rect 80 172 94 206
rect -125 118 0 122
rect -125 88 10 118
rect 442 80 488 82
rect 442 78 446 80
rect 270 76 446 78
rect 10 44 46 62
rect 242 46 446 76
rect 480 46 488 80
rect 242 44 488 46
rect 442 38 488 44
rect -459 -65 -425 -44
rect 588 -118 622 240
rect -100 -162 106 -118
rect 306 -162 494 -118
rect 546 -158 622 -118
rect -78 -324 -64 -294
rect -74 -326 -64 -324
rect -460 -386 -456 -352
rect -422 -386 -418 -352
rect 634 -362 778 -340
rect 1234 -346 1272 -344
rect 1038 -358 1082 -356
rect 488 -368 554 -366
rect 634 -368 792 -362
rect 488 -372 792 -368
rect 530 -382 792 -372
rect 530 -402 674 -382
rect 726 -388 792 -382
rect 1038 -392 1043 -358
rect 1077 -392 1082 -358
rect 1234 -380 1236 -346
rect 1270 -380 1272 -346
rect 1234 -382 1272 -380
rect 1038 -394 1082 -392
rect 222 -484 502 -450
rect -332 -526 -48 -494
rect -378 -530 128 -526
rect -378 -554 -318 -530
rect -84 -562 128 -530
rect 454 -572 502 -484
rect -176 -600 -130 -590
rect -176 -634 -170 -600
rect -136 -620 -130 -600
rect 454 -606 462 -572
rect 496 -606 502 -572
rect 454 -618 502 -606
rect -136 -634 -126 -620
rect -176 -704 -126 -634
rect -258 -740 -126 -704
rect -258 -788 -222 -740
rect 78 -766 81 -729
rect -74 -788 82 -766
rect -258 -802 82 -788
rect -258 -824 -38 -802
rect 214 -978 266 -936
<< viali >>
rect -321 666 -287 700
rect -148 662 -114 696
rect 491 664 525 698
rect 665 664 699 698
rect -239 546 -205 580
rect 579 541 613 575
rect -356 180 -322 214
rect 446 46 480 80
rect -456 -386 -422 -352
rect 1043 -392 1077 -358
rect 1236 -380 1270 -346
rect 822 -490 856 -456
rect -170 -634 -136 -600
rect 462 -606 496 -572
<< metal1 >>
rect -574 1120 1322 1192
rect -574 1004 961 1120
rect 1269 1004 1322 1120
rect -574 938 1322 1004
rect -514 -66 -436 938
rect 102 922 146 938
rect -336 746 30 778
rect -336 708 -308 746
rect 226 742 546 774
rect -336 700 -270 708
rect -336 666 -321 700
rect -287 666 -270 700
rect -336 654 -270 666
rect -164 704 -96 710
rect 518 706 546 742
rect -164 652 -154 704
rect -102 652 -96 704
rect -164 646 -96 652
rect 476 698 546 706
rect 476 664 491 698
rect 525 664 546 698
rect 476 646 546 664
rect 652 706 716 712
rect 652 654 658 706
rect 710 654 716 706
rect 652 648 716 654
rect -254 592 -186 598
rect -254 540 -246 592
rect -194 540 -186 592
rect -254 530 -186 540
rect 564 590 628 596
rect 564 538 570 590
rect 622 538 628 590
rect 564 532 628 538
rect -374 357 -310 364
rect -374 324 -368 357
rect -316 324 -310 357
rect -198 357 -134 364
rect -198 324 -192 357
rect -316 305 -192 324
rect -140 305 -134 357
rect -368 296 -134 305
rect -218 244 -14 258
rect -218 230 36 244
rect -374 224 -308 230
rect -374 172 -366 224
rect -314 172 -308 224
rect -374 166 -308 172
rect -218 -120 -190 230
rect 106 172 402 206
rect 4 108 64 112
rect 4 56 8 108
rect 60 56 64 108
rect 4 52 64 56
rect 368 -10 402 172
rect 430 90 458 422
rect 430 80 498 90
rect 430 46 446 80
rect 480 46 498 80
rect 430 32 498 46
rect -158 -38 402 -10
rect -158 -84 -92 -38
rect -218 -122 -146 -120
rect -218 -124 -190 -122
rect -218 -148 -192 -124
rect -102 -148 -36 -142
rect -102 -200 -96 -148
rect -44 -200 -36 -148
rect -102 -208 -36 -200
rect 368 -212 402 -38
rect 488 -86 554 -30
rect 662 -40 1286 -8
rect 662 -92 692 -40
rect 744 -92 1286 -40
rect 662 -110 1286 -92
rect 446 -128 512 -122
rect 446 -180 454 -128
rect 506 -180 512 -128
rect 446 -186 512 -180
rect -554 -340 -486 -334
rect -554 -392 -547 -340
rect -495 -346 -486 -340
rect 1028 -344 1100 -340
rect -495 -352 -402 -346
rect -495 -386 -456 -352
rect -422 -386 -402 -352
rect -495 -392 -402 -386
rect -554 -396 -402 -392
rect -554 -398 -486 -396
rect -158 -416 -92 -358
rect 488 -412 554 -356
rect 1028 -396 1037 -344
rect 1089 -396 1100 -344
rect 1028 -408 1100 -396
rect 1224 -346 1298 -326
rect 1224 -380 1236 -346
rect 1270 -380 1298 -346
rect 1224 -404 1298 -380
rect 810 -456 868 -442
rect 810 -476 822 -456
rect 386 -490 822 -476
rect 856 -490 868 -456
rect 386 -510 868 -490
rect -414 -582 -356 -576
rect -414 -628 -411 -582
rect -466 -634 -411 -628
rect -359 -634 -356 -582
rect -182 -586 -124 -578
rect -190 -592 -116 -586
rect -466 -640 -356 -634
rect -466 -930 -382 -640
rect -296 -654 -284 -620
rect -190 -644 -179 -592
rect -127 -644 -116 -592
rect -36 -602 28 -536
rect 446 -560 522 -554
rect 446 -612 454 -560
rect 506 -612 522 -560
rect 446 -618 522 -612
rect -190 -650 -116 -644
rect -182 -656 -124 -650
rect 662 -654 1284 -556
rect 662 -930 760 -654
rect -566 -1004 1322 -930
rect -566 -1120 961 -1004
rect 1269 -1120 1322 -1004
rect -566 -1184 1322 -1120
<< via1 >>
rect 961 1004 1269 1120
rect -154 696 -102 704
rect -154 662 -148 696
rect -148 662 -114 696
rect -114 662 -102 696
rect -154 652 -102 662
rect 658 698 710 706
rect 658 664 665 698
rect 665 664 699 698
rect 699 664 710 698
rect 658 654 710 664
rect -246 580 -194 592
rect -246 546 -239 580
rect -239 546 -205 580
rect -205 546 -194 580
rect -246 540 -194 546
rect 570 575 622 590
rect 570 541 579 575
rect 579 541 613 575
rect 613 541 622 575
rect 570 538 622 541
rect -368 305 -316 357
rect -192 305 -140 357
rect -366 214 -314 224
rect -366 180 -356 214
rect -356 180 -322 214
rect -322 180 -314 214
rect -366 172 -314 180
rect -342 -86 -290 -34
rect 8 56 60 108
rect -96 -200 -44 -148
rect 692 -92 744 -40
rect 454 -180 506 -128
rect -547 -392 -495 -340
rect 1037 -358 1089 -344
rect 1037 -392 1043 -358
rect 1043 -392 1077 -358
rect 1077 -392 1089 -358
rect 1037 -396 1089 -392
rect -411 -634 -359 -582
rect -179 -600 -127 -592
rect -179 -634 -170 -600
rect -170 -634 -136 -600
rect -136 -634 -127 -600
rect -179 -644 -127 -634
rect 454 -572 506 -560
rect 454 -606 462 -572
rect 462 -606 496 -572
rect 496 -606 506 -572
rect 454 -612 506 -606
rect 961 -1120 1269 -1004
<< metal2 >>
rect 940 1120 1290 1134
rect 940 1004 961 1120
rect 1269 1004 1290 1120
rect 940 990 1290 1004
rect -566 816 1050 844
rect -124 710 -96 816
rect -164 704 -96 710
rect -164 652 -154 704
rect -102 652 -96 704
rect 650 712 678 816
rect 650 706 716 712
rect 650 692 658 706
rect -164 646 -96 652
rect 652 654 658 692
rect 710 654 716 706
rect 652 648 716 654
rect -254 592 -186 598
rect -254 540 -246 592
rect -194 540 -186 592
rect 564 590 628 596
rect 564 560 570 590
rect -254 530 -186 540
rect 354 538 570 560
rect 622 538 628 590
rect 354 532 628 538
rect -374 357 -310 364
rect -374 326 -368 357
rect -566 305 -368 326
rect -316 305 -310 357
rect -566 298 -310 305
rect -566 296 -368 298
rect -566 290 -374 296
rect -374 224 -308 230
rect -374 172 -366 224
rect -314 172 -308 224
rect -374 166 -308 172
rect -374 44 -346 166
rect -414 16 -346 44
rect -554 -340 -486 -334
rect -554 -392 -547 -340
rect -495 -392 -486 -340
rect -554 -398 -486 -392
rect -554 -1184 -510 -398
rect -414 -568 -386 16
rect -352 -34 -290 -28
rect -352 -86 -342 -34
rect -254 -42 -226 530
rect 136 462 168 504
rect -198 357 -134 364
rect -198 305 -192 357
rect -140 324 -134 357
rect -140 305 180 324
rect -198 296 180 305
rect -2 108 70 120
rect -2 56 8 108
rect 60 56 70 108
rect -2 44 70 56
rect 34 42 70 44
rect -254 -70 34 -42
rect -352 -92 -290 -86
rect -318 -138 -290 -92
rect -318 -142 -74 -138
rect -318 -148 -36 -142
rect -318 -166 -96 -148
rect -102 -200 -96 -166
rect -44 -200 -36 -148
rect -102 -208 -36 -200
rect -414 -582 -350 -568
rect 6 -576 34 -70
rect 138 -572 166 -536
rect -414 -634 -411 -582
rect -359 -634 -350 -582
rect -414 -650 -350 -634
rect -180 -592 34 -576
rect -180 -644 -179 -592
rect -127 -604 34 -592
rect 354 -586 382 532
rect 786 290 1322 326
rect 686 -40 750 -32
rect 686 -92 692 -40
rect 744 -92 750 -40
rect 686 -100 750 -92
rect 446 -128 512 -122
rect 446 -180 454 -128
rect 506 -158 512 -128
rect 686 -158 714 -100
rect 506 -180 714 -158
rect 446 -186 714 -180
rect 786 -336 814 290
rect 786 -344 1098 -336
rect 786 -372 1037 -344
rect 446 -560 522 -554
rect 446 -586 454 -560
rect -127 -644 -126 -604
rect 354 -612 454 -586
rect 506 -612 522 -560
rect 354 -614 522 -612
rect 446 -618 522 -614
rect -180 -660 -126 -644
rect 786 -776 814 -372
rect 1018 -396 1037 -372
rect 1089 -396 1098 -344
rect 1018 -408 1098 -396
rect 162 -804 814 -776
rect 940 -1004 1290 -990
rect 940 -1120 961 -1004
rect 1269 -1120 1290 -1004
rect 940 -1134 1290 -1120
<< via2 >>
rect 967 1034 1023 1090
rect 1047 1034 1103 1090
rect 1127 1034 1183 1090
rect 1207 1034 1263 1090
rect 967 -1090 1023 -1034
rect 1047 -1090 1103 -1034
rect 1127 -1090 1183 -1034
rect 1207 -1090 1263 -1034
<< metal3 >>
rect -574 1090 1322 1192
rect -574 1034 967 1090
rect 1023 1034 1047 1090
rect 1103 1034 1127 1090
rect 1183 1034 1207 1090
rect 1263 1034 1322 1090
rect -574 938 1322 1034
rect -566 -1034 1322 -930
rect -566 -1090 967 -1034
rect 1023 -1090 1047 -1034
rect 1103 -1090 1127 -1034
rect 1183 -1090 1207 -1034
rect 1263 -1090 1322 -1034
rect -566 -1185 1322 -1090
use sky130_fd_pr__pfet_01v8_hvt_UUWA33  1
timestamp 1655322987
transform 1 0 -125 0 1 -222
box -109 -200 109 200
use sky130_fd_pr__pfet_01v8_hvt_UUWA33  2
timestamp 1655322987
transform 1 0 521 0 1 -222
box -109 -200 109 200
use demux  demux_0
timestamp 1655348380
transform 1 0 36 0 1 156
box -76 -122 336 878
use mux  mux_0
timestamp 1655348380
transform 1 0 34 0 1 -900
box -54 -122 366 878
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_0
timestamp 1655322987
transform 1 0 1008 0 1 -606
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1#0  sky130_fd_sc_hd__inv_1_0
timestamp 1655322987
transform 1 0 662 0 1 -604
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1#0  sky130_fd_sc_hd__inv_1_1
timestamp 1655322987
transform 1 0 -534 0 1 -612
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_0
timestamp 1655322987
transform 1 0 -366 0 1 442
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_1
timestamp 1655322987
transform 1 0 458 0 1 442
box -38 -48 314 592
<< labels >>
flabel metal2 s -514 304 -450 312 1 FreeSans 625 0 0 0 IN
port 1 nsew
flabel metal2 s -554 -896 -510 -852 1 FreeSans 625 0 0 0 C
port 2 nsew
flabel metal1 s -438 -834 -394 -778 1 FreeSans 625 0 0 0 VSS
port 3 nsew
flabel metal3 s -484 1060 -440 1116 1 FreeSans 625 0 0 0 VDD
port 4 nsew
flabel metal2 s 1194 306 1258 314 1 FreeSans 625 0 0 0 OUT
port 5 nsew
flabel metal1 s 1246 -392 1290 -336 1 FreeSans 625 0 0 0 buf_out
port 6 nsew
<< end >>
