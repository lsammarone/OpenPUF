magic
tech sky130A
magscale 1 2
timestamp 1656729169
<< nwell >>
rect 120 1707 27826 1940
rect 120 294 27827 1707
rect 217 293 27827 294
<< pmoslvt >>
rect 311 355 711 1645
rect 769 355 1169 1645
rect 1227 355 1627 1645
rect 1685 355 2085 1645
rect 2143 355 2543 1645
rect 2601 355 3001 1645
rect 3059 355 3459 1645
rect 3517 355 3917 1645
rect 3975 355 4375 1645
rect 4433 355 4833 1645
rect 4891 355 5291 1645
rect 5349 355 5749 1645
rect 5807 355 6207 1645
rect 6265 355 6665 1645
rect 6723 355 7123 1645
rect 7181 355 7581 1645
rect 7639 355 8039 1645
rect 8097 355 8497 1645
rect 8555 355 8955 1645
rect 9013 355 9413 1645
rect 9471 355 9871 1645
rect 9929 355 10329 1645
rect 10387 355 10787 1645
rect 10845 355 11245 1645
rect 11303 355 11703 1645
rect 11761 355 12161 1645
rect 12219 355 12619 1645
rect 12677 355 13077 1645
rect 13135 355 13535 1645
rect 13593 355 13993 1645
rect 14051 355 14451 1645
rect 14509 355 14909 1645
rect 14967 355 15367 1645
rect 15425 355 15825 1645
rect 15883 355 16283 1645
rect 16341 355 16741 1645
rect 16799 355 17199 1645
rect 17257 355 17657 1645
rect 17715 355 18115 1645
rect 18173 355 18573 1645
rect 18631 355 19031 1645
rect 19089 355 19489 1645
rect 19547 355 19947 1645
rect 20005 355 20405 1645
rect 20463 355 20863 1645
rect 20921 355 21321 1645
rect 21379 355 21779 1645
rect 21837 355 22237 1645
rect 22295 355 22695 1645
rect 22753 355 23153 1645
rect 23211 355 23611 1645
rect 23669 355 24069 1645
rect 24127 355 24527 1645
rect 24585 355 24985 1645
rect 25043 355 25443 1645
rect 25501 355 25901 1645
rect 25959 355 26359 1645
rect 26417 355 26817 1645
rect 26875 355 27275 1645
rect 27333 355 27733 1645
<< pdiff >>
rect 253 1629 311 1645
rect 253 1595 265 1629
rect 299 1595 311 1629
rect 253 1561 311 1595
rect 253 1527 265 1561
rect 299 1527 311 1561
rect 253 1493 311 1527
rect 253 1459 265 1493
rect 299 1459 311 1493
rect 253 1425 311 1459
rect 253 1391 265 1425
rect 299 1391 311 1425
rect 253 1357 311 1391
rect 253 1323 265 1357
rect 299 1323 311 1357
rect 253 1289 311 1323
rect 253 1255 265 1289
rect 299 1255 311 1289
rect 253 1221 311 1255
rect 253 1187 265 1221
rect 299 1187 311 1221
rect 253 1153 311 1187
rect 253 1119 265 1153
rect 299 1119 311 1153
rect 253 1085 311 1119
rect 253 1051 265 1085
rect 299 1051 311 1085
rect 253 1017 311 1051
rect 253 983 265 1017
rect 299 983 311 1017
rect 253 949 311 983
rect 253 915 265 949
rect 299 915 311 949
rect 253 881 311 915
rect 253 847 265 881
rect 299 847 311 881
rect 253 813 311 847
rect 253 779 265 813
rect 299 779 311 813
rect 253 745 311 779
rect 253 711 265 745
rect 299 711 311 745
rect 253 677 311 711
rect 253 643 265 677
rect 299 643 311 677
rect 253 609 311 643
rect 253 575 265 609
rect 299 575 311 609
rect 253 541 311 575
rect 253 507 265 541
rect 299 507 311 541
rect 253 473 311 507
rect 253 439 265 473
rect 299 439 311 473
rect 253 405 311 439
rect 253 371 265 405
rect 299 371 311 405
rect 253 355 311 371
rect 711 1629 769 1645
rect 711 1595 723 1629
rect 757 1595 769 1629
rect 711 1561 769 1595
rect 711 1527 723 1561
rect 757 1527 769 1561
rect 711 1493 769 1527
rect 711 1459 723 1493
rect 757 1459 769 1493
rect 711 1425 769 1459
rect 711 1391 723 1425
rect 757 1391 769 1425
rect 711 1357 769 1391
rect 711 1323 723 1357
rect 757 1323 769 1357
rect 711 1289 769 1323
rect 711 1255 723 1289
rect 757 1255 769 1289
rect 711 1221 769 1255
rect 711 1187 723 1221
rect 757 1187 769 1221
rect 711 1153 769 1187
rect 711 1119 723 1153
rect 757 1119 769 1153
rect 711 1085 769 1119
rect 711 1051 723 1085
rect 757 1051 769 1085
rect 711 1017 769 1051
rect 711 983 723 1017
rect 757 983 769 1017
rect 711 949 769 983
rect 711 915 723 949
rect 757 915 769 949
rect 711 881 769 915
rect 711 847 723 881
rect 757 847 769 881
rect 711 813 769 847
rect 711 779 723 813
rect 757 779 769 813
rect 711 745 769 779
rect 711 711 723 745
rect 757 711 769 745
rect 711 677 769 711
rect 711 643 723 677
rect 757 643 769 677
rect 711 609 769 643
rect 711 575 723 609
rect 757 575 769 609
rect 711 541 769 575
rect 711 507 723 541
rect 757 507 769 541
rect 711 473 769 507
rect 711 439 723 473
rect 757 439 769 473
rect 711 405 769 439
rect 711 371 723 405
rect 757 371 769 405
rect 711 355 769 371
rect 1169 1629 1227 1645
rect 1169 1595 1181 1629
rect 1215 1595 1227 1629
rect 1169 1561 1227 1595
rect 1169 1527 1181 1561
rect 1215 1527 1227 1561
rect 1169 1493 1227 1527
rect 1169 1459 1181 1493
rect 1215 1459 1227 1493
rect 1169 1425 1227 1459
rect 1169 1391 1181 1425
rect 1215 1391 1227 1425
rect 1169 1357 1227 1391
rect 1169 1323 1181 1357
rect 1215 1323 1227 1357
rect 1169 1289 1227 1323
rect 1169 1255 1181 1289
rect 1215 1255 1227 1289
rect 1169 1221 1227 1255
rect 1169 1187 1181 1221
rect 1215 1187 1227 1221
rect 1169 1153 1227 1187
rect 1169 1119 1181 1153
rect 1215 1119 1227 1153
rect 1169 1085 1227 1119
rect 1169 1051 1181 1085
rect 1215 1051 1227 1085
rect 1169 1017 1227 1051
rect 1169 983 1181 1017
rect 1215 983 1227 1017
rect 1169 949 1227 983
rect 1169 915 1181 949
rect 1215 915 1227 949
rect 1169 881 1227 915
rect 1169 847 1181 881
rect 1215 847 1227 881
rect 1169 813 1227 847
rect 1169 779 1181 813
rect 1215 779 1227 813
rect 1169 745 1227 779
rect 1169 711 1181 745
rect 1215 711 1227 745
rect 1169 677 1227 711
rect 1169 643 1181 677
rect 1215 643 1227 677
rect 1169 609 1227 643
rect 1169 575 1181 609
rect 1215 575 1227 609
rect 1169 541 1227 575
rect 1169 507 1181 541
rect 1215 507 1227 541
rect 1169 473 1227 507
rect 1169 439 1181 473
rect 1215 439 1227 473
rect 1169 405 1227 439
rect 1169 371 1181 405
rect 1215 371 1227 405
rect 1169 355 1227 371
rect 1627 1629 1685 1645
rect 1627 1595 1639 1629
rect 1673 1595 1685 1629
rect 1627 1561 1685 1595
rect 1627 1527 1639 1561
rect 1673 1527 1685 1561
rect 1627 1493 1685 1527
rect 1627 1459 1639 1493
rect 1673 1459 1685 1493
rect 1627 1425 1685 1459
rect 1627 1391 1639 1425
rect 1673 1391 1685 1425
rect 1627 1357 1685 1391
rect 1627 1323 1639 1357
rect 1673 1323 1685 1357
rect 1627 1289 1685 1323
rect 1627 1255 1639 1289
rect 1673 1255 1685 1289
rect 1627 1221 1685 1255
rect 1627 1187 1639 1221
rect 1673 1187 1685 1221
rect 1627 1153 1685 1187
rect 1627 1119 1639 1153
rect 1673 1119 1685 1153
rect 1627 1085 1685 1119
rect 1627 1051 1639 1085
rect 1673 1051 1685 1085
rect 1627 1017 1685 1051
rect 1627 983 1639 1017
rect 1673 983 1685 1017
rect 1627 949 1685 983
rect 1627 915 1639 949
rect 1673 915 1685 949
rect 1627 881 1685 915
rect 1627 847 1639 881
rect 1673 847 1685 881
rect 1627 813 1685 847
rect 1627 779 1639 813
rect 1673 779 1685 813
rect 1627 745 1685 779
rect 1627 711 1639 745
rect 1673 711 1685 745
rect 1627 677 1685 711
rect 1627 643 1639 677
rect 1673 643 1685 677
rect 1627 609 1685 643
rect 1627 575 1639 609
rect 1673 575 1685 609
rect 1627 541 1685 575
rect 1627 507 1639 541
rect 1673 507 1685 541
rect 1627 473 1685 507
rect 1627 439 1639 473
rect 1673 439 1685 473
rect 1627 405 1685 439
rect 1627 371 1639 405
rect 1673 371 1685 405
rect 1627 355 1685 371
rect 2085 1629 2143 1645
rect 2085 1595 2097 1629
rect 2131 1595 2143 1629
rect 2085 1561 2143 1595
rect 2085 1527 2097 1561
rect 2131 1527 2143 1561
rect 2085 1493 2143 1527
rect 2085 1459 2097 1493
rect 2131 1459 2143 1493
rect 2085 1425 2143 1459
rect 2085 1391 2097 1425
rect 2131 1391 2143 1425
rect 2085 1357 2143 1391
rect 2085 1323 2097 1357
rect 2131 1323 2143 1357
rect 2085 1289 2143 1323
rect 2085 1255 2097 1289
rect 2131 1255 2143 1289
rect 2085 1221 2143 1255
rect 2085 1187 2097 1221
rect 2131 1187 2143 1221
rect 2085 1153 2143 1187
rect 2085 1119 2097 1153
rect 2131 1119 2143 1153
rect 2085 1085 2143 1119
rect 2085 1051 2097 1085
rect 2131 1051 2143 1085
rect 2085 1017 2143 1051
rect 2085 983 2097 1017
rect 2131 983 2143 1017
rect 2085 949 2143 983
rect 2085 915 2097 949
rect 2131 915 2143 949
rect 2085 881 2143 915
rect 2085 847 2097 881
rect 2131 847 2143 881
rect 2085 813 2143 847
rect 2085 779 2097 813
rect 2131 779 2143 813
rect 2085 745 2143 779
rect 2085 711 2097 745
rect 2131 711 2143 745
rect 2085 677 2143 711
rect 2085 643 2097 677
rect 2131 643 2143 677
rect 2085 609 2143 643
rect 2085 575 2097 609
rect 2131 575 2143 609
rect 2085 541 2143 575
rect 2085 507 2097 541
rect 2131 507 2143 541
rect 2085 473 2143 507
rect 2085 439 2097 473
rect 2131 439 2143 473
rect 2085 405 2143 439
rect 2085 371 2097 405
rect 2131 371 2143 405
rect 2085 355 2143 371
rect 2543 1629 2601 1645
rect 2543 1595 2555 1629
rect 2589 1595 2601 1629
rect 2543 1561 2601 1595
rect 2543 1527 2555 1561
rect 2589 1527 2601 1561
rect 2543 1493 2601 1527
rect 2543 1459 2555 1493
rect 2589 1459 2601 1493
rect 2543 1425 2601 1459
rect 2543 1391 2555 1425
rect 2589 1391 2601 1425
rect 2543 1357 2601 1391
rect 2543 1323 2555 1357
rect 2589 1323 2601 1357
rect 2543 1289 2601 1323
rect 2543 1255 2555 1289
rect 2589 1255 2601 1289
rect 2543 1221 2601 1255
rect 2543 1187 2555 1221
rect 2589 1187 2601 1221
rect 2543 1153 2601 1187
rect 2543 1119 2555 1153
rect 2589 1119 2601 1153
rect 2543 1085 2601 1119
rect 2543 1051 2555 1085
rect 2589 1051 2601 1085
rect 2543 1017 2601 1051
rect 2543 983 2555 1017
rect 2589 983 2601 1017
rect 2543 949 2601 983
rect 2543 915 2555 949
rect 2589 915 2601 949
rect 2543 881 2601 915
rect 2543 847 2555 881
rect 2589 847 2601 881
rect 2543 813 2601 847
rect 2543 779 2555 813
rect 2589 779 2601 813
rect 2543 745 2601 779
rect 2543 711 2555 745
rect 2589 711 2601 745
rect 2543 677 2601 711
rect 2543 643 2555 677
rect 2589 643 2601 677
rect 2543 609 2601 643
rect 2543 575 2555 609
rect 2589 575 2601 609
rect 2543 541 2601 575
rect 2543 507 2555 541
rect 2589 507 2601 541
rect 2543 473 2601 507
rect 2543 439 2555 473
rect 2589 439 2601 473
rect 2543 405 2601 439
rect 2543 371 2555 405
rect 2589 371 2601 405
rect 2543 355 2601 371
rect 3001 1629 3059 1645
rect 3001 1595 3013 1629
rect 3047 1595 3059 1629
rect 3001 1561 3059 1595
rect 3001 1527 3013 1561
rect 3047 1527 3059 1561
rect 3001 1493 3059 1527
rect 3001 1459 3013 1493
rect 3047 1459 3059 1493
rect 3001 1425 3059 1459
rect 3001 1391 3013 1425
rect 3047 1391 3059 1425
rect 3001 1357 3059 1391
rect 3001 1323 3013 1357
rect 3047 1323 3059 1357
rect 3001 1289 3059 1323
rect 3001 1255 3013 1289
rect 3047 1255 3059 1289
rect 3001 1221 3059 1255
rect 3001 1187 3013 1221
rect 3047 1187 3059 1221
rect 3001 1153 3059 1187
rect 3001 1119 3013 1153
rect 3047 1119 3059 1153
rect 3001 1085 3059 1119
rect 3001 1051 3013 1085
rect 3047 1051 3059 1085
rect 3001 1017 3059 1051
rect 3001 983 3013 1017
rect 3047 983 3059 1017
rect 3001 949 3059 983
rect 3001 915 3013 949
rect 3047 915 3059 949
rect 3001 881 3059 915
rect 3001 847 3013 881
rect 3047 847 3059 881
rect 3001 813 3059 847
rect 3001 779 3013 813
rect 3047 779 3059 813
rect 3001 745 3059 779
rect 3001 711 3013 745
rect 3047 711 3059 745
rect 3001 677 3059 711
rect 3001 643 3013 677
rect 3047 643 3059 677
rect 3001 609 3059 643
rect 3001 575 3013 609
rect 3047 575 3059 609
rect 3001 541 3059 575
rect 3001 507 3013 541
rect 3047 507 3059 541
rect 3001 473 3059 507
rect 3001 439 3013 473
rect 3047 439 3059 473
rect 3001 405 3059 439
rect 3001 371 3013 405
rect 3047 371 3059 405
rect 3001 355 3059 371
rect 3459 1629 3517 1645
rect 3459 1595 3471 1629
rect 3505 1595 3517 1629
rect 3459 1561 3517 1595
rect 3459 1527 3471 1561
rect 3505 1527 3517 1561
rect 3459 1493 3517 1527
rect 3459 1459 3471 1493
rect 3505 1459 3517 1493
rect 3459 1425 3517 1459
rect 3459 1391 3471 1425
rect 3505 1391 3517 1425
rect 3459 1357 3517 1391
rect 3459 1323 3471 1357
rect 3505 1323 3517 1357
rect 3459 1289 3517 1323
rect 3459 1255 3471 1289
rect 3505 1255 3517 1289
rect 3459 1221 3517 1255
rect 3459 1187 3471 1221
rect 3505 1187 3517 1221
rect 3459 1153 3517 1187
rect 3459 1119 3471 1153
rect 3505 1119 3517 1153
rect 3459 1085 3517 1119
rect 3459 1051 3471 1085
rect 3505 1051 3517 1085
rect 3459 1017 3517 1051
rect 3459 983 3471 1017
rect 3505 983 3517 1017
rect 3459 949 3517 983
rect 3459 915 3471 949
rect 3505 915 3517 949
rect 3459 881 3517 915
rect 3459 847 3471 881
rect 3505 847 3517 881
rect 3459 813 3517 847
rect 3459 779 3471 813
rect 3505 779 3517 813
rect 3459 745 3517 779
rect 3459 711 3471 745
rect 3505 711 3517 745
rect 3459 677 3517 711
rect 3459 643 3471 677
rect 3505 643 3517 677
rect 3459 609 3517 643
rect 3459 575 3471 609
rect 3505 575 3517 609
rect 3459 541 3517 575
rect 3459 507 3471 541
rect 3505 507 3517 541
rect 3459 473 3517 507
rect 3459 439 3471 473
rect 3505 439 3517 473
rect 3459 405 3517 439
rect 3459 371 3471 405
rect 3505 371 3517 405
rect 3459 355 3517 371
rect 3917 1629 3975 1645
rect 3917 1595 3929 1629
rect 3963 1595 3975 1629
rect 3917 1561 3975 1595
rect 3917 1527 3929 1561
rect 3963 1527 3975 1561
rect 3917 1493 3975 1527
rect 3917 1459 3929 1493
rect 3963 1459 3975 1493
rect 3917 1425 3975 1459
rect 3917 1391 3929 1425
rect 3963 1391 3975 1425
rect 3917 1357 3975 1391
rect 3917 1323 3929 1357
rect 3963 1323 3975 1357
rect 3917 1289 3975 1323
rect 3917 1255 3929 1289
rect 3963 1255 3975 1289
rect 3917 1221 3975 1255
rect 3917 1187 3929 1221
rect 3963 1187 3975 1221
rect 3917 1153 3975 1187
rect 3917 1119 3929 1153
rect 3963 1119 3975 1153
rect 3917 1085 3975 1119
rect 3917 1051 3929 1085
rect 3963 1051 3975 1085
rect 3917 1017 3975 1051
rect 3917 983 3929 1017
rect 3963 983 3975 1017
rect 3917 949 3975 983
rect 3917 915 3929 949
rect 3963 915 3975 949
rect 3917 881 3975 915
rect 3917 847 3929 881
rect 3963 847 3975 881
rect 3917 813 3975 847
rect 3917 779 3929 813
rect 3963 779 3975 813
rect 3917 745 3975 779
rect 3917 711 3929 745
rect 3963 711 3975 745
rect 3917 677 3975 711
rect 3917 643 3929 677
rect 3963 643 3975 677
rect 3917 609 3975 643
rect 3917 575 3929 609
rect 3963 575 3975 609
rect 3917 541 3975 575
rect 3917 507 3929 541
rect 3963 507 3975 541
rect 3917 473 3975 507
rect 3917 439 3929 473
rect 3963 439 3975 473
rect 3917 405 3975 439
rect 3917 371 3929 405
rect 3963 371 3975 405
rect 3917 355 3975 371
rect 4375 1629 4433 1645
rect 4375 1595 4387 1629
rect 4421 1595 4433 1629
rect 4375 1561 4433 1595
rect 4375 1527 4387 1561
rect 4421 1527 4433 1561
rect 4375 1493 4433 1527
rect 4375 1459 4387 1493
rect 4421 1459 4433 1493
rect 4375 1425 4433 1459
rect 4375 1391 4387 1425
rect 4421 1391 4433 1425
rect 4375 1357 4433 1391
rect 4375 1323 4387 1357
rect 4421 1323 4433 1357
rect 4375 1289 4433 1323
rect 4375 1255 4387 1289
rect 4421 1255 4433 1289
rect 4375 1221 4433 1255
rect 4375 1187 4387 1221
rect 4421 1187 4433 1221
rect 4375 1153 4433 1187
rect 4375 1119 4387 1153
rect 4421 1119 4433 1153
rect 4375 1085 4433 1119
rect 4375 1051 4387 1085
rect 4421 1051 4433 1085
rect 4375 1017 4433 1051
rect 4375 983 4387 1017
rect 4421 983 4433 1017
rect 4375 949 4433 983
rect 4375 915 4387 949
rect 4421 915 4433 949
rect 4375 881 4433 915
rect 4375 847 4387 881
rect 4421 847 4433 881
rect 4375 813 4433 847
rect 4375 779 4387 813
rect 4421 779 4433 813
rect 4375 745 4433 779
rect 4375 711 4387 745
rect 4421 711 4433 745
rect 4375 677 4433 711
rect 4375 643 4387 677
rect 4421 643 4433 677
rect 4375 609 4433 643
rect 4375 575 4387 609
rect 4421 575 4433 609
rect 4375 541 4433 575
rect 4375 507 4387 541
rect 4421 507 4433 541
rect 4375 473 4433 507
rect 4375 439 4387 473
rect 4421 439 4433 473
rect 4375 405 4433 439
rect 4375 371 4387 405
rect 4421 371 4433 405
rect 4375 355 4433 371
rect 4833 1629 4891 1645
rect 4833 1595 4845 1629
rect 4879 1595 4891 1629
rect 4833 1561 4891 1595
rect 4833 1527 4845 1561
rect 4879 1527 4891 1561
rect 4833 1493 4891 1527
rect 4833 1459 4845 1493
rect 4879 1459 4891 1493
rect 4833 1425 4891 1459
rect 4833 1391 4845 1425
rect 4879 1391 4891 1425
rect 4833 1357 4891 1391
rect 4833 1323 4845 1357
rect 4879 1323 4891 1357
rect 4833 1289 4891 1323
rect 4833 1255 4845 1289
rect 4879 1255 4891 1289
rect 4833 1221 4891 1255
rect 4833 1187 4845 1221
rect 4879 1187 4891 1221
rect 4833 1153 4891 1187
rect 4833 1119 4845 1153
rect 4879 1119 4891 1153
rect 4833 1085 4891 1119
rect 4833 1051 4845 1085
rect 4879 1051 4891 1085
rect 4833 1017 4891 1051
rect 4833 983 4845 1017
rect 4879 983 4891 1017
rect 4833 949 4891 983
rect 4833 915 4845 949
rect 4879 915 4891 949
rect 4833 881 4891 915
rect 4833 847 4845 881
rect 4879 847 4891 881
rect 4833 813 4891 847
rect 4833 779 4845 813
rect 4879 779 4891 813
rect 4833 745 4891 779
rect 4833 711 4845 745
rect 4879 711 4891 745
rect 4833 677 4891 711
rect 4833 643 4845 677
rect 4879 643 4891 677
rect 4833 609 4891 643
rect 4833 575 4845 609
rect 4879 575 4891 609
rect 4833 541 4891 575
rect 4833 507 4845 541
rect 4879 507 4891 541
rect 4833 473 4891 507
rect 4833 439 4845 473
rect 4879 439 4891 473
rect 4833 405 4891 439
rect 4833 371 4845 405
rect 4879 371 4891 405
rect 4833 355 4891 371
rect 5291 1629 5349 1645
rect 5291 1595 5303 1629
rect 5337 1595 5349 1629
rect 5291 1561 5349 1595
rect 5291 1527 5303 1561
rect 5337 1527 5349 1561
rect 5291 1493 5349 1527
rect 5291 1459 5303 1493
rect 5337 1459 5349 1493
rect 5291 1425 5349 1459
rect 5291 1391 5303 1425
rect 5337 1391 5349 1425
rect 5291 1357 5349 1391
rect 5291 1323 5303 1357
rect 5337 1323 5349 1357
rect 5291 1289 5349 1323
rect 5291 1255 5303 1289
rect 5337 1255 5349 1289
rect 5291 1221 5349 1255
rect 5291 1187 5303 1221
rect 5337 1187 5349 1221
rect 5291 1153 5349 1187
rect 5291 1119 5303 1153
rect 5337 1119 5349 1153
rect 5291 1085 5349 1119
rect 5291 1051 5303 1085
rect 5337 1051 5349 1085
rect 5291 1017 5349 1051
rect 5291 983 5303 1017
rect 5337 983 5349 1017
rect 5291 949 5349 983
rect 5291 915 5303 949
rect 5337 915 5349 949
rect 5291 881 5349 915
rect 5291 847 5303 881
rect 5337 847 5349 881
rect 5291 813 5349 847
rect 5291 779 5303 813
rect 5337 779 5349 813
rect 5291 745 5349 779
rect 5291 711 5303 745
rect 5337 711 5349 745
rect 5291 677 5349 711
rect 5291 643 5303 677
rect 5337 643 5349 677
rect 5291 609 5349 643
rect 5291 575 5303 609
rect 5337 575 5349 609
rect 5291 541 5349 575
rect 5291 507 5303 541
rect 5337 507 5349 541
rect 5291 473 5349 507
rect 5291 439 5303 473
rect 5337 439 5349 473
rect 5291 405 5349 439
rect 5291 371 5303 405
rect 5337 371 5349 405
rect 5291 355 5349 371
rect 5749 1629 5807 1645
rect 5749 1595 5761 1629
rect 5795 1595 5807 1629
rect 5749 1561 5807 1595
rect 5749 1527 5761 1561
rect 5795 1527 5807 1561
rect 5749 1493 5807 1527
rect 5749 1459 5761 1493
rect 5795 1459 5807 1493
rect 5749 1425 5807 1459
rect 5749 1391 5761 1425
rect 5795 1391 5807 1425
rect 5749 1357 5807 1391
rect 5749 1323 5761 1357
rect 5795 1323 5807 1357
rect 5749 1289 5807 1323
rect 5749 1255 5761 1289
rect 5795 1255 5807 1289
rect 5749 1221 5807 1255
rect 5749 1187 5761 1221
rect 5795 1187 5807 1221
rect 5749 1153 5807 1187
rect 5749 1119 5761 1153
rect 5795 1119 5807 1153
rect 5749 1085 5807 1119
rect 5749 1051 5761 1085
rect 5795 1051 5807 1085
rect 5749 1017 5807 1051
rect 5749 983 5761 1017
rect 5795 983 5807 1017
rect 5749 949 5807 983
rect 5749 915 5761 949
rect 5795 915 5807 949
rect 5749 881 5807 915
rect 5749 847 5761 881
rect 5795 847 5807 881
rect 5749 813 5807 847
rect 5749 779 5761 813
rect 5795 779 5807 813
rect 5749 745 5807 779
rect 5749 711 5761 745
rect 5795 711 5807 745
rect 5749 677 5807 711
rect 5749 643 5761 677
rect 5795 643 5807 677
rect 5749 609 5807 643
rect 5749 575 5761 609
rect 5795 575 5807 609
rect 5749 541 5807 575
rect 5749 507 5761 541
rect 5795 507 5807 541
rect 5749 473 5807 507
rect 5749 439 5761 473
rect 5795 439 5807 473
rect 5749 405 5807 439
rect 5749 371 5761 405
rect 5795 371 5807 405
rect 5749 355 5807 371
rect 6207 1629 6265 1645
rect 6207 1595 6219 1629
rect 6253 1595 6265 1629
rect 6207 1561 6265 1595
rect 6207 1527 6219 1561
rect 6253 1527 6265 1561
rect 6207 1493 6265 1527
rect 6207 1459 6219 1493
rect 6253 1459 6265 1493
rect 6207 1425 6265 1459
rect 6207 1391 6219 1425
rect 6253 1391 6265 1425
rect 6207 1357 6265 1391
rect 6207 1323 6219 1357
rect 6253 1323 6265 1357
rect 6207 1289 6265 1323
rect 6207 1255 6219 1289
rect 6253 1255 6265 1289
rect 6207 1221 6265 1255
rect 6207 1187 6219 1221
rect 6253 1187 6265 1221
rect 6207 1153 6265 1187
rect 6207 1119 6219 1153
rect 6253 1119 6265 1153
rect 6207 1085 6265 1119
rect 6207 1051 6219 1085
rect 6253 1051 6265 1085
rect 6207 1017 6265 1051
rect 6207 983 6219 1017
rect 6253 983 6265 1017
rect 6207 949 6265 983
rect 6207 915 6219 949
rect 6253 915 6265 949
rect 6207 881 6265 915
rect 6207 847 6219 881
rect 6253 847 6265 881
rect 6207 813 6265 847
rect 6207 779 6219 813
rect 6253 779 6265 813
rect 6207 745 6265 779
rect 6207 711 6219 745
rect 6253 711 6265 745
rect 6207 677 6265 711
rect 6207 643 6219 677
rect 6253 643 6265 677
rect 6207 609 6265 643
rect 6207 575 6219 609
rect 6253 575 6265 609
rect 6207 541 6265 575
rect 6207 507 6219 541
rect 6253 507 6265 541
rect 6207 473 6265 507
rect 6207 439 6219 473
rect 6253 439 6265 473
rect 6207 405 6265 439
rect 6207 371 6219 405
rect 6253 371 6265 405
rect 6207 355 6265 371
rect 6665 1629 6723 1645
rect 6665 1595 6677 1629
rect 6711 1595 6723 1629
rect 6665 1561 6723 1595
rect 6665 1527 6677 1561
rect 6711 1527 6723 1561
rect 6665 1493 6723 1527
rect 6665 1459 6677 1493
rect 6711 1459 6723 1493
rect 6665 1425 6723 1459
rect 6665 1391 6677 1425
rect 6711 1391 6723 1425
rect 6665 1357 6723 1391
rect 6665 1323 6677 1357
rect 6711 1323 6723 1357
rect 6665 1289 6723 1323
rect 6665 1255 6677 1289
rect 6711 1255 6723 1289
rect 6665 1221 6723 1255
rect 6665 1187 6677 1221
rect 6711 1187 6723 1221
rect 6665 1153 6723 1187
rect 6665 1119 6677 1153
rect 6711 1119 6723 1153
rect 6665 1085 6723 1119
rect 6665 1051 6677 1085
rect 6711 1051 6723 1085
rect 6665 1017 6723 1051
rect 6665 983 6677 1017
rect 6711 983 6723 1017
rect 6665 949 6723 983
rect 6665 915 6677 949
rect 6711 915 6723 949
rect 6665 881 6723 915
rect 6665 847 6677 881
rect 6711 847 6723 881
rect 6665 813 6723 847
rect 6665 779 6677 813
rect 6711 779 6723 813
rect 6665 745 6723 779
rect 6665 711 6677 745
rect 6711 711 6723 745
rect 6665 677 6723 711
rect 6665 643 6677 677
rect 6711 643 6723 677
rect 6665 609 6723 643
rect 6665 575 6677 609
rect 6711 575 6723 609
rect 6665 541 6723 575
rect 6665 507 6677 541
rect 6711 507 6723 541
rect 6665 473 6723 507
rect 6665 439 6677 473
rect 6711 439 6723 473
rect 6665 405 6723 439
rect 6665 371 6677 405
rect 6711 371 6723 405
rect 6665 355 6723 371
rect 7123 1629 7181 1645
rect 7123 1595 7135 1629
rect 7169 1595 7181 1629
rect 7123 1561 7181 1595
rect 7123 1527 7135 1561
rect 7169 1527 7181 1561
rect 7123 1493 7181 1527
rect 7123 1459 7135 1493
rect 7169 1459 7181 1493
rect 7123 1425 7181 1459
rect 7123 1391 7135 1425
rect 7169 1391 7181 1425
rect 7123 1357 7181 1391
rect 7123 1323 7135 1357
rect 7169 1323 7181 1357
rect 7123 1289 7181 1323
rect 7123 1255 7135 1289
rect 7169 1255 7181 1289
rect 7123 1221 7181 1255
rect 7123 1187 7135 1221
rect 7169 1187 7181 1221
rect 7123 1153 7181 1187
rect 7123 1119 7135 1153
rect 7169 1119 7181 1153
rect 7123 1085 7181 1119
rect 7123 1051 7135 1085
rect 7169 1051 7181 1085
rect 7123 1017 7181 1051
rect 7123 983 7135 1017
rect 7169 983 7181 1017
rect 7123 949 7181 983
rect 7123 915 7135 949
rect 7169 915 7181 949
rect 7123 881 7181 915
rect 7123 847 7135 881
rect 7169 847 7181 881
rect 7123 813 7181 847
rect 7123 779 7135 813
rect 7169 779 7181 813
rect 7123 745 7181 779
rect 7123 711 7135 745
rect 7169 711 7181 745
rect 7123 677 7181 711
rect 7123 643 7135 677
rect 7169 643 7181 677
rect 7123 609 7181 643
rect 7123 575 7135 609
rect 7169 575 7181 609
rect 7123 541 7181 575
rect 7123 507 7135 541
rect 7169 507 7181 541
rect 7123 473 7181 507
rect 7123 439 7135 473
rect 7169 439 7181 473
rect 7123 405 7181 439
rect 7123 371 7135 405
rect 7169 371 7181 405
rect 7123 355 7181 371
rect 7581 1629 7639 1645
rect 7581 1595 7593 1629
rect 7627 1595 7639 1629
rect 7581 1561 7639 1595
rect 7581 1527 7593 1561
rect 7627 1527 7639 1561
rect 7581 1493 7639 1527
rect 7581 1459 7593 1493
rect 7627 1459 7639 1493
rect 7581 1425 7639 1459
rect 7581 1391 7593 1425
rect 7627 1391 7639 1425
rect 7581 1357 7639 1391
rect 7581 1323 7593 1357
rect 7627 1323 7639 1357
rect 7581 1289 7639 1323
rect 7581 1255 7593 1289
rect 7627 1255 7639 1289
rect 7581 1221 7639 1255
rect 7581 1187 7593 1221
rect 7627 1187 7639 1221
rect 7581 1153 7639 1187
rect 7581 1119 7593 1153
rect 7627 1119 7639 1153
rect 7581 1085 7639 1119
rect 7581 1051 7593 1085
rect 7627 1051 7639 1085
rect 7581 1017 7639 1051
rect 7581 983 7593 1017
rect 7627 983 7639 1017
rect 7581 949 7639 983
rect 7581 915 7593 949
rect 7627 915 7639 949
rect 7581 881 7639 915
rect 7581 847 7593 881
rect 7627 847 7639 881
rect 7581 813 7639 847
rect 7581 779 7593 813
rect 7627 779 7639 813
rect 7581 745 7639 779
rect 7581 711 7593 745
rect 7627 711 7639 745
rect 7581 677 7639 711
rect 7581 643 7593 677
rect 7627 643 7639 677
rect 7581 609 7639 643
rect 7581 575 7593 609
rect 7627 575 7639 609
rect 7581 541 7639 575
rect 7581 507 7593 541
rect 7627 507 7639 541
rect 7581 473 7639 507
rect 7581 439 7593 473
rect 7627 439 7639 473
rect 7581 405 7639 439
rect 7581 371 7593 405
rect 7627 371 7639 405
rect 7581 355 7639 371
rect 8039 1629 8097 1645
rect 8039 1595 8051 1629
rect 8085 1595 8097 1629
rect 8039 1561 8097 1595
rect 8039 1527 8051 1561
rect 8085 1527 8097 1561
rect 8039 1493 8097 1527
rect 8039 1459 8051 1493
rect 8085 1459 8097 1493
rect 8039 1425 8097 1459
rect 8039 1391 8051 1425
rect 8085 1391 8097 1425
rect 8039 1357 8097 1391
rect 8039 1323 8051 1357
rect 8085 1323 8097 1357
rect 8039 1289 8097 1323
rect 8039 1255 8051 1289
rect 8085 1255 8097 1289
rect 8039 1221 8097 1255
rect 8039 1187 8051 1221
rect 8085 1187 8097 1221
rect 8039 1153 8097 1187
rect 8039 1119 8051 1153
rect 8085 1119 8097 1153
rect 8039 1085 8097 1119
rect 8039 1051 8051 1085
rect 8085 1051 8097 1085
rect 8039 1017 8097 1051
rect 8039 983 8051 1017
rect 8085 983 8097 1017
rect 8039 949 8097 983
rect 8039 915 8051 949
rect 8085 915 8097 949
rect 8039 881 8097 915
rect 8039 847 8051 881
rect 8085 847 8097 881
rect 8039 813 8097 847
rect 8039 779 8051 813
rect 8085 779 8097 813
rect 8039 745 8097 779
rect 8039 711 8051 745
rect 8085 711 8097 745
rect 8039 677 8097 711
rect 8039 643 8051 677
rect 8085 643 8097 677
rect 8039 609 8097 643
rect 8039 575 8051 609
rect 8085 575 8097 609
rect 8039 541 8097 575
rect 8039 507 8051 541
rect 8085 507 8097 541
rect 8039 473 8097 507
rect 8039 439 8051 473
rect 8085 439 8097 473
rect 8039 405 8097 439
rect 8039 371 8051 405
rect 8085 371 8097 405
rect 8039 355 8097 371
rect 8497 1629 8555 1645
rect 8497 1595 8509 1629
rect 8543 1595 8555 1629
rect 8497 1561 8555 1595
rect 8497 1527 8509 1561
rect 8543 1527 8555 1561
rect 8497 1493 8555 1527
rect 8497 1459 8509 1493
rect 8543 1459 8555 1493
rect 8497 1425 8555 1459
rect 8497 1391 8509 1425
rect 8543 1391 8555 1425
rect 8497 1357 8555 1391
rect 8497 1323 8509 1357
rect 8543 1323 8555 1357
rect 8497 1289 8555 1323
rect 8497 1255 8509 1289
rect 8543 1255 8555 1289
rect 8497 1221 8555 1255
rect 8497 1187 8509 1221
rect 8543 1187 8555 1221
rect 8497 1153 8555 1187
rect 8497 1119 8509 1153
rect 8543 1119 8555 1153
rect 8497 1085 8555 1119
rect 8497 1051 8509 1085
rect 8543 1051 8555 1085
rect 8497 1017 8555 1051
rect 8497 983 8509 1017
rect 8543 983 8555 1017
rect 8497 949 8555 983
rect 8497 915 8509 949
rect 8543 915 8555 949
rect 8497 881 8555 915
rect 8497 847 8509 881
rect 8543 847 8555 881
rect 8497 813 8555 847
rect 8497 779 8509 813
rect 8543 779 8555 813
rect 8497 745 8555 779
rect 8497 711 8509 745
rect 8543 711 8555 745
rect 8497 677 8555 711
rect 8497 643 8509 677
rect 8543 643 8555 677
rect 8497 609 8555 643
rect 8497 575 8509 609
rect 8543 575 8555 609
rect 8497 541 8555 575
rect 8497 507 8509 541
rect 8543 507 8555 541
rect 8497 473 8555 507
rect 8497 439 8509 473
rect 8543 439 8555 473
rect 8497 405 8555 439
rect 8497 371 8509 405
rect 8543 371 8555 405
rect 8497 355 8555 371
rect 8955 1629 9013 1645
rect 8955 1595 8967 1629
rect 9001 1595 9013 1629
rect 8955 1561 9013 1595
rect 8955 1527 8967 1561
rect 9001 1527 9013 1561
rect 8955 1493 9013 1527
rect 8955 1459 8967 1493
rect 9001 1459 9013 1493
rect 8955 1425 9013 1459
rect 8955 1391 8967 1425
rect 9001 1391 9013 1425
rect 8955 1357 9013 1391
rect 8955 1323 8967 1357
rect 9001 1323 9013 1357
rect 8955 1289 9013 1323
rect 8955 1255 8967 1289
rect 9001 1255 9013 1289
rect 8955 1221 9013 1255
rect 8955 1187 8967 1221
rect 9001 1187 9013 1221
rect 8955 1153 9013 1187
rect 8955 1119 8967 1153
rect 9001 1119 9013 1153
rect 8955 1085 9013 1119
rect 8955 1051 8967 1085
rect 9001 1051 9013 1085
rect 8955 1017 9013 1051
rect 8955 983 8967 1017
rect 9001 983 9013 1017
rect 8955 949 9013 983
rect 8955 915 8967 949
rect 9001 915 9013 949
rect 8955 881 9013 915
rect 8955 847 8967 881
rect 9001 847 9013 881
rect 8955 813 9013 847
rect 8955 779 8967 813
rect 9001 779 9013 813
rect 8955 745 9013 779
rect 8955 711 8967 745
rect 9001 711 9013 745
rect 8955 677 9013 711
rect 8955 643 8967 677
rect 9001 643 9013 677
rect 8955 609 9013 643
rect 8955 575 8967 609
rect 9001 575 9013 609
rect 8955 541 9013 575
rect 8955 507 8967 541
rect 9001 507 9013 541
rect 8955 473 9013 507
rect 8955 439 8967 473
rect 9001 439 9013 473
rect 8955 405 9013 439
rect 8955 371 8967 405
rect 9001 371 9013 405
rect 8955 355 9013 371
rect 9413 1629 9471 1645
rect 9413 1595 9425 1629
rect 9459 1595 9471 1629
rect 9413 1561 9471 1595
rect 9413 1527 9425 1561
rect 9459 1527 9471 1561
rect 9413 1493 9471 1527
rect 9413 1459 9425 1493
rect 9459 1459 9471 1493
rect 9413 1425 9471 1459
rect 9413 1391 9425 1425
rect 9459 1391 9471 1425
rect 9413 1357 9471 1391
rect 9413 1323 9425 1357
rect 9459 1323 9471 1357
rect 9413 1289 9471 1323
rect 9413 1255 9425 1289
rect 9459 1255 9471 1289
rect 9413 1221 9471 1255
rect 9413 1187 9425 1221
rect 9459 1187 9471 1221
rect 9413 1153 9471 1187
rect 9413 1119 9425 1153
rect 9459 1119 9471 1153
rect 9413 1085 9471 1119
rect 9413 1051 9425 1085
rect 9459 1051 9471 1085
rect 9413 1017 9471 1051
rect 9413 983 9425 1017
rect 9459 983 9471 1017
rect 9413 949 9471 983
rect 9413 915 9425 949
rect 9459 915 9471 949
rect 9413 881 9471 915
rect 9413 847 9425 881
rect 9459 847 9471 881
rect 9413 813 9471 847
rect 9413 779 9425 813
rect 9459 779 9471 813
rect 9413 745 9471 779
rect 9413 711 9425 745
rect 9459 711 9471 745
rect 9413 677 9471 711
rect 9413 643 9425 677
rect 9459 643 9471 677
rect 9413 609 9471 643
rect 9413 575 9425 609
rect 9459 575 9471 609
rect 9413 541 9471 575
rect 9413 507 9425 541
rect 9459 507 9471 541
rect 9413 473 9471 507
rect 9413 439 9425 473
rect 9459 439 9471 473
rect 9413 405 9471 439
rect 9413 371 9425 405
rect 9459 371 9471 405
rect 9413 355 9471 371
rect 9871 1629 9929 1645
rect 9871 1595 9883 1629
rect 9917 1595 9929 1629
rect 9871 1561 9929 1595
rect 9871 1527 9883 1561
rect 9917 1527 9929 1561
rect 9871 1493 9929 1527
rect 9871 1459 9883 1493
rect 9917 1459 9929 1493
rect 9871 1425 9929 1459
rect 9871 1391 9883 1425
rect 9917 1391 9929 1425
rect 9871 1357 9929 1391
rect 9871 1323 9883 1357
rect 9917 1323 9929 1357
rect 9871 1289 9929 1323
rect 9871 1255 9883 1289
rect 9917 1255 9929 1289
rect 9871 1221 9929 1255
rect 9871 1187 9883 1221
rect 9917 1187 9929 1221
rect 9871 1153 9929 1187
rect 9871 1119 9883 1153
rect 9917 1119 9929 1153
rect 9871 1085 9929 1119
rect 9871 1051 9883 1085
rect 9917 1051 9929 1085
rect 9871 1017 9929 1051
rect 9871 983 9883 1017
rect 9917 983 9929 1017
rect 9871 949 9929 983
rect 9871 915 9883 949
rect 9917 915 9929 949
rect 9871 881 9929 915
rect 9871 847 9883 881
rect 9917 847 9929 881
rect 9871 813 9929 847
rect 9871 779 9883 813
rect 9917 779 9929 813
rect 9871 745 9929 779
rect 9871 711 9883 745
rect 9917 711 9929 745
rect 9871 677 9929 711
rect 9871 643 9883 677
rect 9917 643 9929 677
rect 9871 609 9929 643
rect 9871 575 9883 609
rect 9917 575 9929 609
rect 9871 541 9929 575
rect 9871 507 9883 541
rect 9917 507 9929 541
rect 9871 473 9929 507
rect 9871 439 9883 473
rect 9917 439 9929 473
rect 9871 405 9929 439
rect 9871 371 9883 405
rect 9917 371 9929 405
rect 9871 355 9929 371
rect 10329 1629 10387 1645
rect 10329 1595 10341 1629
rect 10375 1595 10387 1629
rect 10329 1561 10387 1595
rect 10329 1527 10341 1561
rect 10375 1527 10387 1561
rect 10329 1493 10387 1527
rect 10329 1459 10341 1493
rect 10375 1459 10387 1493
rect 10329 1425 10387 1459
rect 10329 1391 10341 1425
rect 10375 1391 10387 1425
rect 10329 1357 10387 1391
rect 10329 1323 10341 1357
rect 10375 1323 10387 1357
rect 10329 1289 10387 1323
rect 10329 1255 10341 1289
rect 10375 1255 10387 1289
rect 10329 1221 10387 1255
rect 10329 1187 10341 1221
rect 10375 1187 10387 1221
rect 10329 1153 10387 1187
rect 10329 1119 10341 1153
rect 10375 1119 10387 1153
rect 10329 1085 10387 1119
rect 10329 1051 10341 1085
rect 10375 1051 10387 1085
rect 10329 1017 10387 1051
rect 10329 983 10341 1017
rect 10375 983 10387 1017
rect 10329 949 10387 983
rect 10329 915 10341 949
rect 10375 915 10387 949
rect 10329 881 10387 915
rect 10329 847 10341 881
rect 10375 847 10387 881
rect 10329 813 10387 847
rect 10329 779 10341 813
rect 10375 779 10387 813
rect 10329 745 10387 779
rect 10329 711 10341 745
rect 10375 711 10387 745
rect 10329 677 10387 711
rect 10329 643 10341 677
rect 10375 643 10387 677
rect 10329 609 10387 643
rect 10329 575 10341 609
rect 10375 575 10387 609
rect 10329 541 10387 575
rect 10329 507 10341 541
rect 10375 507 10387 541
rect 10329 473 10387 507
rect 10329 439 10341 473
rect 10375 439 10387 473
rect 10329 405 10387 439
rect 10329 371 10341 405
rect 10375 371 10387 405
rect 10329 355 10387 371
rect 10787 1629 10845 1645
rect 10787 1595 10799 1629
rect 10833 1595 10845 1629
rect 10787 1561 10845 1595
rect 10787 1527 10799 1561
rect 10833 1527 10845 1561
rect 10787 1493 10845 1527
rect 10787 1459 10799 1493
rect 10833 1459 10845 1493
rect 10787 1425 10845 1459
rect 10787 1391 10799 1425
rect 10833 1391 10845 1425
rect 10787 1357 10845 1391
rect 10787 1323 10799 1357
rect 10833 1323 10845 1357
rect 10787 1289 10845 1323
rect 10787 1255 10799 1289
rect 10833 1255 10845 1289
rect 10787 1221 10845 1255
rect 10787 1187 10799 1221
rect 10833 1187 10845 1221
rect 10787 1153 10845 1187
rect 10787 1119 10799 1153
rect 10833 1119 10845 1153
rect 10787 1085 10845 1119
rect 10787 1051 10799 1085
rect 10833 1051 10845 1085
rect 10787 1017 10845 1051
rect 10787 983 10799 1017
rect 10833 983 10845 1017
rect 10787 949 10845 983
rect 10787 915 10799 949
rect 10833 915 10845 949
rect 10787 881 10845 915
rect 10787 847 10799 881
rect 10833 847 10845 881
rect 10787 813 10845 847
rect 10787 779 10799 813
rect 10833 779 10845 813
rect 10787 745 10845 779
rect 10787 711 10799 745
rect 10833 711 10845 745
rect 10787 677 10845 711
rect 10787 643 10799 677
rect 10833 643 10845 677
rect 10787 609 10845 643
rect 10787 575 10799 609
rect 10833 575 10845 609
rect 10787 541 10845 575
rect 10787 507 10799 541
rect 10833 507 10845 541
rect 10787 473 10845 507
rect 10787 439 10799 473
rect 10833 439 10845 473
rect 10787 405 10845 439
rect 10787 371 10799 405
rect 10833 371 10845 405
rect 10787 355 10845 371
rect 11245 1629 11303 1645
rect 11245 1595 11257 1629
rect 11291 1595 11303 1629
rect 11245 1561 11303 1595
rect 11245 1527 11257 1561
rect 11291 1527 11303 1561
rect 11245 1493 11303 1527
rect 11245 1459 11257 1493
rect 11291 1459 11303 1493
rect 11245 1425 11303 1459
rect 11245 1391 11257 1425
rect 11291 1391 11303 1425
rect 11245 1357 11303 1391
rect 11245 1323 11257 1357
rect 11291 1323 11303 1357
rect 11245 1289 11303 1323
rect 11245 1255 11257 1289
rect 11291 1255 11303 1289
rect 11245 1221 11303 1255
rect 11245 1187 11257 1221
rect 11291 1187 11303 1221
rect 11245 1153 11303 1187
rect 11245 1119 11257 1153
rect 11291 1119 11303 1153
rect 11245 1085 11303 1119
rect 11245 1051 11257 1085
rect 11291 1051 11303 1085
rect 11245 1017 11303 1051
rect 11245 983 11257 1017
rect 11291 983 11303 1017
rect 11245 949 11303 983
rect 11245 915 11257 949
rect 11291 915 11303 949
rect 11245 881 11303 915
rect 11245 847 11257 881
rect 11291 847 11303 881
rect 11245 813 11303 847
rect 11245 779 11257 813
rect 11291 779 11303 813
rect 11245 745 11303 779
rect 11245 711 11257 745
rect 11291 711 11303 745
rect 11245 677 11303 711
rect 11245 643 11257 677
rect 11291 643 11303 677
rect 11245 609 11303 643
rect 11245 575 11257 609
rect 11291 575 11303 609
rect 11245 541 11303 575
rect 11245 507 11257 541
rect 11291 507 11303 541
rect 11245 473 11303 507
rect 11245 439 11257 473
rect 11291 439 11303 473
rect 11245 405 11303 439
rect 11245 371 11257 405
rect 11291 371 11303 405
rect 11245 355 11303 371
rect 11703 1629 11761 1645
rect 11703 1595 11715 1629
rect 11749 1595 11761 1629
rect 11703 1561 11761 1595
rect 11703 1527 11715 1561
rect 11749 1527 11761 1561
rect 11703 1493 11761 1527
rect 11703 1459 11715 1493
rect 11749 1459 11761 1493
rect 11703 1425 11761 1459
rect 11703 1391 11715 1425
rect 11749 1391 11761 1425
rect 11703 1357 11761 1391
rect 11703 1323 11715 1357
rect 11749 1323 11761 1357
rect 11703 1289 11761 1323
rect 11703 1255 11715 1289
rect 11749 1255 11761 1289
rect 11703 1221 11761 1255
rect 11703 1187 11715 1221
rect 11749 1187 11761 1221
rect 11703 1153 11761 1187
rect 11703 1119 11715 1153
rect 11749 1119 11761 1153
rect 11703 1085 11761 1119
rect 11703 1051 11715 1085
rect 11749 1051 11761 1085
rect 11703 1017 11761 1051
rect 11703 983 11715 1017
rect 11749 983 11761 1017
rect 11703 949 11761 983
rect 11703 915 11715 949
rect 11749 915 11761 949
rect 11703 881 11761 915
rect 11703 847 11715 881
rect 11749 847 11761 881
rect 11703 813 11761 847
rect 11703 779 11715 813
rect 11749 779 11761 813
rect 11703 745 11761 779
rect 11703 711 11715 745
rect 11749 711 11761 745
rect 11703 677 11761 711
rect 11703 643 11715 677
rect 11749 643 11761 677
rect 11703 609 11761 643
rect 11703 575 11715 609
rect 11749 575 11761 609
rect 11703 541 11761 575
rect 11703 507 11715 541
rect 11749 507 11761 541
rect 11703 473 11761 507
rect 11703 439 11715 473
rect 11749 439 11761 473
rect 11703 405 11761 439
rect 11703 371 11715 405
rect 11749 371 11761 405
rect 11703 355 11761 371
rect 12161 1629 12219 1645
rect 12161 1595 12173 1629
rect 12207 1595 12219 1629
rect 12161 1561 12219 1595
rect 12161 1527 12173 1561
rect 12207 1527 12219 1561
rect 12161 1493 12219 1527
rect 12161 1459 12173 1493
rect 12207 1459 12219 1493
rect 12161 1425 12219 1459
rect 12161 1391 12173 1425
rect 12207 1391 12219 1425
rect 12161 1357 12219 1391
rect 12161 1323 12173 1357
rect 12207 1323 12219 1357
rect 12161 1289 12219 1323
rect 12161 1255 12173 1289
rect 12207 1255 12219 1289
rect 12161 1221 12219 1255
rect 12161 1187 12173 1221
rect 12207 1187 12219 1221
rect 12161 1153 12219 1187
rect 12161 1119 12173 1153
rect 12207 1119 12219 1153
rect 12161 1085 12219 1119
rect 12161 1051 12173 1085
rect 12207 1051 12219 1085
rect 12161 1017 12219 1051
rect 12161 983 12173 1017
rect 12207 983 12219 1017
rect 12161 949 12219 983
rect 12161 915 12173 949
rect 12207 915 12219 949
rect 12161 881 12219 915
rect 12161 847 12173 881
rect 12207 847 12219 881
rect 12161 813 12219 847
rect 12161 779 12173 813
rect 12207 779 12219 813
rect 12161 745 12219 779
rect 12161 711 12173 745
rect 12207 711 12219 745
rect 12161 677 12219 711
rect 12161 643 12173 677
rect 12207 643 12219 677
rect 12161 609 12219 643
rect 12161 575 12173 609
rect 12207 575 12219 609
rect 12161 541 12219 575
rect 12161 507 12173 541
rect 12207 507 12219 541
rect 12161 473 12219 507
rect 12161 439 12173 473
rect 12207 439 12219 473
rect 12161 405 12219 439
rect 12161 371 12173 405
rect 12207 371 12219 405
rect 12161 355 12219 371
rect 12619 1629 12677 1645
rect 12619 1595 12631 1629
rect 12665 1595 12677 1629
rect 12619 1561 12677 1595
rect 12619 1527 12631 1561
rect 12665 1527 12677 1561
rect 12619 1493 12677 1527
rect 12619 1459 12631 1493
rect 12665 1459 12677 1493
rect 12619 1425 12677 1459
rect 12619 1391 12631 1425
rect 12665 1391 12677 1425
rect 12619 1357 12677 1391
rect 12619 1323 12631 1357
rect 12665 1323 12677 1357
rect 12619 1289 12677 1323
rect 12619 1255 12631 1289
rect 12665 1255 12677 1289
rect 12619 1221 12677 1255
rect 12619 1187 12631 1221
rect 12665 1187 12677 1221
rect 12619 1153 12677 1187
rect 12619 1119 12631 1153
rect 12665 1119 12677 1153
rect 12619 1085 12677 1119
rect 12619 1051 12631 1085
rect 12665 1051 12677 1085
rect 12619 1017 12677 1051
rect 12619 983 12631 1017
rect 12665 983 12677 1017
rect 12619 949 12677 983
rect 12619 915 12631 949
rect 12665 915 12677 949
rect 12619 881 12677 915
rect 12619 847 12631 881
rect 12665 847 12677 881
rect 12619 813 12677 847
rect 12619 779 12631 813
rect 12665 779 12677 813
rect 12619 745 12677 779
rect 12619 711 12631 745
rect 12665 711 12677 745
rect 12619 677 12677 711
rect 12619 643 12631 677
rect 12665 643 12677 677
rect 12619 609 12677 643
rect 12619 575 12631 609
rect 12665 575 12677 609
rect 12619 541 12677 575
rect 12619 507 12631 541
rect 12665 507 12677 541
rect 12619 473 12677 507
rect 12619 439 12631 473
rect 12665 439 12677 473
rect 12619 405 12677 439
rect 12619 371 12631 405
rect 12665 371 12677 405
rect 12619 355 12677 371
rect 13077 1629 13135 1645
rect 13077 1595 13089 1629
rect 13123 1595 13135 1629
rect 13077 1561 13135 1595
rect 13077 1527 13089 1561
rect 13123 1527 13135 1561
rect 13077 1493 13135 1527
rect 13077 1459 13089 1493
rect 13123 1459 13135 1493
rect 13077 1425 13135 1459
rect 13077 1391 13089 1425
rect 13123 1391 13135 1425
rect 13077 1357 13135 1391
rect 13077 1323 13089 1357
rect 13123 1323 13135 1357
rect 13077 1289 13135 1323
rect 13077 1255 13089 1289
rect 13123 1255 13135 1289
rect 13077 1221 13135 1255
rect 13077 1187 13089 1221
rect 13123 1187 13135 1221
rect 13077 1153 13135 1187
rect 13077 1119 13089 1153
rect 13123 1119 13135 1153
rect 13077 1085 13135 1119
rect 13077 1051 13089 1085
rect 13123 1051 13135 1085
rect 13077 1017 13135 1051
rect 13077 983 13089 1017
rect 13123 983 13135 1017
rect 13077 949 13135 983
rect 13077 915 13089 949
rect 13123 915 13135 949
rect 13077 881 13135 915
rect 13077 847 13089 881
rect 13123 847 13135 881
rect 13077 813 13135 847
rect 13077 779 13089 813
rect 13123 779 13135 813
rect 13077 745 13135 779
rect 13077 711 13089 745
rect 13123 711 13135 745
rect 13077 677 13135 711
rect 13077 643 13089 677
rect 13123 643 13135 677
rect 13077 609 13135 643
rect 13077 575 13089 609
rect 13123 575 13135 609
rect 13077 541 13135 575
rect 13077 507 13089 541
rect 13123 507 13135 541
rect 13077 473 13135 507
rect 13077 439 13089 473
rect 13123 439 13135 473
rect 13077 405 13135 439
rect 13077 371 13089 405
rect 13123 371 13135 405
rect 13077 355 13135 371
rect 13535 1629 13593 1645
rect 13535 1595 13547 1629
rect 13581 1595 13593 1629
rect 13535 1561 13593 1595
rect 13535 1527 13547 1561
rect 13581 1527 13593 1561
rect 13535 1493 13593 1527
rect 13535 1459 13547 1493
rect 13581 1459 13593 1493
rect 13535 1425 13593 1459
rect 13535 1391 13547 1425
rect 13581 1391 13593 1425
rect 13535 1357 13593 1391
rect 13535 1323 13547 1357
rect 13581 1323 13593 1357
rect 13535 1289 13593 1323
rect 13535 1255 13547 1289
rect 13581 1255 13593 1289
rect 13535 1221 13593 1255
rect 13535 1187 13547 1221
rect 13581 1187 13593 1221
rect 13535 1153 13593 1187
rect 13535 1119 13547 1153
rect 13581 1119 13593 1153
rect 13535 1085 13593 1119
rect 13535 1051 13547 1085
rect 13581 1051 13593 1085
rect 13535 1017 13593 1051
rect 13535 983 13547 1017
rect 13581 983 13593 1017
rect 13535 949 13593 983
rect 13535 915 13547 949
rect 13581 915 13593 949
rect 13535 881 13593 915
rect 13535 847 13547 881
rect 13581 847 13593 881
rect 13535 813 13593 847
rect 13535 779 13547 813
rect 13581 779 13593 813
rect 13535 745 13593 779
rect 13535 711 13547 745
rect 13581 711 13593 745
rect 13535 677 13593 711
rect 13535 643 13547 677
rect 13581 643 13593 677
rect 13535 609 13593 643
rect 13535 575 13547 609
rect 13581 575 13593 609
rect 13535 541 13593 575
rect 13535 507 13547 541
rect 13581 507 13593 541
rect 13535 473 13593 507
rect 13535 439 13547 473
rect 13581 439 13593 473
rect 13535 405 13593 439
rect 13535 371 13547 405
rect 13581 371 13593 405
rect 13535 355 13593 371
rect 13993 1629 14051 1645
rect 13993 1595 14005 1629
rect 14039 1595 14051 1629
rect 13993 1561 14051 1595
rect 13993 1527 14005 1561
rect 14039 1527 14051 1561
rect 13993 1493 14051 1527
rect 13993 1459 14005 1493
rect 14039 1459 14051 1493
rect 13993 1425 14051 1459
rect 13993 1391 14005 1425
rect 14039 1391 14051 1425
rect 13993 1357 14051 1391
rect 13993 1323 14005 1357
rect 14039 1323 14051 1357
rect 13993 1289 14051 1323
rect 13993 1255 14005 1289
rect 14039 1255 14051 1289
rect 13993 1221 14051 1255
rect 13993 1187 14005 1221
rect 14039 1187 14051 1221
rect 13993 1153 14051 1187
rect 13993 1119 14005 1153
rect 14039 1119 14051 1153
rect 13993 1085 14051 1119
rect 13993 1051 14005 1085
rect 14039 1051 14051 1085
rect 13993 1017 14051 1051
rect 13993 983 14005 1017
rect 14039 983 14051 1017
rect 13993 949 14051 983
rect 13993 915 14005 949
rect 14039 915 14051 949
rect 13993 881 14051 915
rect 13993 847 14005 881
rect 14039 847 14051 881
rect 13993 813 14051 847
rect 13993 779 14005 813
rect 14039 779 14051 813
rect 13993 745 14051 779
rect 13993 711 14005 745
rect 14039 711 14051 745
rect 13993 677 14051 711
rect 13993 643 14005 677
rect 14039 643 14051 677
rect 13993 609 14051 643
rect 13993 575 14005 609
rect 14039 575 14051 609
rect 13993 541 14051 575
rect 13993 507 14005 541
rect 14039 507 14051 541
rect 13993 473 14051 507
rect 13993 439 14005 473
rect 14039 439 14051 473
rect 13993 405 14051 439
rect 13993 371 14005 405
rect 14039 371 14051 405
rect 13993 355 14051 371
rect 14451 1629 14509 1645
rect 14451 1595 14463 1629
rect 14497 1595 14509 1629
rect 14451 1561 14509 1595
rect 14451 1527 14463 1561
rect 14497 1527 14509 1561
rect 14451 1493 14509 1527
rect 14451 1459 14463 1493
rect 14497 1459 14509 1493
rect 14451 1425 14509 1459
rect 14451 1391 14463 1425
rect 14497 1391 14509 1425
rect 14451 1357 14509 1391
rect 14451 1323 14463 1357
rect 14497 1323 14509 1357
rect 14451 1289 14509 1323
rect 14451 1255 14463 1289
rect 14497 1255 14509 1289
rect 14451 1221 14509 1255
rect 14451 1187 14463 1221
rect 14497 1187 14509 1221
rect 14451 1153 14509 1187
rect 14451 1119 14463 1153
rect 14497 1119 14509 1153
rect 14451 1085 14509 1119
rect 14451 1051 14463 1085
rect 14497 1051 14509 1085
rect 14451 1017 14509 1051
rect 14451 983 14463 1017
rect 14497 983 14509 1017
rect 14451 949 14509 983
rect 14451 915 14463 949
rect 14497 915 14509 949
rect 14451 881 14509 915
rect 14451 847 14463 881
rect 14497 847 14509 881
rect 14451 813 14509 847
rect 14451 779 14463 813
rect 14497 779 14509 813
rect 14451 745 14509 779
rect 14451 711 14463 745
rect 14497 711 14509 745
rect 14451 677 14509 711
rect 14451 643 14463 677
rect 14497 643 14509 677
rect 14451 609 14509 643
rect 14451 575 14463 609
rect 14497 575 14509 609
rect 14451 541 14509 575
rect 14451 507 14463 541
rect 14497 507 14509 541
rect 14451 473 14509 507
rect 14451 439 14463 473
rect 14497 439 14509 473
rect 14451 405 14509 439
rect 14451 371 14463 405
rect 14497 371 14509 405
rect 14451 355 14509 371
rect 14909 1629 14967 1645
rect 14909 1595 14921 1629
rect 14955 1595 14967 1629
rect 14909 1561 14967 1595
rect 14909 1527 14921 1561
rect 14955 1527 14967 1561
rect 14909 1493 14967 1527
rect 14909 1459 14921 1493
rect 14955 1459 14967 1493
rect 14909 1425 14967 1459
rect 14909 1391 14921 1425
rect 14955 1391 14967 1425
rect 14909 1357 14967 1391
rect 14909 1323 14921 1357
rect 14955 1323 14967 1357
rect 14909 1289 14967 1323
rect 14909 1255 14921 1289
rect 14955 1255 14967 1289
rect 14909 1221 14967 1255
rect 14909 1187 14921 1221
rect 14955 1187 14967 1221
rect 14909 1153 14967 1187
rect 14909 1119 14921 1153
rect 14955 1119 14967 1153
rect 14909 1085 14967 1119
rect 14909 1051 14921 1085
rect 14955 1051 14967 1085
rect 14909 1017 14967 1051
rect 14909 983 14921 1017
rect 14955 983 14967 1017
rect 14909 949 14967 983
rect 14909 915 14921 949
rect 14955 915 14967 949
rect 14909 881 14967 915
rect 14909 847 14921 881
rect 14955 847 14967 881
rect 14909 813 14967 847
rect 14909 779 14921 813
rect 14955 779 14967 813
rect 14909 745 14967 779
rect 14909 711 14921 745
rect 14955 711 14967 745
rect 14909 677 14967 711
rect 14909 643 14921 677
rect 14955 643 14967 677
rect 14909 609 14967 643
rect 14909 575 14921 609
rect 14955 575 14967 609
rect 14909 541 14967 575
rect 14909 507 14921 541
rect 14955 507 14967 541
rect 14909 473 14967 507
rect 14909 439 14921 473
rect 14955 439 14967 473
rect 14909 405 14967 439
rect 14909 371 14921 405
rect 14955 371 14967 405
rect 14909 355 14967 371
rect 15367 1629 15425 1645
rect 15367 1595 15379 1629
rect 15413 1595 15425 1629
rect 15367 1561 15425 1595
rect 15367 1527 15379 1561
rect 15413 1527 15425 1561
rect 15367 1493 15425 1527
rect 15367 1459 15379 1493
rect 15413 1459 15425 1493
rect 15367 1425 15425 1459
rect 15367 1391 15379 1425
rect 15413 1391 15425 1425
rect 15367 1357 15425 1391
rect 15367 1323 15379 1357
rect 15413 1323 15425 1357
rect 15367 1289 15425 1323
rect 15367 1255 15379 1289
rect 15413 1255 15425 1289
rect 15367 1221 15425 1255
rect 15367 1187 15379 1221
rect 15413 1187 15425 1221
rect 15367 1153 15425 1187
rect 15367 1119 15379 1153
rect 15413 1119 15425 1153
rect 15367 1085 15425 1119
rect 15367 1051 15379 1085
rect 15413 1051 15425 1085
rect 15367 1017 15425 1051
rect 15367 983 15379 1017
rect 15413 983 15425 1017
rect 15367 949 15425 983
rect 15367 915 15379 949
rect 15413 915 15425 949
rect 15367 881 15425 915
rect 15367 847 15379 881
rect 15413 847 15425 881
rect 15367 813 15425 847
rect 15367 779 15379 813
rect 15413 779 15425 813
rect 15367 745 15425 779
rect 15367 711 15379 745
rect 15413 711 15425 745
rect 15367 677 15425 711
rect 15367 643 15379 677
rect 15413 643 15425 677
rect 15367 609 15425 643
rect 15367 575 15379 609
rect 15413 575 15425 609
rect 15367 541 15425 575
rect 15367 507 15379 541
rect 15413 507 15425 541
rect 15367 473 15425 507
rect 15367 439 15379 473
rect 15413 439 15425 473
rect 15367 405 15425 439
rect 15367 371 15379 405
rect 15413 371 15425 405
rect 15367 355 15425 371
rect 15825 1629 15883 1645
rect 15825 1595 15837 1629
rect 15871 1595 15883 1629
rect 15825 1561 15883 1595
rect 15825 1527 15837 1561
rect 15871 1527 15883 1561
rect 15825 1493 15883 1527
rect 15825 1459 15837 1493
rect 15871 1459 15883 1493
rect 15825 1425 15883 1459
rect 15825 1391 15837 1425
rect 15871 1391 15883 1425
rect 15825 1357 15883 1391
rect 15825 1323 15837 1357
rect 15871 1323 15883 1357
rect 15825 1289 15883 1323
rect 15825 1255 15837 1289
rect 15871 1255 15883 1289
rect 15825 1221 15883 1255
rect 15825 1187 15837 1221
rect 15871 1187 15883 1221
rect 15825 1153 15883 1187
rect 15825 1119 15837 1153
rect 15871 1119 15883 1153
rect 15825 1085 15883 1119
rect 15825 1051 15837 1085
rect 15871 1051 15883 1085
rect 15825 1017 15883 1051
rect 15825 983 15837 1017
rect 15871 983 15883 1017
rect 15825 949 15883 983
rect 15825 915 15837 949
rect 15871 915 15883 949
rect 15825 881 15883 915
rect 15825 847 15837 881
rect 15871 847 15883 881
rect 15825 813 15883 847
rect 15825 779 15837 813
rect 15871 779 15883 813
rect 15825 745 15883 779
rect 15825 711 15837 745
rect 15871 711 15883 745
rect 15825 677 15883 711
rect 15825 643 15837 677
rect 15871 643 15883 677
rect 15825 609 15883 643
rect 15825 575 15837 609
rect 15871 575 15883 609
rect 15825 541 15883 575
rect 15825 507 15837 541
rect 15871 507 15883 541
rect 15825 473 15883 507
rect 15825 439 15837 473
rect 15871 439 15883 473
rect 15825 405 15883 439
rect 15825 371 15837 405
rect 15871 371 15883 405
rect 15825 355 15883 371
rect 16283 1629 16341 1645
rect 16283 1595 16295 1629
rect 16329 1595 16341 1629
rect 16283 1561 16341 1595
rect 16283 1527 16295 1561
rect 16329 1527 16341 1561
rect 16283 1493 16341 1527
rect 16283 1459 16295 1493
rect 16329 1459 16341 1493
rect 16283 1425 16341 1459
rect 16283 1391 16295 1425
rect 16329 1391 16341 1425
rect 16283 1357 16341 1391
rect 16283 1323 16295 1357
rect 16329 1323 16341 1357
rect 16283 1289 16341 1323
rect 16283 1255 16295 1289
rect 16329 1255 16341 1289
rect 16283 1221 16341 1255
rect 16283 1187 16295 1221
rect 16329 1187 16341 1221
rect 16283 1153 16341 1187
rect 16283 1119 16295 1153
rect 16329 1119 16341 1153
rect 16283 1085 16341 1119
rect 16283 1051 16295 1085
rect 16329 1051 16341 1085
rect 16283 1017 16341 1051
rect 16283 983 16295 1017
rect 16329 983 16341 1017
rect 16283 949 16341 983
rect 16283 915 16295 949
rect 16329 915 16341 949
rect 16283 881 16341 915
rect 16283 847 16295 881
rect 16329 847 16341 881
rect 16283 813 16341 847
rect 16283 779 16295 813
rect 16329 779 16341 813
rect 16283 745 16341 779
rect 16283 711 16295 745
rect 16329 711 16341 745
rect 16283 677 16341 711
rect 16283 643 16295 677
rect 16329 643 16341 677
rect 16283 609 16341 643
rect 16283 575 16295 609
rect 16329 575 16341 609
rect 16283 541 16341 575
rect 16283 507 16295 541
rect 16329 507 16341 541
rect 16283 473 16341 507
rect 16283 439 16295 473
rect 16329 439 16341 473
rect 16283 405 16341 439
rect 16283 371 16295 405
rect 16329 371 16341 405
rect 16283 355 16341 371
rect 16741 1629 16799 1645
rect 16741 1595 16753 1629
rect 16787 1595 16799 1629
rect 16741 1561 16799 1595
rect 16741 1527 16753 1561
rect 16787 1527 16799 1561
rect 16741 1493 16799 1527
rect 16741 1459 16753 1493
rect 16787 1459 16799 1493
rect 16741 1425 16799 1459
rect 16741 1391 16753 1425
rect 16787 1391 16799 1425
rect 16741 1357 16799 1391
rect 16741 1323 16753 1357
rect 16787 1323 16799 1357
rect 16741 1289 16799 1323
rect 16741 1255 16753 1289
rect 16787 1255 16799 1289
rect 16741 1221 16799 1255
rect 16741 1187 16753 1221
rect 16787 1187 16799 1221
rect 16741 1153 16799 1187
rect 16741 1119 16753 1153
rect 16787 1119 16799 1153
rect 16741 1085 16799 1119
rect 16741 1051 16753 1085
rect 16787 1051 16799 1085
rect 16741 1017 16799 1051
rect 16741 983 16753 1017
rect 16787 983 16799 1017
rect 16741 949 16799 983
rect 16741 915 16753 949
rect 16787 915 16799 949
rect 16741 881 16799 915
rect 16741 847 16753 881
rect 16787 847 16799 881
rect 16741 813 16799 847
rect 16741 779 16753 813
rect 16787 779 16799 813
rect 16741 745 16799 779
rect 16741 711 16753 745
rect 16787 711 16799 745
rect 16741 677 16799 711
rect 16741 643 16753 677
rect 16787 643 16799 677
rect 16741 609 16799 643
rect 16741 575 16753 609
rect 16787 575 16799 609
rect 16741 541 16799 575
rect 16741 507 16753 541
rect 16787 507 16799 541
rect 16741 473 16799 507
rect 16741 439 16753 473
rect 16787 439 16799 473
rect 16741 405 16799 439
rect 16741 371 16753 405
rect 16787 371 16799 405
rect 16741 355 16799 371
rect 17199 1629 17257 1645
rect 17199 1595 17211 1629
rect 17245 1595 17257 1629
rect 17199 1561 17257 1595
rect 17199 1527 17211 1561
rect 17245 1527 17257 1561
rect 17199 1493 17257 1527
rect 17199 1459 17211 1493
rect 17245 1459 17257 1493
rect 17199 1425 17257 1459
rect 17199 1391 17211 1425
rect 17245 1391 17257 1425
rect 17199 1357 17257 1391
rect 17199 1323 17211 1357
rect 17245 1323 17257 1357
rect 17199 1289 17257 1323
rect 17199 1255 17211 1289
rect 17245 1255 17257 1289
rect 17199 1221 17257 1255
rect 17199 1187 17211 1221
rect 17245 1187 17257 1221
rect 17199 1153 17257 1187
rect 17199 1119 17211 1153
rect 17245 1119 17257 1153
rect 17199 1085 17257 1119
rect 17199 1051 17211 1085
rect 17245 1051 17257 1085
rect 17199 1017 17257 1051
rect 17199 983 17211 1017
rect 17245 983 17257 1017
rect 17199 949 17257 983
rect 17199 915 17211 949
rect 17245 915 17257 949
rect 17199 881 17257 915
rect 17199 847 17211 881
rect 17245 847 17257 881
rect 17199 813 17257 847
rect 17199 779 17211 813
rect 17245 779 17257 813
rect 17199 745 17257 779
rect 17199 711 17211 745
rect 17245 711 17257 745
rect 17199 677 17257 711
rect 17199 643 17211 677
rect 17245 643 17257 677
rect 17199 609 17257 643
rect 17199 575 17211 609
rect 17245 575 17257 609
rect 17199 541 17257 575
rect 17199 507 17211 541
rect 17245 507 17257 541
rect 17199 473 17257 507
rect 17199 439 17211 473
rect 17245 439 17257 473
rect 17199 405 17257 439
rect 17199 371 17211 405
rect 17245 371 17257 405
rect 17199 355 17257 371
rect 17657 1629 17715 1645
rect 17657 1595 17669 1629
rect 17703 1595 17715 1629
rect 17657 1561 17715 1595
rect 17657 1527 17669 1561
rect 17703 1527 17715 1561
rect 17657 1493 17715 1527
rect 17657 1459 17669 1493
rect 17703 1459 17715 1493
rect 17657 1425 17715 1459
rect 17657 1391 17669 1425
rect 17703 1391 17715 1425
rect 17657 1357 17715 1391
rect 17657 1323 17669 1357
rect 17703 1323 17715 1357
rect 17657 1289 17715 1323
rect 17657 1255 17669 1289
rect 17703 1255 17715 1289
rect 17657 1221 17715 1255
rect 17657 1187 17669 1221
rect 17703 1187 17715 1221
rect 17657 1153 17715 1187
rect 17657 1119 17669 1153
rect 17703 1119 17715 1153
rect 17657 1085 17715 1119
rect 17657 1051 17669 1085
rect 17703 1051 17715 1085
rect 17657 1017 17715 1051
rect 17657 983 17669 1017
rect 17703 983 17715 1017
rect 17657 949 17715 983
rect 17657 915 17669 949
rect 17703 915 17715 949
rect 17657 881 17715 915
rect 17657 847 17669 881
rect 17703 847 17715 881
rect 17657 813 17715 847
rect 17657 779 17669 813
rect 17703 779 17715 813
rect 17657 745 17715 779
rect 17657 711 17669 745
rect 17703 711 17715 745
rect 17657 677 17715 711
rect 17657 643 17669 677
rect 17703 643 17715 677
rect 17657 609 17715 643
rect 17657 575 17669 609
rect 17703 575 17715 609
rect 17657 541 17715 575
rect 17657 507 17669 541
rect 17703 507 17715 541
rect 17657 473 17715 507
rect 17657 439 17669 473
rect 17703 439 17715 473
rect 17657 405 17715 439
rect 17657 371 17669 405
rect 17703 371 17715 405
rect 17657 355 17715 371
rect 18115 1629 18173 1645
rect 18115 1595 18127 1629
rect 18161 1595 18173 1629
rect 18115 1561 18173 1595
rect 18115 1527 18127 1561
rect 18161 1527 18173 1561
rect 18115 1493 18173 1527
rect 18115 1459 18127 1493
rect 18161 1459 18173 1493
rect 18115 1425 18173 1459
rect 18115 1391 18127 1425
rect 18161 1391 18173 1425
rect 18115 1357 18173 1391
rect 18115 1323 18127 1357
rect 18161 1323 18173 1357
rect 18115 1289 18173 1323
rect 18115 1255 18127 1289
rect 18161 1255 18173 1289
rect 18115 1221 18173 1255
rect 18115 1187 18127 1221
rect 18161 1187 18173 1221
rect 18115 1153 18173 1187
rect 18115 1119 18127 1153
rect 18161 1119 18173 1153
rect 18115 1085 18173 1119
rect 18115 1051 18127 1085
rect 18161 1051 18173 1085
rect 18115 1017 18173 1051
rect 18115 983 18127 1017
rect 18161 983 18173 1017
rect 18115 949 18173 983
rect 18115 915 18127 949
rect 18161 915 18173 949
rect 18115 881 18173 915
rect 18115 847 18127 881
rect 18161 847 18173 881
rect 18115 813 18173 847
rect 18115 779 18127 813
rect 18161 779 18173 813
rect 18115 745 18173 779
rect 18115 711 18127 745
rect 18161 711 18173 745
rect 18115 677 18173 711
rect 18115 643 18127 677
rect 18161 643 18173 677
rect 18115 609 18173 643
rect 18115 575 18127 609
rect 18161 575 18173 609
rect 18115 541 18173 575
rect 18115 507 18127 541
rect 18161 507 18173 541
rect 18115 473 18173 507
rect 18115 439 18127 473
rect 18161 439 18173 473
rect 18115 405 18173 439
rect 18115 371 18127 405
rect 18161 371 18173 405
rect 18115 355 18173 371
rect 18573 1629 18631 1645
rect 18573 1595 18585 1629
rect 18619 1595 18631 1629
rect 18573 1561 18631 1595
rect 18573 1527 18585 1561
rect 18619 1527 18631 1561
rect 18573 1493 18631 1527
rect 18573 1459 18585 1493
rect 18619 1459 18631 1493
rect 18573 1425 18631 1459
rect 18573 1391 18585 1425
rect 18619 1391 18631 1425
rect 18573 1357 18631 1391
rect 18573 1323 18585 1357
rect 18619 1323 18631 1357
rect 18573 1289 18631 1323
rect 18573 1255 18585 1289
rect 18619 1255 18631 1289
rect 18573 1221 18631 1255
rect 18573 1187 18585 1221
rect 18619 1187 18631 1221
rect 18573 1153 18631 1187
rect 18573 1119 18585 1153
rect 18619 1119 18631 1153
rect 18573 1085 18631 1119
rect 18573 1051 18585 1085
rect 18619 1051 18631 1085
rect 18573 1017 18631 1051
rect 18573 983 18585 1017
rect 18619 983 18631 1017
rect 18573 949 18631 983
rect 18573 915 18585 949
rect 18619 915 18631 949
rect 18573 881 18631 915
rect 18573 847 18585 881
rect 18619 847 18631 881
rect 18573 813 18631 847
rect 18573 779 18585 813
rect 18619 779 18631 813
rect 18573 745 18631 779
rect 18573 711 18585 745
rect 18619 711 18631 745
rect 18573 677 18631 711
rect 18573 643 18585 677
rect 18619 643 18631 677
rect 18573 609 18631 643
rect 18573 575 18585 609
rect 18619 575 18631 609
rect 18573 541 18631 575
rect 18573 507 18585 541
rect 18619 507 18631 541
rect 18573 473 18631 507
rect 18573 439 18585 473
rect 18619 439 18631 473
rect 18573 405 18631 439
rect 18573 371 18585 405
rect 18619 371 18631 405
rect 18573 355 18631 371
rect 19031 1629 19089 1645
rect 19031 1595 19043 1629
rect 19077 1595 19089 1629
rect 19031 1561 19089 1595
rect 19031 1527 19043 1561
rect 19077 1527 19089 1561
rect 19031 1493 19089 1527
rect 19031 1459 19043 1493
rect 19077 1459 19089 1493
rect 19031 1425 19089 1459
rect 19031 1391 19043 1425
rect 19077 1391 19089 1425
rect 19031 1357 19089 1391
rect 19031 1323 19043 1357
rect 19077 1323 19089 1357
rect 19031 1289 19089 1323
rect 19031 1255 19043 1289
rect 19077 1255 19089 1289
rect 19031 1221 19089 1255
rect 19031 1187 19043 1221
rect 19077 1187 19089 1221
rect 19031 1153 19089 1187
rect 19031 1119 19043 1153
rect 19077 1119 19089 1153
rect 19031 1085 19089 1119
rect 19031 1051 19043 1085
rect 19077 1051 19089 1085
rect 19031 1017 19089 1051
rect 19031 983 19043 1017
rect 19077 983 19089 1017
rect 19031 949 19089 983
rect 19031 915 19043 949
rect 19077 915 19089 949
rect 19031 881 19089 915
rect 19031 847 19043 881
rect 19077 847 19089 881
rect 19031 813 19089 847
rect 19031 779 19043 813
rect 19077 779 19089 813
rect 19031 745 19089 779
rect 19031 711 19043 745
rect 19077 711 19089 745
rect 19031 677 19089 711
rect 19031 643 19043 677
rect 19077 643 19089 677
rect 19031 609 19089 643
rect 19031 575 19043 609
rect 19077 575 19089 609
rect 19031 541 19089 575
rect 19031 507 19043 541
rect 19077 507 19089 541
rect 19031 473 19089 507
rect 19031 439 19043 473
rect 19077 439 19089 473
rect 19031 405 19089 439
rect 19031 371 19043 405
rect 19077 371 19089 405
rect 19031 355 19089 371
rect 19489 1629 19547 1645
rect 19489 1595 19501 1629
rect 19535 1595 19547 1629
rect 19489 1561 19547 1595
rect 19489 1527 19501 1561
rect 19535 1527 19547 1561
rect 19489 1493 19547 1527
rect 19489 1459 19501 1493
rect 19535 1459 19547 1493
rect 19489 1425 19547 1459
rect 19489 1391 19501 1425
rect 19535 1391 19547 1425
rect 19489 1357 19547 1391
rect 19489 1323 19501 1357
rect 19535 1323 19547 1357
rect 19489 1289 19547 1323
rect 19489 1255 19501 1289
rect 19535 1255 19547 1289
rect 19489 1221 19547 1255
rect 19489 1187 19501 1221
rect 19535 1187 19547 1221
rect 19489 1153 19547 1187
rect 19489 1119 19501 1153
rect 19535 1119 19547 1153
rect 19489 1085 19547 1119
rect 19489 1051 19501 1085
rect 19535 1051 19547 1085
rect 19489 1017 19547 1051
rect 19489 983 19501 1017
rect 19535 983 19547 1017
rect 19489 949 19547 983
rect 19489 915 19501 949
rect 19535 915 19547 949
rect 19489 881 19547 915
rect 19489 847 19501 881
rect 19535 847 19547 881
rect 19489 813 19547 847
rect 19489 779 19501 813
rect 19535 779 19547 813
rect 19489 745 19547 779
rect 19489 711 19501 745
rect 19535 711 19547 745
rect 19489 677 19547 711
rect 19489 643 19501 677
rect 19535 643 19547 677
rect 19489 609 19547 643
rect 19489 575 19501 609
rect 19535 575 19547 609
rect 19489 541 19547 575
rect 19489 507 19501 541
rect 19535 507 19547 541
rect 19489 473 19547 507
rect 19489 439 19501 473
rect 19535 439 19547 473
rect 19489 405 19547 439
rect 19489 371 19501 405
rect 19535 371 19547 405
rect 19489 355 19547 371
rect 19947 1629 20005 1645
rect 19947 1595 19959 1629
rect 19993 1595 20005 1629
rect 19947 1561 20005 1595
rect 19947 1527 19959 1561
rect 19993 1527 20005 1561
rect 19947 1493 20005 1527
rect 19947 1459 19959 1493
rect 19993 1459 20005 1493
rect 19947 1425 20005 1459
rect 19947 1391 19959 1425
rect 19993 1391 20005 1425
rect 19947 1357 20005 1391
rect 19947 1323 19959 1357
rect 19993 1323 20005 1357
rect 19947 1289 20005 1323
rect 19947 1255 19959 1289
rect 19993 1255 20005 1289
rect 19947 1221 20005 1255
rect 19947 1187 19959 1221
rect 19993 1187 20005 1221
rect 19947 1153 20005 1187
rect 19947 1119 19959 1153
rect 19993 1119 20005 1153
rect 19947 1085 20005 1119
rect 19947 1051 19959 1085
rect 19993 1051 20005 1085
rect 19947 1017 20005 1051
rect 19947 983 19959 1017
rect 19993 983 20005 1017
rect 19947 949 20005 983
rect 19947 915 19959 949
rect 19993 915 20005 949
rect 19947 881 20005 915
rect 19947 847 19959 881
rect 19993 847 20005 881
rect 19947 813 20005 847
rect 19947 779 19959 813
rect 19993 779 20005 813
rect 19947 745 20005 779
rect 19947 711 19959 745
rect 19993 711 20005 745
rect 19947 677 20005 711
rect 19947 643 19959 677
rect 19993 643 20005 677
rect 19947 609 20005 643
rect 19947 575 19959 609
rect 19993 575 20005 609
rect 19947 541 20005 575
rect 19947 507 19959 541
rect 19993 507 20005 541
rect 19947 473 20005 507
rect 19947 439 19959 473
rect 19993 439 20005 473
rect 19947 405 20005 439
rect 19947 371 19959 405
rect 19993 371 20005 405
rect 19947 355 20005 371
rect 20405 1629 20463 1645
rect 20405 1595 20417 1629
rect 20451 1595 20463 1629
rect 20405 1561 20463 1595
rect 20405 1527 20417 1561
rect 20451 1527 20463 1561
rect 20405 1493 20463 1527
rect 20405 1459 20417 1493
rect 20451 1459 20463 1493
rect 20405 1425 20463 1459
rect 20405 1391 20417 1425
rect 20451 1391 20463 1425
rect 20405 1357 20463 1391
rect 20405 1323 20417 1357
rect 20451 1323 20463 1357
rect 20405 1289 20463 1323
rect 20405 1255 20417 1289
rect 20451 1255 20463 1289
rect 20405 1221 20463 1255
rect 20405 1187 20417 1221
rect 20451 1187 20463 1221
rect 20405 1153 20463 1187
rect 20405 1119 20417 1153
rect 20451 1119 20463 1153
rect 20405 1085 20463 1119
rect 20405 1051 20417 1085
rect 20451 1051 20463 1085
rect 20405 1017 20463 1051
rect 20405 983 20417 1017
rect 20451 983 20463 1017
rect 20405 949 20463 983
rect 20405 915 20417 949
rect 20451 915 20463 949
rect 20405 881 20463 915
rect 20405 847 20417 881
rect 20451 847 20463 881
rect 20405 813 20463 847
rect 20405 779 20417 813
rect 20451 779 20463 813
rect 20405 745 20463 779
rect 20405 711 20417 745
rect 20451 711 20463 745
rect 20405 677 20463 711
rect 20405 643 20417 677
rect 20451 643 20463 677
rect 20405 609 20463 643
rect 20405 575 20417 609
rect 20451 575 20463 609
rect 20405 541 20463 575
rect 20405 507 20417 541
rect 20451 507 20463 541
rect 20405 473 20463 507
rect 20405 439 20417 473
rect 20451 439 20463 473
rect 20405 405 20463 439
rect 20405 371 20417 405
rect 20451 371 20463 405
rect 20405 355 20463 371
rect 20863 1629 20921 1645
rect 20863 1595 20875 1629
rect 20909 1595 20921 1629
rect 20863 1561 20921 1595
rect 20863 1527 20875 1561
rect 20909 1527 20921 1561
rect 20863 1493 20921 1527
rect 20863 1459 20875 1493
rect 20909 1459 20921 1493
rect 20863 1425 20921 1459
rect 20863 1391 20875 1425
rect 20909 1391 20921 1425
rect 20863 1357 20921 1391
rect 20863 1323 20875 1357
rect 20909 1323 20921 1357
rect 20863 1289 20921 1323
rect 20863 1255 20875 1289
rect 20909 1255 20921 1289
rect 20863 1221 20921 1255
rect 20863 1187 20875 1221
rect 20909 1187 20921 1221
rect 20863 1153 20921 1187
rect 20863 1119 20875 1153
rect 20909 1119 20921 1153
rect 20863 1085 20921 1119
rect 20863 1051 20875 1085
rect 20909 1051 20921 1085
rect 20863 1017 20921 1051
rect 20863 983 20875 1017
rect 20909 983 20921 1017
rect 20863 949 20921 983
rect 20863 915 20875 949
rect 20909 915 20921 949
rect 20863 881 20921 915
rect 20863 847 20875 881
rect 20909 847 20921 881
rect 20863 813 20921 847
rect 20863 779 20875 813
rect 20909 779 20921 813
rect 20863 745 20921 779
rect 20863 711 20875 745
rect 20909 711 20921 745
rect 20863 677 20921 711
rect 20863 643 20875 677
rect 20909 643 20921 677
rect 20863 609 20921 643
rect 20863 575 20875 609
rect 20909 575 20921 609
rect 20863 541 20921 575
rect 20863 507 20875 541
rect 20909 507 20921 541
rect 20863 473 20921 507
rect 20863 439 20875 473
rect 20909 439 20921 473
rect 20863 405 20921 439
rect 20863 371 20875 405
rect 20909 371 20921 405
rect 20863 355 20921 371
rect 21321 1629 21379 1645
rect 21321 1595 21333 1629
rect 21367 1595 21379 1629
rect 21321 1561 21379 1595
rect 21321 1527 21333 1561
rect 21367 1527 21379 1561
rect 21321 1493 21379 1527
rect 21321 1459 21333 1493
rect 21367 1459 21379 1493
rect 21321 1425 21379 1459
rect 21321 1391 21333 1425
rect 21367 1391 21379 1425
rect 21321 1357 21379 1391
rect 21321 1323 21333 1357
rect 21367 1323 21379 1357
rect 21321 1289 21379 1323
rect 21321 1255 21333 1289
rect 21367 1255 21379 1289
rect 21321 1221 21379 1255
rect 21321 1187 21333 1221
rect 21367 1187 21379 1221
rect 21321 1153 21379 1187
rect 21321 1119 21333 1153
rect 21367 1119 21379 1153
rect 21321 1085 21379 1119
rect 21321 1051 21333 1085
rect 21367 1051 21379 1085
rect 21321 1017 21379 1051
rect 21321 983 21333 1017
rect 21367 983 21379 1017
rect 21321 949 21379 983
rect 21321 915 21333 949
rect 21367 915 21379 949
rect 21321 881 21379 915
rect 21321 847 21333 881
rect 21367 847 21379 881
rect 21321 813 21379 847
rect 21321 779 21333 813
rect 21367 779 21379 813
rect 21321 745 21379 779
rect 21321 711 21333 745
rect 21367 711 21379 745
rect 21321 677 21379 711
rect 21321 643 21333 677
rect 21367 643 21379 677
rect 21321 609 21379 643
rect 21321 575 21333 609
rect 21367 575 21379 609
rect 21321 541 21379 575
rect 21321 507 21333 541
rect 21367 507 21379 541
rect 21321 473 21379 507
rect 21321 439 21333 473
rect 21367 439 21379 473
rect 21321 405 21379 439
rect 21321 371 21333 405
rect 21367 371 21379 405
rect 21321 355 21379 371
rect 21779 1629 21837 1645
rect 21779 1595 21791 1629
rect 21825 1595 21837 1629
rect 21779 1561 21837 1595
rect 21779 1527 21791 1561
rect 21825 1527 21837 1561
rect 21779 1493 21837 1527
rect 21779 1459 21791 1493
rect 21825 1459 21837 1493
rect 21779 1425 21837 1459
rect 21779 1391 21791 1425
rect 21825 1391 21837 1425
rect 21779 1357 21837 1391
rect 21779 1323 21791 1357
rect 21825 1323 21837 1357
rect 21779 1289 21837 1323
rect 21779 1255 21791 1289
rect 21825 1255 21837 1289
rect 21779 1221 21837 1255
rect 21779 1187 21791 1221
rect 21825 1187 21837 1221
rect 21779 1153 21837 1187
rect 21779 1119 21791 1153
rect 21825 1119 21837 1153
rect 21779 1085 21837 1119
rect 21779 1051 21791 1085
rect 21825 1051 21837 1085
rect 21779 1017 21837 1051
rect 21779 983 21791 1017
rect 21825 983 21837 1017
rect 21779 949 21837 983
rect 21779 915 21791 949
rect 21825 915 21837 949
rect 21779 881 21837 915
rect 21779 847 21791 881
rect 21825 847 21837 881
rect 21779 813 21837 847
rect 21779 779 21791 813
rect 21825 779 21837 813
rect 21779 745 21837 779
rect 21779 711 21791 745
rect 21825 711 21837 745
rect 21779 677 21837 711
rect 21779 643 21791 677
rect 21825 643 21837 677
rect 21779 609 21837 643
rect 21779 575 21791 609
rect 21825 575 21837 609
rect 21779 541 21837 575
rect 21779 507 21791 541
rect 21825 507 21837 541
rect 21779 473 21837 507
rect 21779 439 21791 473
rect 21825 439 21837 473
rect 21779 405 21837 439
rect 21779 371 21791 405
rect 21825 371 21837 405
rect 21779 355 21837 371
rect 22237 1629 22295 1645
rect 22237 1595 22249 1629
rect 22283 1595 22295 1629
rect 22237 1561 22295 1595
rect 22237 1527 22249 1561
rect 22283 1527 22295 1561
rect 22237 1493 22295 1527
rect 22237 1459 22249 1493
rect 22283 1459 22295 1493
rect 22237 1425 22295 1459
rect 22237 1391 22249 1425
rect 22283 1391 22295 1425
rect 22237 1357 22295 1391
rect 22237 1323 22249 1357
rect 22283 1323 22295 1357
rect 22237 1289 22295 1323
rect 22237 1255 22249 1289
rect 22283 1255 22295 1289
rect 22237 1221 22295 1255
rect 22237 1187 22249 1221
rect 22283 1187 22295 1221
rect 22237 1153 22295 1187
rect 22237 1119 22249 1153
rect 22283 1119 22295 1153
rect 22237 1085 22295 1119
rect 22237 1051 22249 1085
rect 22283 1051 22295 1085
rect 22237 1017 22295 1051
rect 22237 983 22249 1017
rect 22283 983 22295 1017
rect 22237 949 22295 983
rect 22237 915 22249 949
rect 22283 915 22295 949
rect 22237 881 22295 915
rect 22237 847 22249 881
rect 22283 847 22295 881
rect 22237 813 22295 847
rect 22237 779 22249 813
rect 22283 779 22295 813
rect 22237 745 22295 779
rect 22237 711 22249 745
rect 22283 711 22295 745
rect 22237 677 22295 711
rect 22237 643 22249 677
rect 22283 643 22295 677
rect 22237 609 22295 643
rect 22237 575 22249 609
rect 22283 575 22295 609
rect 22237 541 22295 575
rect 22237 507 22249 541
rect 22283 507 22295 541
rect 22237 473 22295 507
rect 22237 439 22249 473
rect 22283 439 22295 473
rect 22237 405 22295 439
rect 22237 371 22249 405
rect 22283 371 22295 405
rect 22237 355 22295 371
rect 22695 1629 22753 1645
rect 22695 1595 22707 1629
rect 22741 1595 22753 1629
rect 22695 1561 22753 1595
rect 22695 1527 22707 1561
rect 22741 1527 22753 1561
rect 22695 1493 22753 1527
rect 22695 1459 22707 1493
rect 22741 1459 22753 1493
rect 22695 1425 22753 1459
rect 22695 1391 22707 1425
rect 22741 1391 22753 1425
rect 22695 1357 22753 1391
rect 22695 1323 22707 1357
rect 22741 1323 22753 1357
rect 22695 1289 22753 1323
rect 22695 1255 22707 1289
rect 22741 1255 22753 1289
rect 22695 1221 22753 1255
rect 22695 1187 22707 1221
rect 22741 1187 22753 1221
rect 22695 1153 22753 1187
rect 22695 1119 22707 1153
rect 22741 1119 22753 1153
rect 22695 1085 22753 1119
rect 22695 1051 22707 1085
rect 22741 1051 22753 1085
rect 22695 1017 22753 1051
rect 22695 983 22707 1017
rect 22741 983 22753 1017
rect 22695 949 22753 983
rect 22695 915 22707 949
rect 22741 915 22753 949
rect 22695 881 22753 915
rect 22695 847 22707 881
rect 22741 847 22753 881
rect 22695 813 22753 847
rect 22695 779 22707 813
rect 22741 779 22753 813
rect 22695 745 22753 779
rect 22695 711 22707 745
rect 22741 711 22753 745
rect 22695 677 22753 711
rect 22695 643 22707 677
rect 22741 643 22753 677
rect 22695 609 22753 643
rect 22695 575 22707 609
rect 22741 575 22753 609
rect 22695 541 22753 575
rect 22695 507 22707 541
rect 22741 507 22753 541
rect 22695 473 22753 507
rect 22695 439 22707 473
rect 22741 439 22753 473
rect 22695 405 22753 439
rect 22695 371 22707 405
rect 22741 371 22753 405
rect 22695 355 22753 371
rect 23153 1629 23211 1645
rect 23153 1595 23165 1629
rect 23199 1595 23211 1629
rect 23153 1561 23211 1595
rect 23153 1527 23165 1561
rect 23199 1527 23211 1561
rect 23153 1493 23211 1527
rect 23153 1459 23165 1493
rect 23199 1459 23211 1493
rect 23153 1425 23211 1459
rect 23153 1391 23165 1425
rect 23199 1391 23211 1425
rect 23153 1357 23211 1391
rect 23153 1323 23165 1357
rect 23199 1323 23211 1357
rect 23153 1289 23211 1323
rect 23153 1255 23165 1289
rect 23199 1255 23211 1289
rect 23153 1221 23211 1255
rect 23153 1187 23165 1221
rect 23199 1187 23211 1221
rect 23153 1153 23211 1187
rect 23153 1119 23165 1153
rect 23199 1119 23211 1153
rect 23153 1085 23211 1119
rect 23153 1051 23165 1085
rect 23199 1051 23211 1085
rect 23153 1017 23211 1051
rect 23153 983 23165 1017
rect 23199 983 23211 1017
rect 23153 949 23211 983
rect 23153 915 23165 949
rect 23199 915 23211 949
rect 23153 881 23211 915
rect 23153 847 23165 881
rect 23199 847 23211 881
rect 23153 813 23211 847
rect 23153 779 23165 813
rect 23199 779 23211 813
rect 23153 745 23211 779
rect 23153 711 23165 745
rect 23199 711 23211 745
rect 23153 677 23211 711
rect 23153 643 23165 677
rect 23199 643 23211 677
rect 23153 609 23211 643
rect 23153 575 23165 609
rect 23199 575 23211 609
rect 23153 541 23211 575
rect 23153 507 23165 541
rect 23199 507 23211 541
rect 23153 473 23211 507
rect 23153 439 23165 473
rect 23199 439 23211 473
rect 23153 405 23211 439
rect 23153 371 23165 405
rect 23199 371 23211 405
rect 23153 355 23211 371
rect 23611 1629 23669 1645
rect 23611 1595 23623 1629
rect 23657 1595 23669 1629
rect 23611 1561 23669 1595
rect 23611 1527 23623 1561
rect 23657 1527 23669 1561
rect 23611 1493 23669 1527
rect 23611 1459 23623 1493
rect 23657 1459 23669 1493
rect 23611 1425 23669 1459
rect 23611 1391 23623 1425
rect 23657 1391 23669 1425
rect 23611 1357 23669 1391
rect 23611 1323 23623 1357
rect 23657 1323 23669 1357
rect 23611 1289 23669 1323
rect 23611 1255 23623 1289
rect 23657 1255 23669 1289
rect 23611 1221 23669 1255
rect 23611 1187 23623 1221
rect 23657 1187 23669 1221
rect 23611 1153 23669 1187
rect 23611 1119 23623 1153
rect 23657 1119 23669 1153
rect 23611 1085 23669 1119
rect 23611 1051 23623 1085
rect 23657 1051 23669 1085
rect 23611 1017 23669 1051
rect 23611 983 23623 1017
rect 23657 983 23669 1017
rect 23611 949 23669 983
rect 23611 915 23623 949
rect 23657 915 23669 949
rect 23611 881 23669 915
rect 23611 847 23623 881
rect 23657 847 23669 881
rect 23611 813 23669 847
rect 23611 779 23623 813
rect 23657 779 23669 813
rect 23611 745 23669 779
rect 23611 711 23623 745
rect 23657 711 23669 745
rect 23611 677 23669 711
rect 23611 643 23623 677
rect 23657 643 23669 677
rect 23611 609 23669 643
rect 23611 575 23623 609
rect 23657 575 23669 609
rect 23611 541 23669 575
rect 23611 507 23623 541
rect 23657 507 23669 541
rect 23611 473 23669 507
rect 23611 439 23623 473
rect 23657 439 23669 473
rect 23611 405 23669 439
rect 23611 371 23623 405
rect 23657 371 23669 405
rect 23611 355 23669 371
rect 24069 1629 24127 1645
rect 24069 1595 24081 1629
rect 24115 1595 24127 1629
rect 24069 1561 24127 1595
rect 24069 1527 24081 1561
rect 24115 1527 24127 1561
rect 24069 1493 24127 1527
rect 24069 1459 24081 1493
rect 24115 1459 24127 1493
rect 24069 1425 24127 1459
rect 24069 1391 24081 1425
rect 24115 1391 24127 1425
rect 24069 1357 24127 1391
rect 24069 1323 24081 1357
rect 24115 1323 24127 1357
rect 24069 1289 24127 1323
rect 24069 1255 24081 1289
rect 24115 1255 24127 1289
rect 24069 1221 24127 1255
rect 24069 1187 24081 1221
rect 24115 1187 24127 1221
rect 24069 1153 24127 1187
rect 24069 1119 24081 1153
rect 24115 1119 24127 1153
rect 24069 1085 24127 1119
rect 24069 1051 24081 1085
rect 24115 1051 24127 1085
rect 24069 1017 24127 1051
rect 24069 983 24081 1017
rect 24115 983 24127 1017
rect 24069 949 24127 983
rect 24069 915 24081 949
rect 24115 915 24127 949
rect 24069 881 24127 915
rect 24069 847 24081 881
rect 24115 847 24127 881
rect 24069 813 24127 847
rect 24069 779 24081 813
rect 24115 779 24127 813
rect 24069 745 24127 779
rect 24069 711 24081 745
rect 24115 711 24127 745
rect 24069 677 24127 711
rect 24069 643 24081 677
rect 24115 643 24127 677
rect 24069 609 24127 643
rect 24069 575 24081 609
rect 24115 575 24127 609
rect 24069 541 24127 575
rect 24069 507 24081 541
rect 24115 507 24127 541
rect 24069 473 24127 507
rect 24069 439 24081 473
rect 24115 439 24127 473
rect 24069 405 24127 439
rect 24069 371 24081 405
rect 24115 371 24127 405
rect 24069 355 24127 371
rect 24527 1629 24585 1645
rect 24527 1595 24539 1629
rect 24573 1595 24585 1629
rect 24527 1561 24585 1595
rect 24527 1527 24539 1561
rect 24573 1527 24585 1561
rect 24527 1493 24585 1527
rect 24527 1459 24539 1493
rect 24573 1459 24585 1493
rect 24527 1425 24585 1459
rect 24527 1391 24539 1425
rect 24573 1391 24585 1425
rect 24527 1357 24585 1391
rect 24527 1323 24539 1357
rect 24573 1323 24585 1357
rect 24527 1289 24585 1323
rect 24527 1255 24539 1289
rect 24573 1255 24585 1289
rect 24527 1221 24585 1255
rect 24527 1187 24539 1221
rect 24573 1187 24585 1221
rect 24527 1153 24585 1187
rect 24527 1119 24539 1153
rect 24573 1119 24585 1153
rect 24527 1085 24585 1119
rect 24527 1051 24539 1085
rect 24573 1051 24585 1085
rect 24527 1017 24585 1051
rect 24527 983 24539 1017
rect 24573 983 24585 1017
rect 24527 949 24585 983
rect 24527 915 24539 949
rect 24573 915 24585 949
rect 24527 881 24585 915
rect 24527 847 24539 881
rect 24573 847 24585 881
rect 24527 813 24585 847
rect 24527 779 24539 813
rect 24573 779 24585 813
rect 24527 745 24585 779
rect 24527 711 24539 745
rect 24573 711 24585 745
rect 24527 677 24585 711
rect 24527 643 24539 677
rect 24573 643 24585 677
rect 24527 609 24585 643
rect 24527 575 24539 609
rect 24573 575 24585 609
rect 24527 541 24585 575
rect 24527 507 24539 541
rect 24573 507 24585 541
rect 24527 473 24585 507
rect 24527 439 24539 473
rect 24573 439 24585 473
rect 24527 405 24585 439
rect 24527 371 24539 405
rect 24573 371 24585 405
rect 24527 355 24585 371
rect 24985 1629 25043 1645
rect 24985 1595 24997 1629
rect 25031 1595 25043 1629
rect 24985 1561 25043 1595
rect 24985 1527 24997 1561
rect 25031 1527 25043 1561
rect 24985 1493 25043 1527
rect 24985 1459 24997 1493
rect 25031 1459 25043 1493
rect 24985 1425 25043 1459
rect 24985 1391 24997 1425
rect 25031 1391 25043 1425
rect 24985 1357 25043 1391
rect 24985 1323 24997 1357
rect 25031 1323 25043 1357
rect 24985 1289 25043 1323
rect 24985 1255 24997 1289
rect 25031 1255 25043 1289
rect 24985 1221 25043 1255
rect 24985 1187 24997 1221
rect 25031 1187 25043 1221
rect 24985 1153 25043 1187
rect 24985 1119 24997 1153
rect 25031 1119 25043 1153
rect 24985 1085 25043 1119
rect 24985 1051 24997 1085
rect 25031 1051 25043 1085
rect 24985 1017 25043 1051
rect 24985 983 24997 1017
rect 25031 983 25043 1017
rect 24985 949 25043 983
rect 24985 915 24997 949
rect 25031 915 25043 949
rect 24985 881 25043 915
rect 24985 847 24997 881
rect 25031 847 25043 881
rect 24985 813 25043 847
rect 24985 779 24997 813
rect 25031 779 25043 813
rect 24985 745 25043 779
rect 24985 711 24997 745
rect 25031 711 25043 745
rect 24985 677 25043 711
rect 24985 643 24997 677
rect 25031 643 25043 677
rect 24985 609 25043 643
rect 24985 575 24997 609
rect 25031 575 25043 609
rect 24985 541 25043 575
rect 24985 507 24997 541
rect 25031 507 25043 541
rect 24985 473 25043 507
rect 24985 439 24997 473
rect 25031 439 25043 473
rect 24985 405 25043 439
rect 24985 371 24997 405
rect 25031 371 25043 405
rect 24985 355 25043 371
rect 25443 1629 25501 1645
rect 25443 1595 25455 1629
rect 25489 1595 25501 1629
rect 25443 1561 25501 1595
rect 25443 1527 25455 1561
rect 25489 1527 25501 1561
rect 25443 1493 25501 1527
rect 25443 1459 25455 1493
rect 25489 1459 25501 1493
rect 25443 1425 25501 1459
rect 25443 1391 25455 1425
rect 25489 1391 25501 1425
rect 25443 1357 25501 1391
rect 25443 1323 25455 1357
rect 25489 1323 25501 1357
rect 25443 1289 25501 1323
rect 25443 1255 25455 1289
rect 25489 1255 25501 1289
rect 25443 1221 25501 1255
rect 25443 1187 25455 1221
rect 25489 1187 25501 1221
rect 25443 1153 25501 1187
rect 25443 1119 25455 1153
rect 25489 1119 25501 1153
rect 25443 1085 25501 1119
rect 25443 1051 25455 1085
rect 25489 1051 25501 1085
rect 25443 1017 25501 1051
rect 25443 983 25455 1017
rect 25489 983 25501 1017
rect 25443 949 25501 983
rect 25443 915 25455 949
rect 25489 915 25501 949
rect 25443 881 25501 915
rect 25443 847 25455 881
rect 25489 847 25501 881
rect 25443 813 25501 847
rect 25443 779 25455 813
rect 25489 779 25501 813
rect 25443 745 25501 779
rect 25443 711 25455 745
rect 25489 711 25501 745
rect 25443 677 25501 711
rect 25443 643 25455 677
rect 25489 643 25501 677
rect 25443 609 25501 643
rect 25443 575 25455 609
rect 25489 575 25501 609
rect 25443 541 25501 575
rect 25443 507 25455 541
rect 25489 507 25501 541
rect 25443 473 25501 507
rect 25443 439 25455 473
rect 25489 439 25501 473
rect 25443 405 25501 439
rect 25443 371 25455 405
rect 25489 371 25501 405
rect 25443 355 25501 371
rect 25901 1629 25959 1645
rect 25901 1595 25913 1629
rect 25947 1595 25959 1629
rect 25901 1561 25959 1595
rect 25901 1527 25913 1561
rect 25947 1527 25959 1561
rect 25901 1493 25959 1527
rect 25901 1459 25913 1493
rect 25947 1459 25959 1493
rect 25901 1425 25959 1459
rect 25901 1391 25913 1425
rect 25947 1391 25959 1425
rect 25901 1357 25959 1391
rect 25901 1323 25913 1357
rect 25947 1323 25959 1357
rect 25901 1289 25959 1323
rect 25901 1255 25913 1289
rect 25947 1255 25959 1289
rect 25901 1221 25959 1255
rect 25901 1187 25913 1221
rect 25947 1187 25959 1221
rect 25901 1153 25959 1187
rect 25901 1119 25913 1153
rect 25947 1119 25959 1153
rect 25901 1085 25959 1119
rect 25901 1051 25913 1085
rect 25947 1051 25959 1085
rect 25901 1017 25959 1051
rect 25901 983 25913 1017
rect 25947 983 25959 1017
rect 25901 949 25959 983
rect 25901 915 25913 949
rect 25947 915 25959 949
rect 25901 881 25959 915
rect 25901 847 25913 881
rect 25947 847 25959 881
rect 25901 813 25959 847
rect 25901 779 25913 813
rect 25947 779 25959 813
rect 25901 745 25959 779
rect 25901 711 25913 745
rect 25947 711 25959 745
rect 25901 677 25959 711
rect 25901 643 25913 677
rect 25947 643 25959 677
rect 25901 609 25959 643
rect 25901 575 25913 609
rect 25947 575 25959 609
rect 25901 541 25959 575
rect 25901 507 25913 541
rect 25947 507 25959 541
rect 25901 473 25959 507
rect 25901 439 25913 473
rect 25947 439 25959 473
rect 25901 405 25959 439
rect 25901 371 25913 405
rect 25947 371 25959 405
rect 25901 355 25959 371
rect 26359 1629 26417 1645
rect 26359 1595 26371 1629
rect 26405 1595 26417 1629
rect 26359 1561 26417 1595
rect 26359 1527 26371 1561
rect 26405 1527 26417 1561
rect 26359 1493 26417 1527
rect 26359 1459 26371 1493
rect 26405 1459 26417 1493
rect 26359 1425 26417 1459
rect 26359 1391 26371 1425
rect 26405 1391 26417 1425
rect 26359 1357 26417 1391
rect 26359 1323 26371 1357
rect 26405 1323 26417 1357
rect 26359 1289 26417 1323
rect 26359 1255 26371 1289
rect 26405 1255 26417 1289
rect 26359 1221 26417 1255
rect 26359 1187 26371 1221
rect 26405 1187 26417 1221
rect 26359 1153 26417 1187
rect 26359 1119 26371 1153
rect 26405 1119 26417 1153
rect 26359 1085 26417 1119
rect 26359 1051 26371 1085
rect 26405 1051 26417 1085
rect 26359 1017 26417 1051
rect 26359 983 26371 1017
rect 26405 983 26417 1017
rect 26359 949 26417 983
rect 26359 915 26371 949
rect 26405 915 26417 949
rect 26359 881 26417 915
rect 26359 847 26371 881
rect 26405 847 26417 881
rect 26359 813 26417 847
rect 26359 779 26371 813
rect 26405 779 26417 813
rect 26359 745 26417 779
rect 26359 711 26371 745
rect 26405 711 26417 745
rect 26359 677 26417 711
rect 26359 643 26371 677
rect 26405 643 26417 677
rect 26359 609 26417 643
rect 26359 575 26371 609
rect 26405 575 26417 609
rect 26359 541 26417 575
rect 26359 507 26371 541
rect 26405 507 26417 541
rect 26359 473 26417 507
rect 26359 439 26371 473
rect 26405 439 26417 473
rect 26359 405 26417 439
rect 26359 371 26371 405
rect 26405 371 26417 405
rect 26359 355 26417 371
rect 26817 1629 26875 1645
rect 26817 1595 26829 1629
rect 26863 1595 26875 1629
rect 26817 1561 26875 1595
rect 26817 1527 26829 1561
rect 26863 1527 26875 1561
rect 26817 1493 26875 1527
rect 26817 1459 26829 1493
rect 26863 1459 26875 1493
rect 26817 1425 26875 1459
rect 26817 1391 26829 1425
rect 26863 1391 26875 1425
rect 26817 1357 26875 1391
rect 26817 1323 26829 1357
rect 26863 1323 26875 1357
rect 26817 1289 26875 1323
rect 26817 1255 26829 1289
rect 26863 1255 26875 1289
rect 26817 1221 26875 1255
rect 26817 1187 26829 1221
rect 26863 1187 26875 1221
rect 26817 1153 26875 1187
rect 26817 1119 26829 1153
rect 26863 1119 26875 1153
rect 26817 1085 26875 1119
rect 26817 1051 26829 1085
rect 26863 1051 26875 1085
rect 26817 1017 26875 1051
rect 26817 983 26829 1017
rect 26863 983 26875 1017
rect 26817 949 26875 983
rect 26817 915 26829 949
rect 26863 915 26875 949
rect 26817 881 26875 915
rect 26817 847 26829 881
rect 26863 847 26875 881
rect 26817 813 26875 847
rect 26817 779 26829 813
rect 26863 779 26875 813
rect 26817 745 26875 779
rect 26817 711 26829 745
rect 26863 711 26875 745
rect 26817 677 26875 711
rect 26817 643 26829 677
rect 26863 643 26875 677
rect 26817 609 26875 643
rect 26817 575 26829 609
rect 26863 575 26875 609
rect 26817 541 26875 575
rect 26817 507 26829 541
rect 26863 507 26875 541
rect 26817 473 26875 507
rect 26817 439 26829 473
rect 26863 439 26875 473
rect 26817 405 26875 439
rect 26817 371 26829 405
rect 26863 371 26875 405
rect 26817 355 26875 371
rect 27275 1629 27333 1645
rect 27275 1595 27287 1629
rect 27321 1595 27333 1629
rect 27275 1561 27333 1595
rect 27275 1527 27287 1561
rect 27321 1527 27333 1561
rect 27275 1493 27333 1527
rect 27275 1459 27287 1493
rect 27321 1459 27333 1493
rect 27275 1425 27333 1459
rect 27275 1391 27287 1425
rect 27321 1391 27333 1425
rect 27275 1357 27333 1391
rect 27275 1323 27287 1357
rect 27321 1323 27333 1357
rect 27275 1289 27333 1323
rect 27275 1255 27287 1289
rect 27321 1255 27333 1289
rect 27275 1221 27333 1255
rect 27275 1187 27287 1221
rect 27321 1187 27333 1221
rect 27275 1153 27333 1187
rect 27275 1119 27287 1153
rect 27321 1119 27333 1153
rect 27275 1085 27333 1119
rect 27275 1051 27287 1085
rect 27321 1051 27333 1085
rect 27275 1017 27333 1051
rect 27275 983 27287 1017
rect 27321 983 27333 1017
rect 27275 949 27333 983
rect 27275 915 27287 949
rect 27321 915 27333 949
rect 27275 881 27333 915
rect 27275 847 27287 881
rect 27321 847 27333 881
rect 27275 813 27333 847
rect 27275 779 27287 813
rect 27321 779 27333 813
rect 27275 745 27333 779
rect 27275 711 27287 745
rect 27321 711 27333 745
rect 27275 677 27333 711
rect 27275 643 27287 677
rect 27321 643 27333 677
rect 27275 609 27333 643
rect 27275 575 27287 609
rect 27321 575 27333 609
rect 27275 541 27333 575
rect 27275 507 27287 541
rect 27321 507 27333 541
rect 27275 473 27333 507
rect 27275 439 27287 473
rect 27321 439 27333 473
rect 27275 405 27333 439
rect 27275 371 27287 405
rect 27321 371 27333 405
rect 27275 355 27333 371
rect 27733 1629 27791 1645
rect 27733 1595 27745 1629
rect 27779 1595 27791 1629
rect 27733 1561 27791 1595
rect 27733 1527 27745 1561
rect 27779 1527 27791 1561
rect 27733 1493 27791 1527
rect 27733 1459 27745 1493
rect 27779 1459 27791 1493
rect 27733 1425 27791 1459
rect 27733 1391 27745 1425
rect 27779 1391 27791 1425
rect 27733 1357 27791 1391
rect 27733 1323 27745 1357
rect 27779 1323 27791 1357
rect 27733 1289 27791 1323
rect 27733 1255 27745 1289
rect 27779 1255 27791 1289
rect 27733 1221 27791 1255
rect 27733 1187 27745 1221
rect 27779 1187 27791 1221
rect 27733 1153 27791 1187
rect 27733 1119 27745 1153
rect 27779 1119 27791 1153
rect 27733 1085 27791 1119
rect 27733 1051 27745 1085
rect 27779 1051 27791 1085
rect 27733 1017 27791 1051
rect 27733 983 27745 1017
rect 27779 983 27791 1017
rect 27733 949 27791 983
rect 27733 915 27745 949
rect 27779 915 27791 949
rect 27733 881 27791 915
rect 27733 847 27745 881
rect 27779 847 27791 881
rect 27733 813 27791 847
rect 27733 779 27745 813
rect 27779 779 27791 813
rect 27733 745 27791 779
rect 27733 711 27745 745
rect 27779 711 27791 745
rect 27733 677 27791 711
rect 27733 643 27745 677
rect 27779 643 27791 677
rect 27733 609 27791 643
rect 27733 575 27745 609
rect 27779 575 27791 609
rect 27733 541 27791 575
rect 27733 507 27745 541
rect 27779 507 27791 541
rect 27733 473 27791 507
rect 27733 439 27745 473
rect 27779 439 27791 473
rect 27733 405 27791 439
rect 27733 371 27745 405
rect 27779 371 27791 405
rect 27733 355 27791 371
<< pdiffc >>
rect 265 1595 299 1629
rect 265 1527 299 1561
rect 265 1459 299 1493
rect 265 1391 299 1425
rect 265 1323 299 1357
rect 265 1255 299 1289
rect 265 1187 299 1221
rect 265 1119 299 1153
rect 265 1051 299 1085
rect 265 983 299 1017
rect 265 915 299 949
rect 265 847 299 881
rect 265 779 299 813
rect 265 711 299 745
rect 265 643 299 677
rect 265 575 299 609
rect 265 507 299 541
rect 265 439 299 473
rect 265 371 299 405
rect 723 1595 757 1629
rect 723 1527 757 1561
rect 723 1459 757 1493
rect 723 1391 757 1425
rect 723 1323 757 1357
rect 723 1255 757 1289
rect 723 1187 757 1221
rect 723 1119 757 1153
rect 723 1051 757 1085
rect 723 983 757 1017
rect 723 915 757 949
rect 723 847 757 881
rect 723 779 757 813
rect 723 711 757 745
rect 723 643 757 677
rect 723 575 757 609
rect 723 507 757 541
rect 723 439 757 473
rect 723 371 757 405
rect 1181 1595 1215 1629
rect 1181 1527 1215 1561
rect 1181 1459 1215 1493
rect 1181 1391 1215 1425
rect 1181 1323 1215 1357
rect 1181 1255 1215 1289
rect 1181 1187 1215 1221
rect 1181 1119 1215 1153
rect 1181 1051 1215 1085
rect 1181 983 1215 1017
rect 1181 915 1215 949
rect 1181 847 1215 881
rect 1181 779 1215 813
rect 1181 711 1215 745
rect 1181 643 1215 677
rect 1181 575 1215 609
rect 1181 507 1215 541
rect 1181 439 1215 473
rect 1181 371 1215 405
rect 1639 1595 1673 1629
rect 1639 1527 1673 1561
rect 1639 1459 1673 1493
rect 1639 1391 1673 1425
rect 1639 1323 1673 1357
rect 1639 1255 1673 1289
rect 1639 1187 1673 1221
rect 1639 1119 1673 1153
rect 1639 1051 1673 1085
rect 1639 983 1673 1017
rect 1639 915 1673 949
rect 1639 847 1673 881
rect 1639 779 1673 813
rect 1639 711 1673 745
rect 1639 643 1673 677
rect 1639 575 1673 609
rect 1639 507 1673 541
rect 1639 439 1673 473
rect 1639 371 1673 405
rect 2097 1595 2131 1629
rect 2097 1527 2131 1561
rect 2097 1459 2131 1493
rect 2097 1391 2131 1425
rect 2097 1323 2131 1357
rect 2097 1255 2131 1289
rect 2097 1187 2131 1221
rect 2097 1119 2131 1153
rect 2097 1051 2131 1085
rect 2097 983 2131 1017
rect 2097 915 2131 949
rect 2097 847 2131 881
rect 2097 779 2131 813
rect 2097 711 2131 745
rect 2097 643 2131 677
rect 2097 575 2131 609
rect 2097 507 2131 541
rect 2097 439 2131 473
rect 2097 371 2131 405
rect 2555 1595 2589 1629
rect 2555 1527 2589 1561
rect 2555 1459 2589 1493
rect 2555 1391 2589 1425
rect 2555 1323 2589 1357
rect 2555 1255 2589 1289
rect 2555 1187 2589 1221
rect 2555 1119 2589 1153
rect 2555 1051 2589 1085
rect 2555 983 2589 1017
rect 2555 915 2589 949
rect 2555 847 2589 881
rect 2555 779 2589 813
rect 2555 711 2589 745
rect 2555 643 2589 677
rect 2555 575 2589 609
rect 2555 507 2589 541
rect 2555 439 2589 473
rect 2555 371 2589 405
rect 3013 1595 3047 1629
rect 3013 1527 3047 1561
rect 3013 1459 3047 1493
rect 3013 1391 3047 1425
rect 3013 1323 3047 1357
rect 3013 1255 3047 1289
rect 3013 1187 3047 1221
rect 3013 1119 3047 1153
rect 3013 1051 3047 1085
rect 3013 983 3047 1017
rect 3013 915 3047 949
rect 3013 847 3047 881
rect 3013 779 3047 813
rect 3013 711 3047 745
rect 3013 643 3047 677
rect 3013 575 3047 609
rect 3013 507 3047 541
rect 3013 439 3047 473
rect 3013 371 3047 405
rect 3471 1595 3505 1629
rect 3471 1527 3505 1561
rect 3471 1459 3505 1493
rect 3471 1391 3505 1425
rect 3471 1323 3505 1357
rect 3471 1255 3505 1289
rect 3471 1187 3505 1221
rect 3471 1119 3505 1153
rect 3471 1051 3505 1085
rect 3471 983 3505 1017
rect 3471 915 3505 949
rect 3471 847 3505 881
rect 3471 779 3505 813
rect 3471 711 3505 745
rect 3471 643 3505 677
rect 3471 575 3505 609
rect 3471 507 3505 541
rect 3471 439 3505 473
rect 3471 371 3505 405
rect 3929 1595 3963 1629
rect 3929 1527 3963 1561
rect 3929 1459 3963 1493
rect 3929 1391 3963 1425
rect 3929 1323 3963 1357
rect 3929 1255 3963 1289
rect 3929 1187 3963 1221
rect 3929 1119 3963 1153
rect 3929 1051 3963 1085
rect 3929 983 3963 1017
rect 3929 915 3963 949
rect 3929 847 3963 881
rect 3929 779 3963 813
rect 3929 711 3963 745
rect 3929 643 3963 677
rect 3929 575 3963 609
rect 3929 507 3963 541
rect 3929 439 3963 473
rect 3929 371 3963 405
rect 4387 1595 4421 1629
rect 4387 1527 4421 1561
rect 4387 1459 4421 1493
rect 4387 1391 4421 1425
rect 4387 1323 4421 1357
rect 4387 1255 4421 1289
rect 4387 1187 4421 1221
rect 4387 1119 4421 1153
rect 4387 1051 4421 1085
rect 4387 983 4421 1017
rect 4387 915 4421 949
rect 4387 847 4421 881
rect 4387 779 4421 813
rect 4387 711 4421 745
rect 4387 643 4421 677
rect 4387 575 4421 609
rect 4387 507 4421 541
rect 4387 439 4421 473
rect 4387 371 4421 405
rect 4845 1595 4879 1629
rect 4845 1527 4879 1561
rect 4845 1459 4879 1493
rect 4845 1391 4879 1425
rect 4845 1323 4879 1357
rect 4845 1255 4879 1289
rect 4845 1187 4879 1221
rect 4845 1119 4879 1153
rect 4845 1051 4879 1085
rect 4845 983 4879 1017
rect 4845 915 4879 949
rect 4845 847 4879 881
rect 4845 779 4879 813
rect 4845 711 4879 745
rect 4845 643 4879 677
rect 4845 575 4879 609
rect 4845 507 4879 541
rect 4845 439 4879 473
rect 4845 371 4879 405
rect 5303 1595 5337 1629
rect 5303 1527 5337 1561
rect 5303 1459 5337 1493
rect 5303 1391 5337 1425
rect 5303 1323 5337 1357
rect 5303 1255 5337 1289
rect 5303 1187 5337 1221
rect 5303 1119 5337 1153
rect 5303 1051 5337 1085
rect 5303 983 5337 1017
rect 5303 915 5337 949
rect 5303 847 5337 881
rect 5303 779 5337 813
rect 5303 711 5337 745
rect 5303 643 5337 677
rect 5303 575 5337 609
rect 5303 507 5337 541
rect 5303 439 5337 473
rect 5303 371 5337 405
rect 5761 1595 5795 1629
rect 5761 1527 5795 1561
rect 5761 1459 5795 1493
rect 5761 1391 5795 1425
rect 5761 1323 5795 1357
rect 5761 1255 5795 1289
rect 5761 1187 5795 1221
rect 5761 1119 5795 1153
rect 5761 1051 5795 1085
rect 5761 983 5795 1017
rect 5761 915 5795 949
rect 5761 847 5795 881
rect 5761 779 5795 813
rect 5761 711 5795 745
rect 5761 643 5795 677
rect 5761 575 5795 609
rect 5761 507 5795 541
rect 5761 439 5795 473
rect 5761 371 5795 405
rect 6219 1595 6253 1629
rect 6219 1527 6253 1561
rect 6219 1459 6253 1493
rect 6219 1391 6253 1425
rect 6219 1323 6253 1357
rect 6219 1255 6253 1289
rect 6219 1187 6253 1221
rect 6219 1119 6253 1153
rect 6219 1051 6253 1085
rect 6219 983 6253 1017
rect 6219 915 6253 949
rect 6219 847 6253 881
rect 6219 779 6253 813
rect 6219 711 6253 745
rect 6219 643 6253 677
rect 6219 575 6253 609
rect 6219 507 6253 541
rect 6219 439 6253 473
rect 6219 371 6253 405
rect 6677 1595 6711 1629
rect 6677 1527 6711 1561
rect 6677 1459 6711 1493
rect 6677 1391 6711 1425
rect 6677 1323 6711 1357
rect 6677 1255 6711 1289
rect 6677 1187 6711 1221
rect 6677 1119 6711 1153
rect 6677 1051 6711 1085
rect 6677 983 6711 1017
rect 6677 915 6711 949
rect 6677 847 6711 881
rect 6677 779 6711 813
rect 6677 711 6711 745
rect 6677 643 6711 677
rect 6677 575 6711 609
rect 6677 507 6711 541
rect 6677 439 6711 473
rect 6677 371 6711 405
rect 7135 1595 7169 1629
rect 7135 1527 7169 1561
rect 7135 1459 7169 1493
rect 7135 1391 7169 1425
rect 7135 1323 7169 1357
rect 7135 1255 7169 1289
rect 7135 1187 7169 1221
rect 7135 1119 7169 1153
rect 7135 1051 7169 1085
rect 7135 983 7169 1017
rect 7135 915 7169 949
rect 7135 847 7169 881
rect 7135 779 7169 813
rect 7135 711 7169 745
rect 7135 643 7169 677
rect 7135 575 7169 609
rect 7135 507 7169 541
rect 7135 439 7169 473
rect 7135 371 7169 405
rect 7593 1595 7627 1629
rect 7593 1527 7627 1561
rect 7593 1459 7627 1493
rect 7593 1391 7627 1425
rect 7593 1323 7627 1357
rect 7593 1255 7627 1289
rect 7593 1187 7627 1221
rect 7593 1119 7627 1153
rect 7593 1051 7627 1085
rect 7593 983 7627 1017
rect 7593 915 7627 949
rect 7593 847 7627 881
rect 7593 779 7627 813
rect 7593 711 7627 745
rect 7593 643 7627 677
rect 7593 575 7627 609
rect 7593 507 7627 541
rect 7593 439 7627 473
rect 7593 371 7627 405
rect 8051 1595 8085 1629
rect 8051 1527 8085 1561
rect 8051 1459 8085 1493
rect 8051 1391 8085 1425
rect 8051 1323 8085 1357
rect 8051 1255 8085 1289
rect 8051 1187 8085 1221
rect 8051 1119 8085 1153
rect 8051 1051 8085 1085
rect 8051 983 8085 1017
rect 8051 915 8085 949
rect 8051 847 8085 881
rect 8051 779 8085 813
rect 8051 711 8085 745
rect 8051 643 8085 677
rect 8051 575 8085 609
rect 8051 507 8085 541
rect 8051 439 8085 473
rect 8051 371 8085 405
rect 8509 1595 8543 1629
rect 8509 1527 8543 1561
rect 8509 1459 8543 1493
rect 8509 1391 8543 1425
rect 8509 1323 8543 1357
rect 8509 1255 8543 1289
rect 8509 1187 8543 1221
rect 8509 1119 8543 1153
rect 8509 1051 8543 1085
rect 8509 983 8543 1017
rect 8509 915 8543 949
rect 8509 847 8543 881
rect 8509 779 8543 813
rect 8509 711 8543 745
rect 8509 643 8543 677
rect 8509 575 8543 609
rect 8509 507 8543 541
rect 8509 439 8543 473
rect 8509 371 8543 405
rect 8967 1595 9001 1629
rect 8967 1527 9001 1561
rect 8967 1459 9001 1493
rect 8967 1391 9001 1425
rect 8967 1323 9001 1357
rect 8967 1255 9001 1289
rect 8967 1187 9001 1221
rect 8967 1119 9001 1153
rect 8967 1051 9001 1085
rect 8967 983 9001 1017
rect 8967 915 9001 949
rect 8967 847 9001 881
rect 8967 779 9001 813
rect 8967 711 9001 745
rect 8967 643 9001 677
rect 8967 575 9001 609
rect 8967 507 9001 541
rect 8967 439 9001 473
rect 8967 371 9001 405
rect 9425 1595 9459 1629
rect 9425 1527 9459 1561
rect 9425 1459 9459 1493
rect 9425 1391 9459 1425
rect 9425 1323 9459 1357
rect 9425 1255 9459 1289
rect 9425 1187 9459 1221
rect 9425 1119 9459 1153
rect 9425 1051 9459 1085
rect 9425 983 9459 1017
rect 9425 915 9459 949
rect 9425 847 9459 881
rect 9425 779 9459 813
rect 9425 711 9459 745
rect 9425 643 9459 677
rect 9425 575 9459 609
rect 9425 507 9459 541
rect 9425 439 9459 473
rect 9425 371 9459 405
rect 9883 1595 9917 1629
rect 9883 1527 9917 1561
rect 9883 1459 9917 1493
rect 9883 1391 9917 1425
rect 9883 1323 9917 1357
rect 9883 1255 9917 1289
rect 9883 1187 9917 1221
rect 9883 1119 9917 1153
rect 9883 1051 9917 1085
rect 9883 983 9917 1017
rect 9883 915 9917 949
rect 9883 847 9917 881
rect 9883 779 9917 813
rect 9883 711 9917 745
rect 9883 643 9917 677
rect 9883 575 9917 609
rect 9883 507 9917 541
rect 9883 439 9917 473
rect 9883 371 9917 405
rect 10341 1595 10375 1629
rect 10341 1527 10375 1561
rect 10341 1459 10375 1493
rect 10341 1391 10375 1425
rect 10341 1323 10375 1357
rect 10341 1255 10375 1289
rect 10341 1187 10375 1221
rect 10341 1119 10375 1153
rect 10341 1051 10375 1085
rect 10341 983 10375 1017
rect 10341 915 10375 949
rect 10341 847 10375 881
rect 10341 779 10375 813
rect 10341 711 10375 745
rect 10341 643 10375 677
rect 10341 575 10375 609
rect 10341 507 10375 541
rect 10341 439 10375 473
rect 10341 371 10375 405
rect 10799 1595 10833 1629
rect 10799 1527 10833 1561
rect 10799 1459 10833 1493
rect 10799 1391 10833 1425
rect 10799 1323 10833 1357
rect 10799 1255 10833 1289
rect 10799 1187 10833 1221
rect 10799 1119 10833 1153
rect 10799 1051 10833 1085
rect 10799 983 10833 1017
rect 10799 915 10833 949
rect 10799 847 10833 881
rect 10799 779 10833 813
rect 10799 711 10833 745
rect 10799 643 10833 677
rect 10799 575 10833 609
rect 10799 507 10833 541
rect 10799 439 10833 473
rect 10799 371 10833 405
rect 11257 1595 11291 1629
rect 11257 1527 11291 1561
rect 11257 1459 11291 1493
rect 11257 1391 11291 1425
rect 11257 1323 11291 1357
rect 11257 1255 11291 1289
rect 11257 1187 11291 1221
rect 11257 1119 11291 1153
rect 11257 1051 11291 1085
rect 11257 983 11291 1017
rect 11257 915 11291 949
rect 11257 847 11291 881
rect 11257 779 11291 813
rect 11257 711 11291 745
rect 11257 643 11291 677
rect 11257 575 11291 609
rect 11257 507 11291 541
rect 11257 439 11291 473
rect 11257 371 11291 405
rect 11715 1595 11749 1629
rect 11715 1527 11749 1561
rect 11715 1459 11749 1493
rect 11715 1391 11749 1425
rect 11715 1323 11749 1357
rect 11715 1255 11749 1289
rect 11715 1187 11749 1221
rect 11715 1119 11749 1153
rect 11715 1051 11749 1085
rect 11715 983 11749 1017
rect 11715 915 11749 949
rect 11715 847 11749 881
rect 11715 779 11749 813
rect 11715 711 11749 745
rect 11715 643 11749 677
rect 11715 575 11749 609
rect 11715 507 11749 541
rect 11715 439 11749 473
rect 11715 371 11749 405
rect 12173 1595 12207 1629
rect 12173 1527 12207 1561
rect 12173 1459 12207 1493
rect 12173 1391 12207 1425
rect 12173 1323 12207 1357
rect 12173 1255 12207 1289
rect 12173 1187 12207 1221
rect 12173 1119 12207 1153
rect 12173 1051 12207 1085
rect 12173 983 12207 1017
rect 12173 915 12207 949
rect 12173 847 12207 881
rect 12173 779 12207 813
rect 12173 711 12207 745
rect 12173 643 12207 677
rect 12173 575 12207 609
rect 12173 507 12207 541
rect 12173 439 12207 473
rect 12173 371 12207 405
rect 12631 1595 12665 1629
rect 12631 1527 12665 1561
rect 12631 1459 12665 1493
rect 12631 1391 12665 1425
rect 12631 1323 12665 1357
rect 12631 1255 12665 1289
rect 12631 1187 12665 1221
rect 12631 1119 12665 1153
rect 12631 1051 12665 1085
rect 12631 983 12665 1017
rect 12631 915 12665 949
rect 12631 847 12665 881
rect 12631 779 12665 813
rect 12631 711 12665 745
rect 12631 643 12665 677
rect 12631 575 12665 609
rect 12631 507 12665 541
rect 12631 439 12665 473
rect 12631 371 12665 405
rect 13089 1595 13123 1629
rect 13089 1527 13123 1561
rect 13089 1459 13123 1493
rect 13089 1391 13123 1425
rect 13089 1323 13123 1357
rect 13089 1255 13123 1289
rect 13089 1187 13123 1221
rect 13089 1119 13123 1153
rect 13089 1051 13123 1085
rect 13089 983 13123 1017
rect 13089 915 13123 949
rect 13089 847 13123 881
rect 13089 779 13123 813
rect 13089 711 13123 745
rect 13089 643 13123 677
rect 13089 575 13123 609
rect 13089 507 13123 541
rect 13089 439 13123 473
rect 13089 371 13123 405
rect 13547 1595 13581 1629
rect 13547 1527 13581 1561
rect 13547 1459 13581 1493
rect 13547 1391 13581 1425
rect 13547 1323 13581 1357
rect 13547 1255 13581 1289
rect 13547 1187 13581 1221
rect 13547 1119 13581 1153
rect 13547 1051 13581 1085
rect 13547 983 13581 1017
rect 13547 915 13581 949
rect 13547 847 13581 881
rect 13547 779 13581 813
rect 13547 711 13581 745
rect 13547 643 13581 677
rect 13547 575 13581 609
rect 13547 507 13581 541
rect 13547 439 13581 473
rect 13547 371 13581 405
rect 14005 1595 14039 1629
rect 14005 1527 14039 1561
rect 14005 1459 14039 1493
rect 14005 1391 14039 1425
rect 14005 1323 14039 1357
rect 14005 1255 14039 1289
rect 14005 1187 14039 1221
rect 14005 1119 14039 1153
rect 14005 1051 14039 1085
rect 14005 983 14039 1017
rect 14005 915 14039 949
rect 14005 847 14039 881
rect 14005 779 14039 813
rect 14005 711 14039 745
rect 14005 643 14039 677
rect 14005 575 14039 609
rect 14005 507 14039 541
rect 14005 439 14039 473
rect 14005 371 14039 405
rect 14463 1595 14497 1629
rect 14463 1527 14497 1561
rect 14463 1459 14497 1493
rect 14463 1391 14497 1425
rect 14463 1323 14497 1357
rect 14463 1255 14497 1289
rect 14463 1187 14497 1221
rect 14463 1119 14497 1153
rect 14463 1051 14497 1085
rect 14463 983 14497 1017
rect 14463 915 14497 949
rect 14463 847 14497 881
rect 14463 779 14497 813
rect 14463 711 14497 745
rect 14463 643 14497 677
rect 14463 575 14497 609
rect 14463 507 14497 541
rect 14463 439 14497 473
rect 14463 371 14497 405
rect 14921 1595 14955 1629
rect 14921 1527 14955 1561
rect 14921 1459 14955 1493
rect 14921 1391 14955 1425
rect 14921 1323 14955 1357
rect 14921 1255 14955 1289
rect 14921 1187 14955 1221
rect 14921 1119 14955 1153
rect 14921 1051 14955 1085
rect 14921 983 14955 1017
rect 14921 915 14955 949
rect 14921 847 14955 881
rect 14921 779 14955 813
rect 14921 711 14955 745
rect 14921 643 14955 677
rect 14921 575 14955 609
rect 14921 507 14955 541
rect 14921 439 14955 473
rect 14921 371 14955 405
rect 15379 1595 15413 1629
rect 15379 1527 15413 1561
rect 15379 1459 15413 1493
rect 15379 1391 15413 1425
rect 15379 1323 15413 1357
rect 15379 1255 15413 1289
rect 15379 1187 15413 1221
rect 15379 1119 15413 1153
rect 15379 1051 15413 1085
rect 15379 983 15413 1017
rect 15379 915 15413 949
rect 15379 847 15413 881
rect 15379 779 15413 813
rect 15379 711 15413 745
rect 15379 643 15413 677
rect 15379 575 15413 609
rect 15379 507 15413 541
rect 15379 439 15413 473
rect 15379 371 15413 405
rect 15837 1595 15871 1629
rect 15837 1527 15871 1561
rect 15837 1459 15871 1493
rect 15837 1391 15871 1425
rect 15837 1323 15871 1357
rect 15837 1255 15871 1289
rect 15837 1187 15871 1221
rect 15837 1119 15871 1153
rect 15837 1051 15871 1085
rect 15837 983 15871 1017
rect 15837 915 15871 949
rect 15837 847 15871 881
rect 15837 779 15871 813
rect 15837 711 15871 745
rect 15837 643 15871 677
rect 15837 575 15871 609
rect 15837 507 15871 541
rect 15837 439 15871 473
rect 15837 371 15871 405
rect 16295 1595 16329 1629
rect 16295 1527 16329 1561
rect 16295 1459 16329 1493
rect 16295 1391 16329 1425
rect 16295 1323 16329 1357
rect 16295 1255 16329 1289
rect 16295 1187 16329 1221
rect 16295 1119 16329 1153
rect 16295 1051 16329 1085
rect 16295 983 16329 1017
rect 16295 915 16329 949
rect 16295 847 16329 881
rect 16295 779 16329 813
rect 16295 711 16329 745
rect 16295 643 16329 677
rect 16295 575 16329 609
rect 16295 507 16329 541
rect 16295 439 16329 473
rect 16295 371 16329 405
rect 16753 1595 16787 1629
rect 16753 1527 16787 1561
rect 16753 1459 16787 1493
rect 16753 1391 16787 1425
rect 16753 1323 16787 1357
rect 16753 1255 16787 1289
rect 16753 1187 16787 1221
rect 16753 1119 16787 1153
rect 16753 1051 16787 1085
rect 16753 983 16787 1017
rect 16753 915 16787 949
rect 16753 847 16787 881
rect 16753 779 16787 813
rect 16753 711 16787 745
rect 16753 643 16787 677
rect 16753 575 16787 609
rect 16753 507 16787 541
rect 16753 439 16787 473
rect 16753 371 16787 405
rect 17211 1595 17245 1629
rect 17211 1527 17245 1561
rect 17211 1459 17245 1493
rect 17211 1391 17245 1425
rect 17211 1323 17245 1357
rect 17211 1255 17245 1289
rect 17211 1187 17245 1221
rect 17211 1119 17245 1153
rect 17211 1051 17245 1085
rect 17211 983 17245 1017
rect 17211 915 17245 949
rect 17211 847 17245 881
rect 17211 779 17245 813
rect 17211 711 17245 745
rect 17211 643 17245 677
rect 17211 575 17245 609
rect 17211 507 17245 541
rect 17211 439 17245 473
rect 17211 371 17245 405
rect 17669 1595 17703 1629
rect 17669 1527 17703 1561
rect 17669 1459 17703 1493
rect 17669 1391 17703 1425
rect 17669 1323 17703 1357
rect 17669 1255 17703 1289
rect 17669 1187 17703 1221
rect 17669 1119 17703 1153
rect 17669 1051 17703 1085
rect 17669 983 17703 1017
rect 17669 915 17703 949
rect 17669 847 17703 881
rect 17669 779 17703 813
rect 17669 711 17703 745
rect 17669 643 17703 677
rect 17669 575 17703 609
rect 17669 507 17703 541
rect 17669 439 17703 473
rect 17669 371 17703 405
rect 18127 1595 18161 1629
rect 18127 1527 18161 1561
rect 18127 1459 18161 1493
rect 18127 1391 18161 1425
rect 18127 1323 18161 1357
rect 18127 1255 18161 1289
rect 18127 1187 18161 1221
rect 18127 1119 18161 1153
rect 18127 1051 18161 1085
rect 18127 983 18161 1017
rect 18127 915 18161 949
rect 18127 847 18161 881
rect 18127 779 18161 813
rect 18127 711 18161 745
rect 18127 643 18161 677
rect 18127 575 18161 609
rect 18127 507 18161 541
rect 18127 439 18161 473
rect 18127 371 18161 405
rect 18585 1595 18619 1629
rect 18585 1527 18619 1561
rect 18585 1459 18619 1493
rect 18585 1391 18619 1425
rect 18585 1323 18619 1357
rect 18585 1255 18619 1289
rect 18585 1187 18619 1221
rect 18585 1119 18619 1153
rect 18585 1051 18619 1085
rect 18585 983 18619 1017
rect 18585 915 18619 949
rect 18585 847 18619 881
rect 18585 779 18619 813
rect 18585 711 18619 745
rect 18585 643 18619 677
rect 18585 575 18619 609
rect 18585 507 18619 541
rect 18585 439 18619 473
rect 18585 371 18619 405
rect 19043 1595 19077 1629
rect 19043 1527 19077 1561
rect 19043 1459 19077 1493
rect 19043 1391 19077 1425
rect 19043 1323 19077 1357
rect 19043 1255 19077 1289
rect 19043 1187 19077 1221
rect 19043 1119 19077 1153
rect 19043 1051 19077 1085
rect 19043 983 19077 1017
rect 19043 915 19077 949
rect 19043 847 19077 881
rect 19043 779 19077 813
rect 19043 711 19077 745
rect 19043 643 19077 677
rect 19043 575 19077 609
rect 19043 507 19077 541
rect 19043 439 19077 473
rect 19043 371 19077 405
rect 19501 1595 19535 1629
rect 19501 1527 19535 1561
rect 19501 1459 19535 1493
rect 19501 1391 19535 1425
rect 19501 1323 19535 1357
rect 19501 1255 19535 1289
rect 19501 1187 19535 1221
rect 19501 1119 19535 1153
rect 19501 1051 19535 1085
rect 19501 983 19535 1017
rect 19501 915 19535 949
rect 19501 847 19535 881
rect 19501 779 19535 813
rect 19501 711 19535 745
rect 19501 643 19535 677
rect 19501 575 19535 609
rect 19501 507 19535 541
rect 19501 439 19535 473
rect 19501 371 19535 405
rect 19959 1595 19993 1629
rect 19959 1527 19993 1561
rect 19959 1459 19993 1493
rect 19959 1391 19993 1425
rect 19959 1323 19993 1357
rect 19959 1255 19993 1289
rect 19959 1187 19993 1221
rect 19959 1119 19993 1153
rect 19959 1051 19993 1085
rect 19959 983 19993 1017
rect 19959 915 19993 949
rect 19959 847 19993 881
rect 19959 779 19993 813
rect 19959 711 19993 745
rect 19959 643 19993 677
rect 19959 575 19993 609
rect 19959 507 19993 541
rect 19959 439 19993 473
rect 19959 371 19993 405
rect 20417 1595 20451 1629
rect 20417 1527 20451 1561
rect 20417 1459 20451 1493
rect 20417 1391 20451 1425
rect 20417 1323 20451 1357
rect 20417 1255 20451 1289
rect 20417 1187 20451 1221
rect 20417 1119 20451 1153
rect 20417 1051 20451 1085
rect 20417 983 20451 1017
rect 20417 915 20451 949
rect 20417 847 20451 881
rect 20417 779 20451 813
rect 20417 711 20451 745
rect 20417 643 20451 677
rect 20417 575 20451 609
rect 20417 507 20451 541
rect 20417 439 20451 473
rect 20417 371 20451 405
rect 20875 1595 20909 1629
rect 20875 1527 20909 1561
rect 20875 1459 20909 1493
rect 20875 1391 20909 1425
rect 20875 1323 20909 1357
rect 20875 1255 20909 1289
rect 20875 1187 20909 1221
rect 20875 1119 20909 1153
rect 20875 1051 20909 1085
rect 20875 983 20909 1017
rect 20875 915 20909 949
rect 20875 847 20909 881
rect 20875 779 20909 813
rect 20875 711 20909 745
rect 20875 643 20909 677
rect 20875 575 20909 609
rect 20875 507 20909 541
rect 20875 439 20909 473
rect 20875 371 20909 405
rect 21333 1595 21367 1629
rect 21333 1527 21367 1561
rect 21333 1459 21367 1493
rect 21333 1391 21367 1425
rect 21333 1323 21367 1357
rect 21333 1255 21367 1289
rect 21333 1187 21367 1221
rect 21333 1119 21367 1153
rect 21333 1051 21367 1085
rect 21333 983 21367 1017
rect 21333 915 21367 949
rect 21333 847 21367 881
rect 21333 779 21367 813
rect 21333 711 21367 745
rect 21333 643 21367 677
rect 21333 575 21367 609
rect 21333 507 21367 541
rect 21333 439 21367 473
rect 21333 371 21367 405
rect 21791 1595 21825 1629
rect 21791 1527 21825 1561
rect 21791 1459 21825 1493
rect 21791 1391 21825 1425
rect 21791 1323 21825 1357
rect 21791 1255 21825 1289
rect 21791 1187 21825 1221
rect 21791 1119 21825 1153
rect 21791 1051 21825 1085
rect 21791 983 21825 1017
rect 21791 915 21825 949
rect 21791 847 21825 881
rect 21791 779 21825 813
rect 21791 711 21825 745
rect 21791 643 21825 677
rect 21791 575 21825 609
rect 21791 507 21825 541
rect 21791 439 21825 473
rect 21791 371 21825 405
rect 22249 1595 22283 1629
rect 22249 1527 22283 1561
rect 22249 1459 22283 1493
rect 22249 1391 22283 1425
rect 22249 1323 22283 1357
rect 22249 1255 22283 1289
rect 22249 1187 22283 1221
rect 22249 1119 22283 1153
rect 22249 1051 22283 1085
rect 22249 983 22283 1017
rect 22249 915 22283 949
rect 22249 847 22283 881
rect 22249 779 22283 813
rect 22249 711 22283 745
rect 22249 643 22283 677
rect 22249 575 22283 609
rect 22249 507 22283 541
rect 22249 439 22283 473
rect 22249 371 22283 405
rect 22707 1595 22741 1629
rect 22707 1527 22741 1561
rect 22707 1459 22741 1493
rect 22707 1391 22741 1425
rect 22707 1323 22741 1357
rect 22707 1255 22741 1289
rect 22707 1187 22741 1221
rect 22707 1119 22741 1153
rect 22707 1051 22741 1085
rect 22707 983 22741 1017
rect 22707 915 22741 949
rect 22707 847 22741 881
rect 22707 779 22741 813
rect 22707 711 22741 745
rect 22707 643 22741 677
rect 22707 575 22741 609
rect 22707 507 22741 541
rect 22707 439 22741 473
rect 22707 371 22741 405
rect 23165 1595 23199 1629
rect 23165 1527 23199 1561
rect 23165 1459 23199 1493
rect 23165 1391 23199 1425
rect 23165 1323 23199 1357
rect 23165 1255 23199 1289
rect 23165 1187 23199 1221
rect 23165 1119 23199 1153
rect 23165 1051 23199 1085
rect 23165 983 23199 1017
rect 23165 915 23199 949
rect 23165 847 23199 881
rect 23165 779 23199 813
rect 23165 711 23199 745
rect 23165 643 23199 677
rect 23165 575 23199 609
rect 23165 507 23199 541
rect 23165 439 23199 473
rect 23165 371 23199 405
rect 23623 1595 23657 1629
rect 23623 1527 23657 1561
rect 23623 1459 23657 1493
rect 23623 1391 23657 1425
rect 23623 1323 23657 1357
rect 23623 1255 23657 1289
rect 23623 1187 23657 1221
rect 23623 1119 23657 1153
rect 23623 1051 23657 1085
rect 23623 983 23657 1017
rect 23623 915 23657 949
rect 23623 847 23657 881
rect 23623 779 23657 813
rect 23623 711 23657 745
rect 23623 643 23657 677
rect 23623 575 23657 609
rect 23623 507 23657 541
rect 23623 439 23657 473
rect 23623 371 23657 405
rect 24081 1595 24115 1629
rect 24081 1527 24115 1561
rect 24081 1459 24115 1493
rect 24081 1391 24115 1425
rect 24081 1323 24115 1357
rect 24081 1255 24115 1289
rect 24081 1187 24115 1221
rect 24081 1119 24115 1153
rect 24081 1051 24115 1085
rect 24081 983 24115 1017
rect 24081 915 24115 949
rect 24081 847 24115 881
rect 24081 779 24115 813
rect 24081 711 24115 745
rect 24081 643 24115 677
rect 24081 575 24115 609
rect 24081 507 24115 541
rect 24081 439 24115 473
rect 24081 371 24115 405
rect 24539 1595 24573 1629
rect 24539 1527 24573 1561
rect 24539 1459 24573 1493
rect 24539 1391 24573 1425
rect 24539 1323 24573 1357
rect 24539 1255 24573 1289
rect 24539 1187 24573 1221
rect 24539 1119 24573 1153
rect 24539 1051 24573 1085
rect 24539 983 24573 1017
rect 24539 915 24573 949
rect 24539 847 24573 881
rect 24539 779 24573 813
rect 24539 711 24573 745
rect 24539 643 24573 677
rect 24539 575 24573 609
rect 24539 507 24573 541
rect 24539 439 24573 473
rect 24539 371 24573 405
rect 24997 1595 25031 1629
rect 24997 1527 25031 1561
rect 24997 1459 25031 1493
rect 24997 1391 25031 1425
rect 24997 1323 25031 1357
rect 24997 1255 25031 1289
rect 24997 1187 25031 1221
rect 24997 1119 25031 1153
rect 24997 1051 25031 1085
rect 24997 983 25031 1017
rect 24997 915 25031 949
rect 24997 847 25031 881
rect 24997 779 25031 813
rect 24997 711 25031 745
rect 24997 643 25031 677
rect 24997 575 25031 609
rect 24997 507 25031 541
rect 24997 439 25031 473
rect 24997 371 25031 405
rect 25455 1595 25489 1629
rect 25455 1527 25489 1561
rect 25455 1459 25489 1493
rect 25455 1391 25489 1425
rect 25455 1323 25489 1357
rect 25455 1255 25489 1289
rect 25455 1187 25489 1221
rect 25455 1119 25489 1153
rect 25455 1051 25489 1085
rect 25455 983 25489 1017
rect 25455 915 25489 949
rect 25455 847 25489 881
rect 25455 779 25489 813
rect 25455 711 25489 745
rect 25455 643 25489 677
rect 25455 575 25489 609
rect 25455 507 25489 541
rect 25455 439 25489 473
rect 25455 371 25489 405
rect 25913 1595 25947 1629
rect 25913 1527 25947 1561
rect 25913 1459 25947 1493
rect 25913 1391 25947 1425
rect 25913 1323 25947 1357
rect 25913 1255 25947 1289
rect 25913 1187 25947 1221
rect 25913 1119 25947 1153
rect 25913 1051 25947 1085
rect 25913 983 25947 1017
rect 25913 915 25947 949
rect 25913 847 25947 881
rect 25913 779 25947 813
rect 25913 711 25947 745
rect 25913 643 25947 677
rect 25913 575 25947 609
rect 25913 507 25947 541
rect 25913 439 25947 473
rect 25913 371 25947 405
rect 26371 1595 26405 1629
rect 26371 1527 26405 1561
rect 26371 1459 26405 1493
rect 26371 1391 26405 1425
rect 26371 1323 26405 1357
rect 26371 1255 26405 1289
rect 26371 1187 26405 1221
rect 26371 1119 26405 1153
rect 26371 1051 26405 1085
rect 26371 983 26405 1017
rect 26371 915 26405 949
rect 26371 847 26405 881
rect 26371 779 26405 813
rect 26371 711 26405 745
rect 26371 643 26405 677
rect 26371 575 26405 609
rect 26371 507 26405 541
rect 26371 439 26405 473
rect 26371 371 26405 405
rect 26829 1595 26863 1629
rect 26829 1527 26863 1561
rect 26829 1459 26863 1493
rect 26829 1391 26863 1425
rect 26829 1323 26863 1357
rect 26829 1255 26863 1289
rect 26829 1187 26863 1221
rect 26829 1119 26863 1153
rect 26829 1051 26863 1085
rect 26829 983 26863 1017
rect 26829 915 26863 949
rect 26829 847 26863 881
rect 26829 779 26863 813
rect 26829 711 26863 745
rect 26829 643 26863 677
rect 26829 575 26863 609
rect 26829 507 26863 541
rect 26829 439 26863 473
rect 26829 371 26863 405
rect 27287 1595 27321 1629
rect 27287 1527 27321 1561
rect 27287 1459 27321 1493
rect 27287 1391 27321 1425
rect 27287 1323 27321 1357
rect 27287 1255 27321 1289
rect 27287 1187 27321 1221
rect 27287 1119 27321 1153
rect 27287 1051 27321 1085
rect 27287 983 27321 1017
rect 27287 915 27321 949
rect 27287 847 27321 881
rect 27287 779 27321 813
rect 27287 711 27321 745
rect 27287 643 27321 677
rect 27287 575 27321 609
rect 27287 507 27321 541
rect 27287 439 27321 473
rect 27287 371 27321 405
rect 27745 1595 27779 1629
rect 27745 1527 27779 1561
rect 27745 1459 27779 1493
rect 27745 1391 27779 1425
rect 27745 1323 27779 1357
rect 27745 1255 27779 1289
rect 27745 1187 27779 1221
rect 27745 1119 27779 1153
rect 27745 1051 27779 1085
rect 27745 983 27779 1017
rect 27745 915 27779 949
rect 27745 847 27779 881
rect 27745 779 27779 813
rect 27745 711 27779 745
rect 27745 643 27779 677
rect 27745 575 27779 609
rect 27745 507 27779 541
rect 27745 439 27779 473
rect 27745 371 27779 405
<< nsubdiff >>
rect 1216 1807 1336 1810
rect 158 1757 198 1800
rect 1216 1773 1261 1807
rect 1295 1773 1336 1807
rect 1216 1770 1336 1773
rect 2516 1807 2636 1810
rect 2516 1773 2561 1807
rect 2595 1773 2636 1807
rect 2516 1770 2636 1773
rect 3816 1807 3936 1810
rect 3816 1773 3861 1807
rect 3895 1773 3936 1807
rect 3816 1770 3936 1773
rect 5116 1807 5236 1810
rect 5116 1773 5161 1807
rect 5195 1773 5236 1807
rect 5116 1770 5236 1773
rect 6416 1807 6536 1810
rect 6416 1773 6461 1807
rect 6495 1773 6536 1807
rect 6416 1770 6536 1773
rect 7716 1807 7836 1810
rect 7716 1773 7761 1807
rect 7795 1773 7836 1807
rect 7716 1770 7836 1773
rect 9016 1807 9136 1810
rect 9016 1773 9061 1807
rect 9095 1773 9136 1807
rect 9016 1770 9136 1773
rect 10316 1807 10436 1810
rect 10316 1773 10361 1807
rect 10395 1773 10436 1807
rect 10316 1770 10436 1773
rect 11616 1807 11736 1810
rect 11616 1773 11661 1807
rect 11695 1773 11736 1807
rect 11616 1770 11736 1773
rect 12916 1807 13036 1810
rect 12916 1773 12961 1807
rect 12995 1773 13036 1807
rect 12916 1770 13036 1773
rect 14216 1807 14336 1810
rect 14216 1773 14261 1807
rect 14295 1773 14336 1807
rect 14216 1770 14336 1773
rect 15516 1807 15636 1810
rect 15516 1773 15561 1807
rect 15595 1773 15636 1807
rect 15516 1770 15636 1773
rect 16816 1807 16936 1810
rect 16816 1773 16861 1807
rect 16895 1773 16936 1807
rect 16816 1770 16936 1773
rect 18116 1807 18236 1810
rect 18116 1773 18161 1807
rect 18195 1773 18236 1807
rect 18116 1770 18236 1773
rect 19416 1807 19536 1810
rect 19416 1773 19461 1807
rect 19495 1773 19536 1807
rect 19416 1770 19536 1773
rect 20716 1807 20836 1810
rect 20716 1773 20761 1807
rect 20795 1773 20836 1807
rect 20716 1770 20836 1773
rect 22016 1807 22136 1810
rect 22016 1773 22061 1807
rect 22095 1773 22136 1807
rect 22016 1770 22136 1773
rect 23316 1807 23436 1810
rect 23316 1773 23361 1807
rect 23395 1773 23436 1807
rect 23316 1770 23436 1773
rect 24616 1807 24736 1810
rect 24616 1773 24661 1807
rect 24695 1773 24736 1807
rect 24616 1770 24736 1773
rect 25916 1807 26036 1810
rect 25916 1773 25961 1807
rect 25995 1773 26036 1807
rect 25916 1770 26036 1773
rect 158 1723 161 1757
rect 195 1723 198 1757
rect 158 1680 198 1723
<< nsubdiffcont >>
rect 1261 1773 1295 1807
rect 2561 1773 2595 1807
rect 3861 1773 3895 1807
rect 5161 1773 5195 1807
rect 6461 1773 6495 1807
rect 7761 1773 7795 1807
rect 9061 1773 9095 1807
rect 10361 1773 10395 1807
rect 11661 1773 11695 1807
rect 12961 1773 12995 1807
rect 14261 1773 14295 1807
rect 15561 1773 15595 1807
rect 16861 1773 16895 1807
rect 18161 1773 18195 1807
rect 19461 1773 19495 1807
rect 20761 1773 20795 1807
rect 22061 1773 22095 1807
rect 23361 1773 23395 1807
rect 24661 1773 24695 1807
rect 25961 1773 25995 1807
rect 161 1723 195 1757
<< poly >>
rect 311 1645 711 1671
rect 769 1645 1169 1671
rect 1227 1645 1627 1671
rect 1685 1645 2085 1671
rect 2143 1645 2543 1671
rect 2601 1645 3001 1671
rect 3059 1645 3459 1671
rect 3517 1645 3917 1671
rect 3975 1645 4375 1671
rect 4433 1645 4833 1671
rect 4891 1645 5291 1671
rect 5349 1645 5749 1671
rect 5807 1645 6207 1671
rect 6265 1645 6665 1671
rect 6723 1645 7123 1671
rect 7181 1645 7581 1671
rect 7639 1645 8039 1671
rect 8097 1645 8497 1671
rect 8555 1645 8955 1671
rect 9013 1645 9413 1671
rect 9471 1645 9871 1671
rect 9929 1645 10329 1671
rect 10387 1645 10787 1671
rect 10845 1645 11245 1671
rect 11303 1645 11703 1671
rect 11761 1645 12161 1671
rect 12219 1645 12619 1671
rect 12677 1645 13077 1671
rect 13135 1645 13535 1671
rect 13593 1645 13993 1671
rect 14051 1645 14451 1671
rect 14509 1645 14909 1671
rect 14967 1645 15367 1671
rect 15425 1645 15825 1671
rect 15883 1645 16283 1671
rect 16341 1645 16741 1671
rect 16799 1645 17199 1671
rect 17257 1645 17657 1671
rect 17715 1645 18115 1671
rect 18173 1645 18573 1671
rect 18631 1645 19031 1671
rect 19089 1645 19489 1671
rect 19547 1645 19947 1671
rect 20005 1645 20405 1671
rect 20463 1645 20863 1671
rect 20921 1645 21321 1671
rect 21379 1645 21779 1671
rect 21837 1645 22237 1671
rect 22295 1645 22695 1671
rect 22753 1645 23153 1671
rect 23211 1645 23611 1671
rect 23669 1645 24069 1671
rect 24127 1645 24527 1671
rect 24585 1645 24985 1671
rect 25043 1645 25443 1671
rect 25501 1645 25901 1671
rect 25959 1645 26359 1671
rect 26417 1645 26817 1671
rect 26875 1645 27275 1671
rect 27333 1645 27733 1671
rect 311 329 711 355
rect 769 329 1169 355
rect 1227 329 1627 355
rect 1685 329 2085 355
rect 2143 329 2543 355
rect 2601 329 3001 355
rect 3059 329 3459 355
rect 3517 329 3917 355
rect 3975 329 4375 355
rect 4433 329 4833 355
rect 4891 329 5291 355
rect 5349 329 5749 355
rect 5807 329 6207 355
rect 6265 329 6665 355
rect 6723 329 7123 355
rect 7181 329 7581 355
rect 7639 329 8039 355
rect 8097 329 8497 355
rect 8555 329 8955 355
rect 9013 329 9413 355
rect 9471 329 9871 355
rect 9929 329 10329 355
rect 10387 329 10787 355
rect 10845 329 11245 355
rect 11303 329 11703 355
rect 11761 329 12161 355
rect 12219 329 12619 355
rect 12677 329 13077 355
rect 13135 329 13535 355
rect 13593 329 13993 355
rect 14051 329 14451 355
rect 14509 329 14909 355
rect 14967 329 15367 355
rect 15425 329 15825 355
rect 15883 329 16283 355
rect 16341 329 16741 355
rect 16799 329 17199 355
rect 17257 329 17657 355
rect 17715 329 18115 355
rect 18173 329 18573 355
rect 18631 329 19031 355
rect 19089 329 19489 355
rect 19547 329 19947 355
rect 20005 329 20405 355
rect 20463 329 20863 355
rect 20921 329 21321 355
rect 21379 329 21779 355
rect 21837 329 22237 355
rect 22295 329 22695 355
rect 22753 329 23153 355
rect 23211 329 23611 355
rect 23669 329 24069 355
rect 24127 329 24527 355
rect 24585 329 24985 355
rect 25043 329 25443 355
rect 25501 329 25901 355
rect 25959 329 26359 355
rect 26417 329 26817 355
rect 26875 329 27275 355
rect 27333 329 27733 355
rect 458 184 578 329
rect 914 184 1034 329
rect 1370 184 1490 329
rect 1826 184 1946 329
rect 2282 184 2402 329
rect 2738 184 2858 329
rect 3194 184 3314 329
rect 3650 184 3770 329
rect 4106 184 4226 329
rect 4562 184 4682 329
rect 5018 184 5138 329
rect 5474 184 5594 329
rect 5930 184 6050 329
rect 6386 184 6506 329
rect 6842 184 6962 329
rect 7298 184 7418 329
rect 7754 184 7874 329
rect 8210 184 8330 329
rect 8666 184 8786 329
rect 9122 184 9242 329
rect 9578 184 9698 329
rect 10034 184 10154 329
rect 10490 184 10610 329
rect 10946 184 11066 329
rect 11402 184 11522 329
rect 11858 184 11978 329
rect 12314 184 12434 329
rect 12770 184 12890 329
rect 13226 184 13346 329
rect 13682 184 13802 329
rect 14138 184 14258 329
rect 14594 184 14714 329
rect 15050 184 15170 329
rect 15506 184 15626 329
rect 15962 184 16082 329
rect 16418 184 16538 329
rect 16874 184 16994 329
rect 17330 184 17450 329
rect 17786 184 17906 329
rect 18242 184 18362 329
rect 18698 184 18818 329
rect 19154 184 19274 329
rect 19610 184 19730 329
rect 20066 184 20186 329
rect 20522 184 20642 329
rect 20978 184 21098 329
rect 21434 184 21554 329
rect 21890 184 22010 329
rect 22346 184 22466 329
rect 22802 184 22922 329
rect 23258 184 23378 329
rect 23714 184 23834 329
rect 24170 184 24290 329
rect 24626 184 24746 329
rect 25082 184 25202 329
rect 25538 184 25658 329
rect 25994 184 26114 329
rect 26450 184 26570 329
rect 26906 184 27026 329
rect 27362 184 27482 329
rect 218 151 27826 184
rect 218 117 401 151
rect 435 117 801 151
rect 835 117 1201 151
rect 1235 117 1601 151
rect 1635 117 2001 151
rect 2035 117 2401 151
rect 2435 117 2801 151
rect 2835 117 3201 151
rect 3235 117 3601 151
rect 3635 117 4001 151
rect 4035 117 4401 151
rect 4435 117 4801 151
rect 4835 117 5201 151
rect 5235 117 5601 151
rect 5635 117 6001 151
rect 6035 117 6401 151
rect 6435 117 6801 151
rect 6835 117 7201 151
rect 7235 117 7601 151
rect 7635 117 8001 151
rect 8035 117 8401 151
rect 8435 117 8801 151
rect 8835 117 9201 151
rect 9235 117 9601 151
rect 9635 117 10001 151
rect 10035 117 10401 151
rect 10435 117 10801 151
rect 10835 117 11201 151
rect 11235 117 11601 151
rect 11635 117 12001 151
rect 12035 117 12401 151
rect 12435 117 12801 151
rect 12835 117 13201 151
rect 13235 117 13601 151
rect 13635 117 14001 151
rect 14035 117 14401 151
rect 14435 117 14801 151
rect 14835 117 15201 151
rect 15235 117 15601 151
rect 15635 117 16001 151
rect 16035 117 16401 151
rect 16435 117 16801 151
rect 16835 117 17201 151
rect 17235 117 17601 151
rect 17635 117 18001 151
rect 18035 117 18401 151
rect 18435 117 18801 151
rect 18835 117 19201 151
rect 19235 117 19601 151
rect 19635 117 20001 151
rect 20035 117 20401 151
rect 20435 117 20801 151
rect 20835 117 21201 151
rect 21235 117 21601 151
rect 21635 117 22001 151
rect 22035 117 22401 151
rect 22435 117 22801 151
rect 22835 117 23201 151
rect 23235 117 23601 151
rect 23635 117 24001 151
rect 24035 117 24401 151
rect 24435 117 24801 151
rect 24835 117 25201 151
rect 25235 117 25601 151
rect 25635 117 26001 151
rect 26035 117 26401 151
rect 26435 117 26801 151
rect 26835 117 27201 151
rect 27235 117 27601 151
rect 27635 117 27826 151
rect 218 84 27826 117
<< polycont >>
rect 401 117 435 151
rect 801 117 835 151
rect 1201 117 1235 151
rect 1601 117 1635 151
rect 2001 117 2035 151
rect 2401 117 2435 151
rect 2801 117 2835 151
rect 3201 117 3235 151
rect 3601 117 3635 151
rect 4001 117 4035 151
rect 4401 117 4435 151
rect 4801 117 4835 151
rect 5201 117 5235 151
rect 5601 117 5635 151
rect 6001 117 6035 151
rect 6401 117 6435 151
rect 6801 117 6835 151
rect 7201 117 7235 151
rect 7601 117 7635 151
rect 8001 117 8035 151
rect 8401 117 8435 151
rect 8801 117 8835 151
rect 9201 117 9235 151
rect 9601 117 9635 151
rect 10001 117 10035 151
rect 10401 117 10435 151
rect 10801 117 10835 151
rect 11201 117 11235 151
rect 11601 117 11635 151
rect 12001 117 12035 151
rect 12401 117 12435 151
rect 12801 117 12835 151
rect 13201 117 13235 151
rect 13601 117 13635 151
rect 14001 117 14035 151
rect 14401 117 14435 151
rect 14801 117 14835 151
rect 15201 117 15235 151
rect 15601 117 15635 151
rect 16001 117 16035 151
rect 16401 117 16435 151
rect 16801 117 16835 151
rect 17201 117 17235 151
rect 17601 117 17635 151
rect 18001 117 18035 151
rect 18401 117 18435 151
rect 18801 117 18835 151
rect 19201 117 19235 151
rect 19601 117 19635 151
rect 20001 117 20035 151
rect 20401 117 20435 151
rect 20801 117 20835 151
rect 21201 117 21235 151
rect 21601 117 21635 151
rect 22001 117 22035 151
rect 22401 117 22435 151
rect 22801 117 22835 151
rect 23201 117 23235 151
rect 23601 117 23635 151
rect 24001 117 24035 151
rect 24401 117 24435 151
rect 24801 117 24835 151
rect 25201 117 25235 151
rect 25601 117 25635 151
rect 26001 117 26035 151
rect 26401 117 26435 151
rect 26801 117 26835 151
rect 27201 117 27235 151
rect 27601 117 27635 151
<< locali >>
rect 120 1897 27826 1910
rect 120 1863 401 1897
rect 435 1863 801 1897
rect 835 1863 1201 1897
rect 1235 1863 1601 1897
rect 1635 1863 2001 1897
rect 2035 1863 2401 1897
rect 2435 1863 2801 1897
rect 2835 1863 3201 1897
rect 3235 1863 3601 1897
rect 3635 1863 4001 1897
rect 4035 1863 4401 1897
rect 4435 1863 4801 1897
rect 4835 1863 5201 1897
rect 5235 1863 5601 1897
rect 5635 1863 6001 1897
rect 6035 1863 6401 1897
rect 6435 1863 6801 1897
rect 6835 1863 7201 1897
rect 7235 1863 7601 1897
rect 7635 1863 8001 1897
rect 8035 1863 8401 1897
rect 8435 1863 8801 1897
rect 8835 1863 9201 1897
rect 9235 1863 9601 1897
rect 9635 1863 10001 1897
rect 10035 1863 10401 1897
rect 10435 1863 10801 1897
rect 10835 1863 11201 1897
rect 11235 1863 11601 1897
rect 11635 1863 12001 1897
rect 12035 1863 12401 1897
rect 12435 1863 12801 1897
rect 12835 1863 13201 1897
rect 13235 1863 13601 1897
rect 13635 1863 14001 1897
rect 14035 1863 14401 1897
rect 14435 1863 14801 1897
rect 14835 1863 15201 1897
rect 15235 1863 15601 1897
rect 15635 1863 16001 1897
rect 16035 1863 16401 1897
rect 16435 1863 16801 1897
rect 16835 1863 17201 1897
rect 17235 1863 17601 1897
rect 17635 1863 18001 1897
rect 18035 1863 18401 1897
rect 18435 1863 18801 1897
rect 18835 1863 19201 1897
rect 19235 1863 19601 1897
rect 19635 1863 20001 1897
rect 20035 1863 20401 1897
rect 20435 1863 20801 1897
rect 20835 1863 21201 1897
rect 21235 1863 21601 1897
rect 21635 1863 22001 1897
rect 22035 1863 22401 1897
rect 22435 1863 22801 1897
rect 22835 1863 23201 1897
rect 23235 1863 23601 1897
rect 23635 1863 24001 1897
rect 24035 1863 24401 1897
rect 24435 1863 24801 1897
rect 24835 1863 25201 1897
rect 25235 1863 25601 1897
rect 25635 1863 26001 1897
rect 26035 1863 26401 1897
rect 26435 1863 26801 1897
rect 26835 1863 27201 1897
rect 27235 1863 27601 1897
rect 27635 1863 27826 1897
rect 120 1850 27826 1863
rect 148 1757 208 1850
rect 1196 1807 1356 1850
rect 1196 1773 1261 1807
rect 1295 1773 1356 1807
rect 1196 1770 1356 1773
rect 2496 1807 2656 1850
rect 2496 1773 2561 1807
rect 2595 1773 2656 1807
rect 2496 1770 2656 1773
rect 3796 1807 3956 1850
rect 3796 1773 3861 1807
rect 3895 1773 3956 1807
rect 3796 1770 3956 1773
rect 5096 1807 5256 1850
rect 5096 1773 5161 1807
rect 5195 1773 5256 1807
rect 5096 1770 5256 1773
rect 6396 1807 6556 1850
rect 6396 1773 6461 1807
rect 6495 1773 6556 1807
rect 6396 1770 6556 1773
rect 7696 1807 7856 1850
rect 7696 1773 7761 1807
rect 7795 1773 7856 1807
rect 7696 1770 7856 1773
rect 8996 1807 9156 1850
rect 8996 1773 9061 1807
rect 9095 1773 9156 1807
rect 8996 1770 9156 1773
rect 10296 1807 10456 1850
rect 10296 1773 10361 1807
rect 10395 1773 10456 1807
rect 10296 1770 10456 1773
rect 11596 1807 11756 1850
rect 11596 1773 11661 1807
rect 11695 1773 11756 1807
rect 11596 1770 11756 1773
rect 12896 1807 13056 1850
rect 12896 1773 12961 1807
rect 12995 1773 13056 1807
rect 12896 1770 13056 1773
rect 14196 1807 14356 1850
rect 14196 1773 14261 1807
rect 14295 1773 14356 1807
rect 14196 1770 14356 1773
rect 15496 1807 15656 1850
rect 15496 1773 15561 1807
rect 15595 1773 15656 1807
rect 15496 1770 15656 1773
rect 16796 1807 16956 1850
rect 16796 1773 16861 1807
rect 16895 1773 16956 1807
rect 16796 1770 16956 1773
rect 18096 1807 18256 1850
rect 18096 1773 18161 1807
rect 18195 1773 18256 1807
rect 18096 1770 18256 1773
rect 19396 1807 19556 1850
rect 19396 1773 19461 1807
rect 19495 1773 19556 1807
rect 19396 1770 19556 1773
rect 20696 1807 20856 1850
rect 20696 1773 20761 1807
rect 20795 1773 20856 1807
rect 20696 1770 20856 1773
rect 21996 1807 22156 1850
rect 21996 1773 22061 1807
rect 22095 1773 22156 1807
rect 21996 1770 22156 1773
rect 23296 1807 23456 1850
rect 23296 1773 23361 1807
rect 23395 1773 23456 1807
rect 23296 1770 23456 1773
rect 24596 1807 24756 1850
rect 24596 1773 24661 1807
rect 24695 1773 24756 1807
rect 24596 1770 24756 1773
rect 25896 1807 26056 1850
rect 25896 1773 25961 1807
rect 25995 1773 26056 1807
rect 25896 1770 26056 1773
rect 148 1723 161 1757
rect 195 1723 208 1757
rect 148 1640 208 1723
rect 278 1690 27826 1730
rect 265 1629 299 1649
rect 265 1561 299 1595
rect 265 1493 299 1523
rect 265 1425 299 1451
rect 265 1357 299 1379
rect 265 1289 299 1307
rect 265 1221 299 1235
rect 265 1153 299 1163
rect 265 1085 299 1091
rect 265 1017 299 1019
rect 265 981 299 983
rect 265 909 299 915
rect 265 837 299 847
rect 265 765 299 779
rect 265 693 299 711
rect 265 621 299 643
rect 265 549 299 575
rect 265 477 299 507
rect 265 405 299 439
rect 265 270 299 371
rect 723 1629 757 1690
rect 723 1561 757 1595
rect 723 1493 757 1523
rect 723 1425 757 1451
rect 723 1357 757 1379
rect 723 1289 757 1307
rect 723 1221 757 1235
rect 723 1153 757 1163
rect 723 1085 757 1091
rect 723 1017 757 1019
rect 723 981 757 983
rect 723 909 757 915
rect 723 837 757 847
rect 723 765 757 779
rect 723 693 757 711
rect 723 621 757 643
rect 723 549 757 575
rect 723 477 757 507
rect 723 405 757 439
rect 723 351 757 371
rect 1181 1629 1215 1649
rect 1181 1561 1215 1595
rect 1181 1493 1215 1523
rect 1181 1425 1215 1451
rect 1181 1357 1215 1379
rect 1181 1289 1215 1307
rect 1181 1221 1215 1235
rect 1181 1153 1215 1163
rect 1181 1085 1215 1091
rect 1181 1017 1215 1019
rect 1181 981 1215 983
rect 1181 909 1215 915
rect 1181 837 1215 847
rect 1181 765 1215 779
rect 1181 693 1215 711
rect 1181 621 1215 643
rect 1181 549 1215 575
rect 1181 477 1215 507
rect 1181 405 1215 439
rect 1181 270 1215 371
rect 1639 1629 1673 1690
rect 1639 1561 1673 1595
rect 1639 1493 1673 1523
rect 1639 1425 1673 1451
rect 1639 1357 1673 1379
rect 1639 1289 1673 1307
rect 1639 1221 1673 1235
rect 1639 1153 1673 1163
rect 1639 1085 1673 1091
rect 1639 1017 1673 1019
rect 1639 981 1673 983
rect 1639 909 1673 915
rect 1639 837 1673 847
rect 1639 765 1673 779
rect 1639 693 1673 711
rect 1639 621 1673 643
rect 1639 549 1673 575
rect 1639 477 1673 507
rect 1639 405 1673 439
rect 1639 351 1673 371
rect 2097 1629 2131 1649
rect 2097 1561 2131 1595
rect 2097 1493 2131 1523
rect 2097 1425 2131 1451
rect 2097 1357 2131 1379
rect 2097 1289 2131 1307
rect 2097 1221 2131 1235
rect 2097 1153 2131 1163
rect 2097 1085 2131 1091
rect 2097 1017 2131 1019
rect 2097 981 2131 983
rect 2097 909 2131 915
rect 2097 837 2131 847
rect 2097 765 2131 779
rect 2097 693 2131 711
rect 2097 621 2131 643
rect 2097 549 2131 575
rect 2097 477 2131 507
rect 2097 405 2131 439
rect 2097 270 2131 371
rect 2555 1629 2589 1690
rect 2555 1561 2589 1595
rect 2555 1493 2589 1523
rect 2555 1425 2589 1451
rect 2555 1357 2589 1379
rect 2555 1289 2589 1307
rect 2555 1221 2589 1235
rect 2555 1153 2589 1163
rect 2555 1085 2589 1091
rect 2555 1017 2589 1019
rect 2555 981 2589 983
rect 2555 909 2589 915
rect 2555 837 2589 847
rect 2555 765 2589 779
rect 2555 693 2589 711
rect 2555 621 2589 643
rect 2555 549 2589 575
rect 2555 477 2589 507
rect 2555 405 2589 439
rect 2555 351 2589 371
rect 3013 1629 3047 1649
rect 3013 1561 3047 1595
rect 3013 1493 3047 1523
rect 3013 1425 3047 1451
rect 3013 1357 3047 1379
rect 3013 1289 3047 1307
rect 3013 1221 3047 1235
rect 3013 1153 3047 1163
rect 3013 1085 3047 1091
rect 3013 1017 3047 1019
rect 3013 981 3047 983
rect 3013 909 3047 915
rect 3013 837 3047 847
rect 3013 765 3047 779
rect 3013 693 3047 711
rect 3013 621 3047 643
rect 3013 549 3047 575
rect 3013 477 3047 507
rect 3013 405 3047 439
rect 3013 270 3047 371
rect 3471 1629 3505 1690
rect 3471 1561 3505 1595
rect 3471 1493 3505 1523
rect 3471 1425 3505 1451
rect 3471 1357 3505 1379
rect 3471 1289 3505 1307
rect 3471 1221 3505 1235
rect 3471 1153 3505 1163
rect 3471 1085 3505 1091
rect 3471 1017 3505 1019
rect 3471 981 3505 983
rect 3471 909 3505 915
rect 3471 837 3505 847
rect 3471 765 3505 779
rect 3471 693 3505 711
rect 3471 621 3505 643
rect 3471 549 3505 575
rect 3471 477 3505 507
rect 3471 405 3505 439
rect 3471 351 3505 371
rect 3929 1629 3963 1649
rect 3929 1561 3963 1595
rect 3929 1493 3963 1523
rect 3929 1425 3963 1451
rect 3929 1357 3963 1379
rect 3929 1289 3963 1307
rect 3929 1221 3963 1235
rect 3929 1153 3963 1163
rect 3929 1085 3963 1091
rect 3929 1017 3963 1019
rect 3929 981 3963 983
rect 3929 909 3963 915
rect 3929 837 3963 847
rect 3929 765 3963 779
rect 3929 693 3963 711
rect 3929 621 3963 643
rect 3929 549 3963 575
rect 3929 477 3963 507
rect 3929 405 3963 439
rect 3929 270 3963 371
rect 4387 1629 4421 1690
rect 4387 1561 4421 1595
rect 4387 1493 4421 1523
rect 4387 1425 4421 1451
rect 4387 1357 4421 1379
rect 4387 1289 4421 1307
rect 4387 1221 4421 1235
rect 4387 1153 4421 1163
rect 4387 1085 4421 1091
rect 4387 1017 4421 1019
rect 4387 981 4421 983
rect 4387 909 4421 915
rect 4387 837 4421 847
rect 4387 765 4421 779
rect 4387 693 4421 711
rect 4387 621 4421 643
rect 4387 549 4421 575
rect 4387 477 4421 507
rect 4387 405 4421 439
rect 4387 351 4421 371
rect 4845 1629 4879 1649
rect 4845 1561 4879 1595
rect 4845 1493 4879 1523
rect 4845 1425 4879 1451
rect 4845 1357 4879 1379
rect 4845 1289 4879 1307
rect 4845 1221 4879 1235
rect 4845 1153 4879 1163
rect 4845 1085 4879 1091
rect 4845 1017 4879 1019
rect 4845 981 4879 983
rect 4845 909 4879 915
rect 4845 837 4879 847
rect 4845 765 4879 779
rect 4845 693 4879 711
rect 4845 621 4879 643
rect 4845 549 4879 575
rect 4845 477 4879 507
rect 4845 405 4879 439
rect 4845 270 4879 371
rect 5303 1629 5337 1690
rect 5303 1561 5337 1595
rect 5303 1493 5337 1523
rect 5303 1425 5337 1451
rect 5303 1357 5337 1379
rect 5303 1289 5337 1307
rect 5303 1221 5337 1235
rect 5303 1153 5337 1163
rect 5303 1085 5337 1091
rect 5303 1017 5337 1019
rect 5303 981 5337 983
rect 5303 909 5337 915
rect 5303 837 5337 847
rect 5303 765 5337 779
rect 5303 693 5337 711
rect 5303 621 5337 643
rect 5303 549 5337 575
rect 5303 477 5337 507
rect 5303 405 5337 439
rect 5303 351 5337 371
rect 5761 1629 5795 1649
rect 5761 1561 5795 1595
rect 5761 1493 5795 1523
rect 5761 1425 5795 1451
rect 5761 1357 5795 1379
rect 5761 1289 5795 1307
rect 5761 1221 5795 1235
rect 5761 1153 5795 1163
rect 5761 1085 5795 1091
rect 5761 1017 5795 1019
rect 5761 981 5795 983
rect 5761 909 5795 915
rect 5761 837 5795 847
rect 5761 765 5795 779
rect 5761 693 5795 711
rect 5761 621 5795 643
rect 5761 549 5795 575
rect 5761 477 5795 507
rect 5761 405 5795 439
rect 5761 270 5795 371
rect 6219 1629 6253 1690
rect 6219 1561 6253 1595
rect 6219 1493 6253 1523
rect 6219 1425 6253 1451
rect 6219 1357 6253 1379
rect 6219 1289 6253 1307
rect 6219 1221 6253 1235
rect 6219 1153 6253 1163
rect 6219 1085 6253 1091
rect 6219 1017 6253 1019
rect 6219 981 6253 983
rect 6219 909 6253 915
rect 6219 837 6253 847
rect 6219 765 6253 779
rect 6219 693 6253 711
rect 6219 621 6253 643
rect 6219 549 6253 575
rect 6219 477 6253 507
rect 6219 405 6253 439
rect 6219 351 6253 371
rect 6677 1629 6711 1649
rect 6677 1561 6711 1595
rect 6677 1493 6711 1523
rect 6677 1425 6711 1451
rect 6677 1357 6711 1379
rect 6677 1289 6711 1307
rect 6677 1221 6711 1235
rect 6677 1153 6711 1163
rect 6677 1085 6711 1091
rect 6677 1017 6711 1019
rect 6677 981 6711 983
rect 6677 909 6711 915
rect 6677 837 6711 847
rect 6677 765 6711 779
rect 6677 693 6711 711
rect 6677 621 6711 643
rect 6677 549 6711 575
rect 6677 477 6711 507
rect 6677 405 6711 439
rect 6677 270 6711 371
rect 7135 1629 7169 1690
rect 7135 1561 7169 1595
rect 7135 1493 7169 1523
rect 7135 1425 7169 1451
rect 7135 1357 7169 1379
rect 7135 1289 7169 1307
rect 7135 1221 7169 1235
rect 7135 1153 7169 1163
rect 7135 1085 7169 1091
rect 7135 1017 7169 1019
rect 7135 981 7169 983
rect 7135 909 7169 915
rect 7135 837 7169 847
rect 7135 765 7169 779
rect 7135 693 7169 711
rect 7135 621 7169 643
rect 7135 549 7169 575
rect 7135 477 7169 507
rect 7135 405 7169 439
rect 7135 351 7169 371
rect 7593 1629 7627 1649
rect 7593 1561 7627 1595
rect 7593 1493 7627 1523
rect 7593 1425 7627 1451
rect 7593 1357 7627 1379
rect 7593 1289 7627 1307
rect 7593 1221 7627 1235
rect 7593 1153 7627 1163
rect 7593 1085 7627 1091
rect 7593 1017 7627 1019
rect 7593 981 7627 983
rect 7593 909 7627 915
rect 7593 837 7627 847
rect 7593 765 7627 779
rect 7593 693 7627 711
rect 7593 621 7627 643
rect 7593 549 7627 575
rect 7593 477 7627 507
rect 7593 405 7627 439
rect 7593 270 7627 371
rect 8051 1629 8085 1690
rect 8051 1561 8085 1595
rect 8051 1493 8085 1523
rect 8051 1425 8085 1451
rect 8051 1357 8085 1379
rect 8051 1289 8085 1307
rect 8051 1221 8085 1235
rect 8051 1153 8085 1163
rect 8051 1085 8085 1091
rect 8051 1017 8085 1019
rect 8051 981 8085 983
rect 8051 909 8085 915
rect 8051 837 8085 847
rect 8051 765 8085 779
rect 8051 693 8085 711
rect 8051 621 8085 643
rect 8051 549 8085 575
rect 8051 477 8085 507
rect 8051 405 8085 439
rect 8051 351 8085 371
rect 8509 1629 8543 1649
rect 8509 1561 8543 1595
rect 8509 1493 8543 1523
rect 8509 1425 8543 1451
rect 8509 1357 8543 1379
rect 8509 1289 8543 1307
rect 8509 1221 8543 1235
rect 8509 1153 8543 1163
rect 8509 1085 8543 1091
rect 8509 1017 8543 1019
rect 8509 981 8543 983
rect 8509 909 8543 915
rect 8509 837 8543 847
rect 8509 765 8543 779
rect 8509 693 8543 711
rect 8509 621 8543 643
rect 8509 549 8543 575
rect 8509 477 8543 507
rect 8509 405 8543 439
rect 8509 270 8543 371
rect 8967 1629 9001 1690
rect 8967 1561 9001 1595
rect 8967 1493 9001 1523
rect 8967 1425 9001 1451
rect 8967 1357 9001 1379
rect 8967 1289 9001 1307
rect 8967 1221 9001 1235
rect 8967 1153 9001 1163
rect 8967 1085 9001 1091
rect 8967 1017 9001 1019
rect 8967 981 9001 983
rect 8967 909 9001 915
rect 8967 837 9001 847
rect 8967 765 9001 779
rect 8967 693 9001 711
rect 8967 621 9001 643
rect 8967 549 9001 575
rect 8967 477 9001 507
rect 8967 405 9001 439
rect 8967 351 9001 371
rect 9425 1629 9459 1649
rect 9425 1561 9459 1595
rect 9425 1493 9459 1523
rect 9425 1425 9459 1451
rect 9425 1357 9459 1379
rect 9425 1289 9459 1307
rect 9425 1221 9459 1235
rect 9425 1153 9459 1163
rect 9425 1085 9459 1091
rect 9425 1017 9459 1019
rect 9425 981 9459 983
rect 9425 909 9459 915
rect 9425 837 9459 847
rect 9425 765 9459 779
rect 9425 693 9459 711
rect 9425 621 9459 643
rect 9425 549 9459 575
rect 9425 477 9459 507
rect 9425 405 9459 439
rect 9425 270 9459 371
rect 9883 1629 9917 1690
rect 9883 1561 9917 1595
rect 9883 1493 9917 1523
rect 9883 1425 9917 1451
rect 9883 1357 9917 1379
rect 9883 1289 9917 1307
rect 9883 1221 9917 1235
rect 9883 1153 9917 1163
rect 9883 1085 9917 1091
rect 9883 1017 9917 1019
rect 9883 981 9917 983
rect 9883 909 9917 915
rect 9883 837 9917 847
rect 9883 765 9917 779
rect 9883 693 9917 711
rect 9883 621 9917 643
rect 9883 549 9917 575
rect 9883 477 9917 507
rect 9883 405 9917 439
rect 9883 351 9917 371
rect 10341 1629 10375 1649
rect 10341 1561 10375 1595
rect 10341 1493 10375 1523
rect 10341 1425 10375 1451
rect 10341 1357 10375 1379
rect 10341 1289 10375 1307
rect 10341 1221 10375 1235
rect 10341 1153 10375 1163
rect 10341 1085 10375 1091
rect 10341 1017 10375 1019
rect 10341 981 10375 983
rect 10341 909 10375 915
rect 10341 837 10375 847
rect 10341 765 10375 779
rect 10341 693 10375 711
rect 10341 621 10375 643
rect 10341 549 10375 575
rect 10341 477 10375 507
rect 10341 405 10375 439
rect 10341 270 10375 371
rect 10799 1629 10833 1690
rect 10799 1561 10833 1595
rect 10799 1493 10833 1523
rect 10799 1425 10833 1451
rect 10799 1357 10833 1379
rect 10799 1289 10833 1307
rect 10799 1221 10833 1235
rect 10799 1153 10833 1163
rect 10799 1085 10833 1091
rect 10799 1017 10833 1019
rect 10799 981 10833 983
rect 10799 909 10833 915
rect 10799 837 10833 847
rect 10799 765 10833 779
rect 10799 693 10833 711
rect 10799 621 10833 643
rect 10799 549 10833 575
rect 10799 477 10833 507
rect 10799 405 10833 439
rect 10799 351 10833 371
rect 11257 1629 11291 1649
rect 11257 1561 11291 1595
rect 11257 1493 11291 1523
rect 11257 1425 11291 1451
rect 11257 1357 11291 1379
rect 11257 1289 11291 1307
rect 11257 1221 11291 1235
rect 11257 1153 11291 1163
rect 11257 1085 11291 1091
rect 11257 1017 11291 1019
rect 11257 981 11291 983
rect 11257 909 11291 915
rect 11257 837 11291 847
rect 11257 765 11291 779
rect 11257 693 11291 711
rect 11257 621 11291 643
rect 11257 549 11291 575
rect 11257 477 11291 507
rect 11257 405 11291 439
rect 11257 270 11291 371
rect 11715 1629 11749 1690
rect 11715 1561 11749 1595
rect 11715 1493 11749 1523
rect 11715 1425 11749 1451
rect 11715 1357 11749 1379
rect 11715 1289 11749 1307
rect 11715 1221 11749 1235
rect 11715 1153 11749 1163
rect 11715 1085 11749 1091
rect 11715 1017 11749 1019
rect 11715 981 11749 983
rect 11715 909 11749 915
rect 11715 837 11749 847
rect 11715 765 11749 779
rect 11715 693 11749 711
rect 11715 621 11749 643
rect 11715 549 11749 575
rect 11715 477 11749 507
rect 11715 405 11749 439
rect 11715 351 11749 371
rect 12173 1629 12207 1649
rect 12173 1561 12207 1595
rect 12173 1493 12207 1523
rect 12173 1425 12207 1451
rect 12173 1357 12207 1379
rect 12173 1289 12207 1307
rect 12173 1221 12207 1235
rect 12173 1153 12207 1163
rect 12173 1085 12207 1091
rect 12173 1017 12207 1019
rect 12173 981 12207 983
rect 12173 909 12207 915
rect 12173 837 12207 847
rect 12173 765 12207 779
rect 12173 693 12207 711
rect 12173 621 12207 643
rect 12173 549 12207 575
rect 12173 477 12207 507
rect 12173 405 12207 439
rect 12173 270 12207 371
rect 12631 1629 12665 1690
rect 12631 1561 12665 1595
rect 12631 1493 12665 1523
rect 12631 1425 12665 1451
rect 12631 1357 12665 1379
rect 12631 1289 12665 1307
rect 12631 1221 12665 1235
rect 12631 1153 12665 1163
rect 12631 1085 12665 1091
rect 12631 1017 12665 1019
rect 12631 981 12665 983
rect 12631 909 12665 915
rect 12631 837 12665 847
rect 12631 765 12665 779
rect 12631 693 12665 711
rect 12631 621 12665 643
rect 12631 549 12665 575
rect 12631 477 12665 507
rect 12631 405 12665 439
rect 12631 351 12665 371
rect 13089 1629 13123 1649
rect 13089 1561 13123 1595
rect 13089 1493 13123 1523
rect 13089 1425 13123 1451
rect 13089 1357 13123 1379
rect 13089 1289 13123 1307
rect 13089 1221 13123 1235
rect 13089 1153 13123 1163
rect 13089 1085 13123 1091
rect 13089 1017 13123 1019
rect 13089 981 13123 983
rect 13089 909 13123 915
rect 13089 837 13123 847
rect 13089 765 13123 779
rect 13089 693 13123 711
rect 13089 621 13123 643
rect 13089 549 13123 575
rect 13089 477 13123 507
rect 13089 405 13123 439
rect 13089 270 13123 371
rect 13547 1629 13581 1690
rect 13547 1561 13581 1595
rect 13547 1493 13581 1523
rect 13547 1425 13581 1451
rect 13547 1357 13581 1379
rect 13547 1289 13581 1307
rect 13547 1221 13581 1235
rect 13547 1153 13581 1163
rect 13547 1085 13581 1091
rect 13547 1017 13581 1019
rect 13547 981 13581 983
rect 13547 909 13581 915
rect 13547 837 13581 847
rect 13547 765 13581 779
rect 13547 693 13581 711
rect 13547 621 13581 643
rect 13547 549 13581 575
rect 13547 477 13581 507
rect 13547 405 13581 439
rect 13547 351 13581 371
rect 14005 1629 14039 1649
rect 14005 1561 14039 1595
rect 14005 1493 14039 1523
rect 14005 1425 14039 1451
rect 14005 1357 14039 1379
rect 14005 1289 14039 1307
rect 14005 1221 14039 1235
rect 14005 1153 14039 1163
rect 14005 1085 14039 1091
rect 14005 1017 14039 1019
rect 14005 981 14039 983
rect 14005 909 14039 915
rect 14005 837 14039 847
rect 14005 765 14039 779
rect 14005 693 14039 711
rect 14005 621 14039 643
rect 14005 549 14039 575
rect 14005 477 14039 507
rect 14005 405 14039 439
rect 14005 270 14039 371
rect 14463 1629 14497 1690
rect 14463 1561 14497 1595
rect 14463 1493 14497 1523
rect 14463 1425 14497 1451
rect 14463 1357 14497 1379
rect 14463 1289 14497 1307
rect 14463 1221 14497 1235
rect 14463 1153 14497 1163
rect 14463 1085 14497 1091
rect 14463 1017 14497 1019
rect 14463 981 14497 983
rect 14463 909 14497 915
rect 14463 837 14497 847
rect 14463 765 14497 779
rect 14463 693 14497 711
rect 14463 621 14497 643
rect 14463 549 14497 575
rect 14463 477 14497 507
rect 14463 405 14497 439
rect 14463 351 14497 371
rect 14921 1629 14955 1649
rect 14921 1561 14955 1595
rect 14921 1493 14955 1523
rect 14921 1425 14955 1451
rect 14921 1357 14955 1379
rect 14921 1289 14955 1307
rect 14921 1221 14955 1235
rect 14921 1153 14955 1163
rect 14921 1085 14955 1091
rect 14921 1017 14955 1019
rect 14921 981 14955 983
rect 14921 909 14955 915
rect 14921 837 14955 847
rect 14921 765 14955 779
rect 14921 693 14955 711
rect 14921 621 14955 643
rect 14921 549 14955 575
rect 14921 477 14955 507
rect 14921 405 14955 439
rect 14921 270 14955 371
rect 15379 1629 15413 1690
rect 15379 1561 15413 1595
rect 15379 1493 15413 1523
rect 15379 1425 15413 1451
rect 15379 1357 15413 1379
rect 15379 1289 15413 1307
rect 15379 1221 15413 1235
rect 15379 1153 15413 1163
rect 15379 1085 15413 1091
rect 15379 1017 15413 1019
rect 15379 981 15413 983
rect 15379 909 15413 915
rect 15379 837 15413 847
rect 15379 765 15413 779
rect 15379 693 15413 711
rect 15379 621 15413 643
rect 15379 549 15413 575
rect 15379 477 15413 507
rect 15379 405 15413 439
rect 15379 351 15413 371
rect 15837 1629 15871 1649
rect 15837 1561 15871 1595
rect 15837 1493 15871 1523
rect 15837 1425 15871 1451
rect 15837 1357 15871 1379
rect 15837 1289 15871 1307
rect 15837 1221 15871 1235
rect 15837 1153 15871 1163
rect 15837 1085 15871 1091
rect 15837 1017 15871 1019
rect 15837 981 15871 983
rect 15837 909 15871 915
rect 15837 837 15871 847
rect 15837 765 15871 779
rect 15837 693 15871 711
rect 15837 621 15871 643
rect 15837 549 15871 575
rect 15837 477 15871 507
rect 15837 405 15871 439
rect 15837 270 15871 371
rect 16295 1629 16329 1690
rect 16295 1561 16329 1595
rect 16295 1493 16329 1523
rect 16295 1425 16329 1451
rect 16295 1357 16329 1379
rect 16295 1289 16329 1307
rect 16295 1221 16329 1235
rect 16295 1153 16329 1163
rect 16295 1085 16329 1091
rect 16295 1017 16329 1019
rect 16295 981 16329 983
rect 16295 909 16329 915
rect 16295 837 16329 847
rect 16295 765 16329 779
rect 16295 693 16329 711
rect 16295 621 16329 643
rect 16295 549 16329 575
rect 16295 477 16329 507
rect 16295 405 16329 439
rect 16295 351 16329 371
rect 16753 1629 16787 1649
rect 16753 1561 16787 1595
rect 16753 1493 16787 1523
rect 16753 1425 16787 1451
rect 16753 1357 16787 1379
rect 16753 1289 16787 1307
rect 16753 1221 16787 1235
rect 16753 1153 16787 1163
rect 16753 1085 16787 1091
rect 16753 1017 16787 1019
rect 16753 981 16787 983
rect 16753 909 16787 915
rect 16753 837 16787 847
rect 16753 765 16787 779
rect 16753 693 16787 711
rect 16753 621 16787 643
rect 16753 549 16787 575
rect 16753 477 16787 507
rect 16753 405 16787 439
rect 16753 270 16787 371
rect 17211 1629 17245 1690
rect 17211 1561 17245 1595
rect 17211 1493 17245 1523
rect 17211 1425 17245 1451
rect 17211 1357 17245 1379
rect 17211 1289 17245 1307
rect 17211 1221 17245 1235
rect 17211 1153 17245 1163
rect 17211 1085 17245 1091
rect 17211 1017 17245 1019
rect 17211 981 17245 983
rect 17211 909 17245 915
rect 17211 837 17245 847
rect 17211 765 17245 779
rect 17211 693 17245 711
rect 17211 621 17245 643
rect 17211 549 17245 575
rect 17211 477 17245 507
rect 17211 405 17245 439
rect 17211 351 17245 371
rect 17669 1629 17703 1649
rect 17669 1561 17703 1595
rect 17669 1493 17703 1523
rect 17669 1425 17703 1451
rect 17669 1357 17703 1379
rect 17669 1289 17703 1307
rect 17669 1221 17703 1235
rect 17669 1153 17703 1163
rect 17669 1085 17703 1091
rect 17669 1017 17703 1019
rect 17669 981 17703 983
rect 17669 909 17703 915
rect 17669 837 17703 847
rect 17669 765 17703 779
rect 17669 693 17703 711
rect 17669 621 17703 643
rect 17669 549 17703 575
rect 17669 477 17703 507
rect 17669 405 17703 439
rect 17669 270 17703 371
rect 18127 1629 18161 1690
rect 18127 1561 18161 1595
rect 18127 1493 18161 1523
rect 18127 1425 18161 1451
rect 18127 1357 18161 1379
rect 18127 1289 18161 1307
rect 18127 1221 18161 1235
rect 18127 1153 18161 1163
rect 18127 1085 18161 1091
rect 18127 1017 18161 1019
rect 18127 981 18161 983
rect 18127 909 18161 915
rect 18127 837 18161 847
rect 18127 765 18161 779
rect 18127 693 18161 711
rect 18127 621 18161 643
rect 18127 549 18161 575
rect 18127 477 18161 507
rect 18127 405 18161 439
rect 18127 351 18161 371
rect 18585 1629 18619 1649
rect 18585 1561 18619 1595
rect 18585 1493 18619 1523
rect 18585 1425 18619 1451
rect 18585 1357 18619 1379
rect 18585 1289 18619 1307
rect 18585 1221 18619 1235
rect 18585 1153 18619 1163
rect 18585 1085 18619 1091
rect 18585 1017 18619 1019
rect 18585 981 18619 983
rect 18585 909 18619 915
rect 18585 837 18619 847
rect 18585 765 18619 779
rect 18585 693 18619 711
rect 18585 621 18619 643
rect 18585 549 18619 575
rect 18585 477 18619 507
rect 18585 405 18619 439
rect 18585 270 18619 371
rect 19043 1629 19077 1690
rect 19043 1561 19077 1595
rect 19043 1493 19077 1523
rect 19043 1425 19077 1451
rect 19043 1357 19077 1379
rect 19043 1289 19077 1307
rect 19043 1221 19077 1235
rect 19043 1153 19077 1163
rect 19043 1085 19077 1091
rect 19043 1017 19077 1019
rect 19043 981 19077 983
rect 19043 909 19077 915
rect 19043 837 19077 847
rect 19043 765 19077 779
rect 19043 693 19077 711
rect 19043 621 19077 643
rect 19043 549 19077 575
rect 19043 477 19077 507
rect 19043 405 19077 439
rect 19043 351 19077 371
rect 19501 1629 19535 1649
rect 19501 1561 19535 1595
rect 19501 1493 19535 1523
rect 19501 1425 19535 1451
rect 19501 1357 19535 1379
rect 19501 1289 19535 1307
rect 19501 1221 19535 1235
rect 19501 1153 19535 1163
rect 19501 1085 19535 1091
rect 19501 1017 19535 1019
rect 19501 981 19535 983
rect 19501 909 19535 915
rect 19501 837 19535 847
rect 19501 765 19535 779
rect 19501 693 19535 711
rect 19501 621 19535 643
rect 19501 549 19535 575
rect 19501 477 19535 507
rect 19501 405 19535 439
rect 19501 270 19535 371
rect 19959 1629 19993 1690
rect 19959 1561 19993 1595
rect 19959 1493 19993 1523
rect 19959 1425 19993 1451
rect 19959 1357 19993 1379
rect 19959 1289 19993 1307
rect 19959 1221 19993 1235
rect 19959 1153 19993 1163
rect 19959 1085 19993 1091
rect 19959 1017 19993 1019
rect 19959 981 19993 983
rect 19959 909 19993 915
rect 19959 837 19993 847
rect 19959 765 19993 779
rect 19959 693 19993 711
rect 19959 621 19993 643
rect 19959 549 19993 575
rect 19959 477 19993 507
rect 19959 405 19993 439
rect 19959 351 19993 371
rect 20417 1629 20451 1649
rect 20417 1561 20451 1595
rect 20417 1493 20451 1523
rect 20417 1425 20451 1451
rect 20417 1357 20451 1379
rect 20417 1289 20451 1307
rect 20417 1221 20451 1235
rect 20417 1153 20451 1163
rect 20417 1085 20451 1091
rect 20417 1017 20451 1019
rect 20417 981 20451 983
rect 20417 909 20451 915
rect 20417 837 20451 847
rect 20417 765 20451 779
rect 20417 693 20451 711
rect 20417 621 20451 643
rect 20417 549 20451 575
rect 20417 477 20451 507
rect 20417 405 20451 439
rect 20417 270 20451 371
rect 20875 1629 20909 1690
rect 20875 1561 20909 1595
rect 20875 1493 20909 1523
rect 20875 1425 20909 1451
rect 20875 1357 20909 1379
rect 20875 1289 20909 1307
rect 20875 1221 20909 1235
rect 20875 1153 20909 1163
rect 20875 1085 20909 1091
rect 20875 1017 20909 1019
rect 20875 981 20909 983
rect 20875 909 20909 915
rect 20875 837 20909 847
rect 20875 765 20909 779
rect 20875 693 20909 711
rect 20875 621 20909 643
rect 20875 549 20909 575
rect 20875 477 20909 507
rect 20875 405 20909 439
rect 20875 351 20909 371
rect 21333 1629 21367 1649
rect 21333 1561 21367 1595
rect 21333 1493 21367 1523
rect 21333 1425 21367 1451
rect 21333 1357 21367 1379
rect 21333 1289 21367 1307
rect 21333 1221 21367 1235
rect 21333 1153 21367 1163
rect 21333 1085 21367 1091
rect 21333 1017 21367 1019
rect 21333 981 21367 983
rect 21333 909 21367 915
rect 21333 837 21367 847
rect 21333 765 21367 779
rect 21333 693 21367 711
rect 21333 621 21367 643
rect 21333 549 21367 575
rect 21333 477 21367 507
rect 21333 405 21367 439
rect 21333 270 21367 371
rect 21791 1629 21825 1690
rect 21791 1561 21825 1595
rect 21791 1493 21825 1523
rect 21791 1425 21825 1451
rect 21791 1357 21825 1379
rect 21791 1289 21825 1307
rect 21791 1221 21825 1235
rect 21791 1153 21825 1163
rect 21791 1085 21825 1091
rect 21791 1017 21825 1019
rect 21791 981 21825 983
rect 21791 909 21825 915
rect 21791 837 21825 847
rect 21791 765 21825 779
rect 21791 693 21825 711
rect 21791 621 21825 643
rect 21791 549 21825 575
rect 21791 477 21825 507
rect 21791 405 21825 439
rect 21791 351 21825 371
rect 22249 1629 22283 1649
rect 22249 1561 22283 1595
rect 22249 1493 22283 1523
rect 22249 1425 22283 1451
rect 22249 1357 22283 1379
rect 22249 1289 22283 1307
rect 22249 1221 22283 1235
rect 22249 1153 22283 1163
rect 22249 1085 22283 1091
rect 22249 1017 22283 1019
rect 22249 981 22283 983
rect 22249 909 22283 915
rect 22249 837 22283 847
rect 22249 765 22283 779
rect 22249 693 22283 711
rect 22249 621 22283 643
rect 22249 549 22283 575
rect 22249 477 22283 507
rect 22249 405 22283 439
rect 22249 270 22283 371
rect 22707 1629 22741 1690
rect 22707 1561 22741 1595
rect 22707 1493 22741 1523
rect 22707 1425 22741 1451
rect 22707 1357 22741 1379
rect 22707 1289 22741 1307
rect 22707 1221 22741 1235
rect 22707 1153 22741 1163
rect 22707 1085 22741 1091
rect 22707 1017 22741 1019
rect 22707 981 22741 983
rect 22707 909 22741 915
rect 22707 837 22741 847
rect 22707 765 22741 779
rect 22707 693 22741 711
rect 22707 621 22741 643
rect 22707 549 22741 575
rect 22707 477 22741 507
rect 22707 405 22741 439
rect 22707 351 22741 371
rect 23165 1629 23199 1649
rect 23165 1561 23199 1595
rect 23165 1493 23199 1523
rect 23165 1425 23199 1451
rect 23165 1357 23199 1379
rect 23165 1289 23199 1307
rect 23165 1221 23199 1235
rect 23165 1153 23199 1163
rect 23165 1085 23199 1091
rect 23165 1017 23199 1019
rect 23165 981 23199 983
rect 23165 909 23199 915
rect 23165 837 23199 847
rect 23165 765 23199 779
rect 23165 693 23199 711
rect 23165 621 23199 643
rect 23165 549 23199 575
rect 23165 477 23199 507
rect 23165 405 23199 439
rect 23165 270 23199 371
rect 23623 1629 23657 1690
rect 23623 1561 23657 1595
rect 23623 1493 23657 1523
rect 23623 1425 23657 1451
rect 23623 1357 23657 1379
rect 23623 1289 23657 1307
rect 23623 1221 23657 1235
rect 23623 1153 23657 1163
rect 23623 1085 23657 1091
rect 23623 1017 23657 1019
rect 23623 981 23657 983
rect 23623 909 23657 915
rect 23623 837 23657 847
rect 23623 765 23657 779
rect 23623 693 23657 711
rect 23623 621 23657 643
rect 23623 549 23657 575
rect 23623 477 23657 507
rect 23623 405 23657 439
rect 23623 351 23657 371
rect 24081 1629 24115 1649
rect 24081 1561 24115 1595
rect 24081 1493 24115 1523
rect 24081 1425 24115 1451
rect 24081 1357 24115 1379
rect 24081 1289 24115 1307
rect 24081 1221 24115 1235
rect 24081 1153 24115 1163
rect 24081 1085 24115 1091
rect 24081 1017 24115 1019
rect 24081 981 24115 983
rect 24081 909 24115 915
rect 24081 837 24115 847
rect 24081 765 24115 779
rect 24081 693 24115 711
rect 24081 621 24115 643
rect 24081 549 24115 575
rect 24081 477 24115 507
rect 24081 405 24115 439
rect 24081 270 24115 371
rect 24539 1629 24573 1690
rect 24539 1561 24573 1595
rect 24539 1493 24573 1523
rect 24539 1425 24573 1451
rect 24539 1357 24573 1379
rect 24539 1289 24573 1307
rect 24539 1221 24573 1235
rect 24539 1153 24573 1163
rect 24539 1085 24573 1091
rect 24539 1017 24573 1019
rect 24539 981 24573 983
rect 24539 909 24573 915
rect 24539 837 24573 847
rect 24539 765 24573 779
rect 24539 693 24573 711
rect 24539 621 24573 643
rect 24539 549 24573 575
rect 24539 477 24573 507
rect 24539 405 24573 439
rect 24539 351 24573 371
rect 24997 1629 25031 1649
rect 24997 1561 25031 1595
rect 24997 1493 25031 1523
rect 24997 1425 25031 1451
rect 24997 1357 25031 1379
rect 24997 1289 25031 1307
rect 24997 1221 25031 1235
rect 24997 1153 25031 1163
rect 24997 1085 25031 1091
rect 24997 1017 25031 1019
rect 24997 981 25031 983
rect 24997 909 25031 915
rect 24997 837 25031 847
rect 24997 765 25031 779
rect 24997 693 25031 711
rect 24997 621 25031 643
rect 24997 549 25031 575
rect 24997 477 25031 507
rect 24997 405 25031 439
rect 24997 270 25031 371
rect 25455 1629 25489 1690
rect 25455 1561 25489 1595
rect 25455 1493 25489 1523
rect 25455 1425 25489 1451
rect 25455 1357 25489 1379
rect 25455 1289 25489 1307
rect 25455 1221 25489 1235
rect 25455 1153 25489 1163
rect 25455 1085 25489 1091
rect 25455 1017 25489 1019
rect 25455 981 25489 983
rect 25455 909 25489 915
rect 25455 837 25489 847
rect 25455 765 25489 779
rect 25455 693 25489 711
rect 25455 621 25489 643
rect 25455 549 25489 575
rect 25455 477 25489 507
rect 25455 405 25489 439
rect 25455 351 25489 371
rect 25913 1629 25947 1649
rect 25913 1561 25947 1595
rect 25913 1493 25947 1523
rect 25913 1425 25947 1451
rect 25913 1357 25947 1379
rect 25913 1289 25947 1307
rect 25913 1221 25947 1235
rect 25913 1153 25947 1163
rect 25913 1085 25947 1091
rect 25913 1017 25947 1019
rect 25913 981 25947 983
rect 25913 909 25947 915
rect 25913 837 25947 847
rect 25913 765 25947 779
rect 25913 693 25947 711
rect 25913 621 25947 643
rect 25913 549 25947 575
rect 25913 477 25947 507
rect 25913 405 25947 439
rect 25913 270 25947 371
rect 26371 1629 26405 1690
rect 26371 1561 26405 1595
rect 26371 1493 26405 1523
rect 26371 1425 26405 1451
rect 26371 1357 26405 1379
rect 26371 1289 26405 1307
rect 26371 1221 26405 1235
rect 26371 1153 26405 1163
rect 26371 1085 26405 1091
rect 26371 1017 26405 1019
rect 26371 981 26405 983
rect 26371 909 26405 915
rect 26371 837 26405 847
rect 26371 765 26405 779
rect 26371 693 26405 711
rect 26371 621 26405 643
rect 26371 549 26405 575
rect 26371 477 26405 507
rect 26371 405 26405 439
rect 26371 351 26405 371
rect 26829 1629 26863 1649
rect 26829 1561 26863 1595
rect 26829 1493 26863 1523
rect 26829 1425 26863 1451
rect 26829 1357 26863 1379
rect 26829 1289 26863 1307
rect 26829 1221 26863 1235
rect 26829 1153 26863 1163
rect 26829 1085 26863 1091
rect 26829 1017 26863 1019
rect 26829 981 26863 983
rect 26829 909 26863 915
rect 26829 837 26863 847
rect 26829 765 26863 779
rect 26829 693 26863 711
rect 26829 621 26863 643
rect 26829 549 26863 575
rect 26829 477 26863 507
rect 26829 405 26863 439
rect 26829 270 26863 371
rect 27287 1629 27321 1690
rect 27287 1561 27321 1595
rect 27287 1493 27321 1523
rect 27287 1425 27321 1451
rect 27287 1357 27321 1379
rect 27287 1289 27321 1307
rect 27287 1221 27321 1235
rect 27287 1153 27321 1163
rect 27287 1085 27321 1091
rect 27287 1017 27321 1019
rect 27287 981 27321 983
rect 27287 909 27321 915
rect 27287 837 27321 847
rect 27287 765 27321 779
rect 27287 693 27321 711
rect 27287 621 27321 643
rect 27287 549 27321 575
rect 27287 477 27321 507
rect 27287 405 27321 439
rect 27287 351 27321 371
rect 27745 1629 27779 1649
rect 27745 1561 27779 1595
rect 27745 1493 27779 1523
rect 27745 1425 27779 1451
rect 27745 1357 27779 1379
rect 27745 1289 27779 1307
rect 27745 1221 27779 1235
rect 27745 1153 27779 1163
rect 27745 1085 27779 1091
rect 27745 1017 27779 1019
rect 27745 981 27779 983
rect 27745 909 27779 915
rect 27745 837 27779 847
rect 27745 765 27779 779
rect 27745 693 27779 711
rect 27745 621 27779 643
rect 27745 549 27779 575
rect 27745 477 27779 507
rect 27745 405 27779 439
rect 27745 270 27779 371
rect 218 210 27826 270
rect 218 151 27826 164
rect 218 117 401 151
rect 435 117 801 151
rect 835 117 1201 151
rect 1235 117 1601 151
rect 1635 117 2001 151
rect 2035 117 2401 151
rect 2435 117 2801 151
rect 2835 117 3201 151
rect 3235 117 3601 151
rect 3635 117 4001 151
rect 4035 117 4401 151
rect 4435 117 4801 151
rect 4835 117 5201 151
rect 5235 117 5601 151
rect 5635 117 6001 151
rect 6035 117 6401 151
rect 6435 117 6801 151
rect 6835 117 7201 151
rect 7235 117 7601 151
rect 7635 117 8001 151
rect 8035 117 8401 151
rect 8435 117 8801 151
rect 8835 117 9201 151
rect 9235 117 9601 151
rect 9635 117 10001 151
rect 10035 117 10401 151
rect 10435 117 10801 151
rect 10835 117 11201 151
rect 11235 117 11601 151
rect 11635 117 12001 151
rect 12035 117 12401 151
rect 12435 117 12801 151
rect 12835 117 13201 151
rect 13235 117 13601 151
rect 13635 117 14001 151
rect 14035 117 14401 151
rect 14435 117 14801 151
rect 14835 117 15201 151
rect 15235 117 15601 151
rect 15635 117 16001 151
rect 16035 117 16401 151
rect 16435 117 16801 151
rect 16835 117 17201 151
rect 17235 117 17601 151
rect 17635 117 18001 151
rect 18035 117 18401 151
rect 18435 117 18801 151
rect 18835 117 19201 151
rect 19235 117 19601 151
rect 19635 117 20001 151
rect 20035 117 20401 151
rect 20435 117 20801 151
rect 20835 117 21201 151
rect 21235 117 21601 151
rect 21635 117 22001 151
rect 22035 117 22401 151
rect 22435 117 22801 151
rect 22835 117 23201 151
rect 23235 117 23601 151
rect 23635 117 24001 151
rect 24035 117 24401 151
rect 24435 117 24801 151
rect 24835 117 25201 151
rect 25235 117 25601 151
rect 25635 117 26001 151
rect 26035 117 26401 151
rect 26435 117 26801 151
rect 26835 117 27201 151
rect 27235 117 27601 151
rect 27635 117 27826 151
rect 218 104 27826 117
rect 120 17 27826 30
rect 120 -17 401 17
rect 435 -17 801 17
rect 835 -17 1201 17
rect 1235 -17 1601 17
rect 1635 -17 2001 17
rect 2035 -17 2401 17
rect 2435 -17 2801 17
rect 2835 -17 3201 17
rect 3235 -17 3601 17
rect 3635 -17 4001 17
rect 4035 -17 4401 17
rect 4435 -17 4801 17
rect 4835 -17 5201 17
rect 5235 -17 5601 17
rect 5635 -17 6001 17
rect 6035 -17 6401 17
rect 6435 -17 6801 17
rect 6835 -17 7201 17
rect 7235 -17 7601 17
rect 7635 -17 8001 17
rect 8035 -17 8401 17
rect 8435 -17 8801 17
rect 8835 -17 9201 17
rect 9235 -17 9601 17
rect 9635 -17 10001 17
rect 10035 -17 10401 17
rect 10435 -17 10801 17
rect 10835 -17 11201 17
rect 11235 -17 11601 17
rect 11635 -17 12001 17
rect 12035 -17 12401 17
rect 12435 -17 12801 17
rect 12835 -17 13201 17
rect 13235 -17 13601 17
rect 13635 -17 14001 17
rect 14035 -17 14401 17
rect 14435 -17 14801 17
rect 14835 -17 15201 17
rect 15235 -17 15601 17
rect 15635 -17 16001 17
rect 16035 -17 16401 17
rect 16435 -17 16801 17
rect 16835 -17 17201 17
rect 17235 -17 17601 17
rect 17635 -17 18001 17
rect 18035 -17 18401 17
rect 18435 -17 18801 17
rect 18835 -17 19201 17
rect 19235 -17 19601 17
rect 19635 -17 20001 17
rect 20035 -17 20401 17
rect 20435 -17 20801 17
rect 20835 -17 21201 17
rect 21235 -17 21601 17
rect 21635 -17 22001 17
rect 22035 -17 22401 17
rect 22435 -17 22801 17
rect 22835 -17 23201 17
rect 23235 -17 23601 17
rect 23635 -17 24001 17
rect 24035 -17 24401 17
rect 24435 -17 24801 17
rect 24835 -17 25201 17
rect 25235 -17 25601 17
rect 25635 -17 26001 17
rect 26035 -17 26401 17
rect 26435 -17 26801 17
rect 26835 -17 27201 17
rect 27235 -17 27601 17
rect 27635 -17 27826 17
rect 120 -30 27826 -17
<< viali >>
rect 401 1863 435 1897
rect 801 1863 835 1897
rect 1201 1863 1235 1897
rect 1601 1863 1635 1897
rect 2001 1863 2035 1897
rect 2401 1863 2435 1897
rect 2801 1863 2835 1897
rect 3201 1863 3235 1897
rect 3601 1863 3635 1897
rect 4001 1863 4035 1897
rect 4401 1863 4435 1897
rect 4801 1863 4835 1897
rect 5201 1863 5235 1897
rect 5601 1863 5635 1897
rect 6001 1863 6035 1897
rect 6401 1863 6435 1897
rect 6801 1863 6835 1897
rect 7201 1863 7235 1897
rect 7601 1863 7635 1897
rect 8001 1863 8035 1897
rect 8401 1863 8435 1897
rect 8801 1863 8835 1897
rect 9201 1863 9235 1897
rect 9601 1863 9635 1897
rect 10001 1863 10035 1897
rect 10401 1863 10435 1897
rect 10801 1863 10835 1897
rect 11201 1863 11235 1897
rect 11601 1863 11635 1897
rect 12001 1863 12035 1897
rect 12401 1863 12435 1897
rect 12801 1863 12835 1897
rect 13201 1863 13235 1897
rect 13601 1863 13635 1897
rect 14001 1863 14035 1897
rect 14401 1863 14435 1897
rect 14801 1863 14835 1897
rect 15201 1863 15235 1897
rect 15601 1863 15635 1897
rect 16001 1863 16035 1897
rect 16401 1863 16435 1897
rect 16801 1863 16835 1897
rect 17201 1863 17235 1897
rect 17601 1863 17635 1897
rect 18001 1863 18035 1897
rect 18401 1863 18435 1897
rect 18801 1863 18835 1897
rect 19201 1863 19235 1897
rect 19601 1863 19635 1897
rect 20001 1863 20035 1897
rect 20401 1863 20435 1897
rect 20801 1863 20835 1897
rect 21201 1863 21235 1897
rect 21601 1863 21635 1897
rect 22001 1863 22035 1897
rect 22401 1863 22435 1897
rect 22801 1863 22835 1897
rect 23201 1863 23235 1897
rect 23601 1863 23635 1897
rect 24001 1863 24035 1897
rect 24401 1863 24435 1897
rect 24801 1863 24835 1897
rect 25201 1863 25235 1897
rect 25601 1863 25635 1897
rect 26001 1863 26035 1897
rect 26401 1863 26435 1897
rect 26801 1863 26835 1897
rect 27201 1863 27235 1897
rect 27601 1863 27635 1897
rect 265 1595 299 1629
rect 265 1527 299 1557
rect 265 1523 299 1527
rect 265 1459 299 1485
rect 265 1451 299 1459
rect 265 1391 299 1413
rect 265 1379 299 1391
rect 265 1323 299 1341
rect 265 1307 299 1323
rect 265 1255 299 1269
rect 265 1235 299 1255
rect 265 1187 299 1197
rect 265 1163 299 1187
rect 265 1119 299 1125
rect 265 1091 299 1119
rect 265 1051 299 1053
rect 265 1019 299 1051
rect 265 949 299 981
rect 265 947 299 949
rect 265 881 299 909
rect 265 875 299 881
rect 265 813 299 837
rect 265 803 299 813
rect 265 745 299 765
rect 265 731 299 745
rect 265 677 299 693
rect 265 659 299 677
rect 265 609 299 621
rect 265 587 299 609
rect 265 541 299 549
rect 265 515 299 541
rect 265 473 299 477
rect 265 443 299 473
rect 265 371 299 405
rect 723 1595 757 1629
rect 723 1527 757 1557
rect 723 1523 757 1527
rect 723 1459 757 1485
rect 723 1451 757 1459
rect 723 1391 757 1413
rect 723 1379 757 1391
rect 723 1323 757 1341
rect 723 1307 757 1323
rect 723 1255 757 1269
rect 723 1235 757 1255
rect 723 1187 757 1197
rect 723 1163 757 1187
rect 723 1119 757 1125
rect 723 1091 757 1119
rect 723 1051 757 1053
rect 723 1019 757 1051
rect 723 949 757 981
rect 723 947 757 949
rect 723 881 757 909
rect 723 875 757 881
rect 723 813 757 837
rect 723 803 757 813
rect 723 745 757 765
rect 723 731 757 745
rect 723 677 757 693
rect 723 659 757 677
rect 723 609 757 621
rect 723 587 757 609
rect 723 541 757 549
rect 723 515 757 541
rect 723 473 757 477
rect 723 443 757 473
rect 723 371 757 405
rect 1181 1595 1215 1629
rect 1181 1527 1215 1557
rect 1181 1523 1215 1527
rect 1181 1459 1215 1485
rect 1181 1451 1215 1459
rect 1181 1391 1215 1413
rect 1181 1379 1215 1391
rect 1181 1323 1215 1341
rect 1181 1307 1215 1323
rect 1181 1255 1215 1269
rect 1181 1235 1215 1255
rect 1181 1187 1215 1197
rect 1181 1163 1215 1187
rect 1181 1119 1215 1125
rect 1181 1091 1215 1119
rect 1181 1051 1215 1053
rect 1181 1019 1215 1051
rect 1181 949 1215 981
rect 1181 947 1215 949
rect 1181 881 1215 909
rect 1181 875 1215 881
rect 1181 813 1215 837
rect 1181 803 1215 813
rect 1181 745 1215 765
rect 1181 731 1215 745
rect 1181 677 1215 693
rect 1181 659 1215 677
rect 1181 609 1215 621
rect 1181 587 1215 609
rect 1181 541 1215 549
rect 1181 515 1215 541
rect 1181 473 1215 477
rect 1181 443 1215 473
rect 1181 371 1215 405
rect 1639 1595 1673 1629
rect 1639 1527 1673 1557
rect 1639 1523 1673 1527
rect 1639 1459 1673 1485
rect 1639 1451 1673 1459
rect 1639 1391 1673 1413
rect 1639 1379 1673 1391
rect 1639 1323 1673 1341
rect 1639 1307 1673 1323
rect 1639 1255 1673 1269
rect 1639 1235 1673 1255
rect 1639 1187 1673 1197
rect 1639 1163 1673 1187
rect 1639 1119 1673 1125
rect 1639 1091 1673 1119
rect 1639 1051 1673 1053
rect 1639 1019 1673 1051
rect 1639 949 1673 981
rect 1639 947 1673 949
rect 1639 881 1673 909
rect 1639 875 1673 881
rect 1639 813 1673 837
rect 1639 803 1673 813
rect 1639 745 1673 765
rect 1639 731 1673 745
rect 1639 677 1673 693
rect 1639 659 1673 677
rect 1639 609 1673 621
rect 1639 587 1673 609
rect 1639 541 1673 549
rect 1639 515 1673 541
rect 1639 473 1673 477
rect 1639 443 1673 473
rect 1639 371 1673 405
rect 2097 1595 2131 1629
rect 2097 1527 2131 1557
rect 2097 1523 2131 1527
rect 2097 1459 2131 1485
rect 2097 1451 2131 1459
rect 2097 1391 2131 1413
rect 2097 1379 2131 1391
rect 2097 1323 2131 1341
rect 2097 1307 2131 1323
rect 2097 1255 2131 1269
rect 2097 1235 2131 1255
rect 2097 1187 2131 1197
rect 2097 1163 2131 1187
rect 2097 1119 2131 1125
rect 2097 1091 2131 1119
rect 2097 1051 2131 1053
rect 2097 1019 2131 1051
rect 2097 949 2131 981
rect 2097 947 2131 949
rect 2097 881 2131 909
rect 2097 875 2131 881
rect 2097 813 2131 837
rect 2097 803 2131 813
rect 2097 745 2131 765
rect 2097 731 2131 745
rect 2097 677 2131 693
rect 2097 659 2131 677
rect 2097 609 2131 621
rect 2097 587 2131 609
rect 2097 541 2131 549
rect 2097 515 2131 541
rect 2097 473 2131 477
rect 2097 443 2131 473
rect 2097 371 2131 405
rect 2555 1595 2589 1629
rect 2555 1527 2589 1557
rect 2555 1523 2589 1527
rect 2555 1459 2589 1485
rect 2555 1451 2589 1459
rect 2555 1391 2589 1413
rect 2555 1379 2589 1391
rect 2555 1323 2589 1341
rect 2555 1307 2589 1323
rect 2555 1255 2589 1269
rect 2555 1235 2589 1255
rect 2555 1187 2589 1197
rect 2555 1163 2589 1187
rect 2555 1119 2589 1125
rect 2555 1091 2589 1119
rect 2555 1051 2589 1053
rect 2555 1019 2589 1051
rect 2555 949 2589 981
rect 2555 947 2589 949
rect 2555 881 2589 909
rect 2555 875 2589 881
rect 2555 813 2589 837
rect 2555 803 2589 813
rect 2555 745 2589 765
rect 2555 731 2589 745
rect 2555 677 2589 693
rect 2555 659 2589 677
rect 2555 609 2589 621
rect 2555 587 2589 609
rect 2555 541 2589 549
rect 2555 515 2589 541
rect 2555 473 2589 477
rect 2555 443 2589 473
rect 2555 371 2589 405
rect 3013 1595 3047 1629
rect 3013 1527 3047 1557
rect 3013 1523 3047 1527
rect 3013 1459 3047 1485
rect 3013 1451 3047 1459
rect 3013 1391 3047 1413
rect 3013 1379 3047 1391
rect 3013 1323 3047 1341
rect 3013 1307 3047 1323
rect 3013 1255 3047 1269
rect 3013 1235 3047 1255
rect 3013 1187 3047 1197
rect 3013 1163 3047 1187
rect 3013 1119 3047 1125
rect 3013 1091 3047 1119
rect 3013 1051 3047 1053
rect 3013 1019 3047 1051
rect 3013 949 3047 981
rect 3013 947 3047 949
rect 3013 881 3047 909
rect 3013 875 3047 881
rect 3013 813 3047 837
rect 3013 803 3047 813
rect 3013 745 3047 765
rect 3013 731 3047 745
rect 3013 677 3047 693
rect 3013 659 3047 677
rect 3013 609 3047 621
rect 3013 587 3047 609
rect 3013 541 3047 549
rect 3013 515 3047 541
rect 3013 473 3047 477
rect 3013 443 3047 473
rect 3013 371 3047 405
rect 3471 1595 3505 1629
rect 3471 1527 3505 1557
rect 3471 1523 3505 1527
rect 3471 1459 3505 1485
rect 3471 1451 3505 1459
rect 3471 1391 3505 1413
rect 3471 1379 3505 1391
rect 3471 1323 3505 1341
rect 3471 1307 3505 1323
rect 3471 1255 3505 1269
rect 3471 1235 3505 1255
rect 3471 1187 3505 1197
rect 3471 1163 3505 1187
rect 3471 1119 3505 1125
rect 3471 1091 3505 1119
rect 3471 1051 3505 1053
rect 3471 1019 3505 1051
rect 3471 949 3505 981
rect 3471 947 3505 949
rect 3471 881 3505 909
rect 3471 875 3505 881
rect 3471 813 3505 837
rect 3471 803 3505 813
rect 3471 745 3505 765
rect 3471 731 3505 745
rect 3471 677 3505 693
rect 3471 659 3505 677
rect 3471 609 3505 621
rect 3471 587 3505 609
rect 3471 541 3505 549
rect 3471 515 3505 541
rect 3471 473 3505 477
rect 3471 443 3505 473
rect 3471 371 3505 405
rect 3929 1595 3963 1629
rect 3929 1527 3963 1557
rect 3929 1523 3963 1527
rect 3929 1459 3963 1485
rect 3929 1451 3963 1459
rect 3929 1391 3963 1413
rect 3929 1379 3963 1391
rect 3929 1323 3963 1341
rect 3929 1307 3963 1323
rect 3929 1255 3963 1269
rect 3929 1235 3963 1255
rect 3929 1187 3963 1197
rect 3929 1163 3963 1187
rect 3929 1119 3963 1125
rect 3929 1091 3963 1119
rect 3929 1051 3963 1053
rect 3929 1019 3963 1051
rect 3929 949 3963 981
rect 3929 947 3963 949
rect 3929 881 3963 909
rect 3929 875 3963 881
rect 3929 813 3963 837
rect 3929 803 3963 813
rect 3929 745 3963 765
rect 3929 731 3963 745
rect 3929 677 3963 693
rect 3929 659 3963 677
rect 3929 609 3963 621
rect 3929 587 3963 609
rect 3929 541 3963 549
rect 3929 515 3963 541
rect 3929 473 3963 477
rect 3929 443 3963 473
rect 3929 371 3963 405
rect 4387 1595 4421 1629
rect 4387 1527 4421 1557
rect 4387 1523 4421 1527
rect 4387 1459 4421 1485
rect 4387 1451 4421 1459
rect 4387 1391 4421 1413
rect 4387 1379 4421 1391
rect 4387 1323 4421 1341
rect 4387 1307 4421 1323
rect 4387 1255 4421 1269
rect 4387 1235 4421 1255
rect 4387 1187 4421 1197
rect 4387 1163 4421 1187
rect 4387 1119 4421 1125
rect 4387 1091 4421 1119
rect 4387 1051 4421 1053
rect 4387 1019 4421 1051
rect 4387 949 4421 981
rect 4387 947 4421 949
rect 4387 881 4421 909
rect 4387 875 4421 881
rect 4387 813 4421 837
rect 4387 803 4421 813
rect 4387 745 4421 765
rect 4387 731 4421 745
rect 4387 677 4421 693
rect 4387 659 4421 677
rect 4387 609 4421 621
rect 4387 587 4421 609
rect 4387 541 4421 549
rect 4387 515 4421 541
rect 4387 473 4421 477
rect 4387 443 4421 473
rect 4387 371 4421 405
rect 4845 1595 4879 1629
rect 4845 1527 4879 1557
rect 4845 1523 4879 1527
rect 4845 1459 4879 1485
rect 4845 1451 4879 1459
rect 4845 1391 4879 1413
rect 4845 1379 4879 1391
rect 4845 1323 4879 1341
rect 4845 1307 4879 1323
rect 4845 1255 4879 1269
rect 4845 1235 4879 1255
rect 4845 1187 4879 1197
rect 4845 1163 4879 1187
rect 4845 1119 4879 1125
rect 4845 1091 4879 1119
rect 4845 1051 4879 1053
rect 4845 1019 4879 1051
rect 4845 949 4879 981
rect 4845 947 4879 949
rect 4845 881 4879 909
rect 4845 875 4879 881
rect 4845 813 4879 837
rect 4845 803 4879 813
rect 4845 745 4879 765
rect 4845 731 4879 745
rect 4845 677 4879 693
rect 4845 659 4879 677
rect 4845 609 4879 621
rect 4845 587 4879 609
rect 4845 541 4879 549
rect 4845 515 4879 541
rect 4845 473 4879 477
rect 4845 443 4879 473
rect 4845 371 4879 405
rect 5303 1595 5337 1629
rect 5303 1527 5337 1557
rect 5303 1523 5337 1527
rect 5303 1459 5337 1485
rect 5303 1451 5337 1459
rect 5303 1391 5337 1413
rect 5303 1379 5337 1391
rect 5303 1323 5337 1341
rect 5303 1307 5337 1323
rect 5303 1255 5337 1269
rect 5303 1235 5337 1255
rect 5303 1187 5337 1197
rect 5303 1163 5337 1187
rect 5303 1119 5337 1125
rect 5303 1091 5337 1119
rect 5303 1051 5337 1053
rect 5303 1019 5337 1051
rect 5303 949 5337 981
rect 5303 947 5337 949
rect 5303 881 5337 909
rect 5303 875 5337 881
rect 5303 813 5337 837
rect 5303 803 5337 813
rect 5303 745 5337 765
rect 5303 731 5337 745
rect 5303 677 5337 693
rect 5303 659 5337 677
rect 5303 609 5337 621
rect 5303 587 5337 609
rect 5303 541 5337 549
rect 5303 515 5337 541
rect 5303 473 5337 477
rect 5303 443 5337 473
rect 5303 371 5337 405
rect 5761 1595 5795 1629
rect 5761 1527 5795 1557
rect 5761 1523 5795 1527
rect 5761 1459 5795 1485
rect 5761 1451 5795 1459
rect 5761 1391 5795 1413
rect 5761 1379 5795 1391
rect 5761 1323 5795 1341
rect 5761 1307 5795 1323
rect 5761 1255 5795 1269
rect 5761 1235 5795 1255
rect 5761 1187 5795 1197
rect 5761 1163 5795 1187
rect 5761 1119 5795 1125
rect 5761 1091 5795 1119
rect 5761 1051 5795 1053
rect 5761 1019 5795 1051
rect 5761 949 5795 981
rect 5761 947 5795 949
rect 5761 881 5795 909
rect 5761 875 5795 881
rect 5761 813 5795 837
rect 5761 803 5795 813
rect 5761 745 5795 765
rect 5761 731 5795 745
rect 5761 677 5795 693
rect 5761 659 5795 677
rect 5761 609 5795 621
rect 5761 587 5795 609
rect 5761 541 5795 549
rect 5761 515 5795 541
rect 5761 473 5795 477
rect 5761 443 5795 473
rect 5761 371 5795 405
rect 6219 1595 6253 1629
rect 6219 1527 6253 1557
rect 6219 1523 6253 1527
rect 6219 1459 6253 1485
rect 6219 1451 6253 1459
rect 6219 1391 6253 1413
rect 6219 1379 6253 1391
rect 6219 1323 6253 1341
rect 6219 1307 6253 1323
rect 6219 1255 6253 1269
rect 6219 1235 6253 1255
rect 6219 1187 6253 1197
rect 6219 1163 6253 1187
rect 6219 1119 6253 1125
rect 6219 1091 6253 1119
rect 6219 1051 6253 1053
rect 6219 1019 6253 1051
rect 6219 949 6253 981
rect 6219 947 6253 949
rect 6219 881 6253 909
rect 6219 875 6253 881
rect 6219 813 6253 837
rect 6219 803 6253 813
rect 6219 745 6253 765
rect 6219 731 6253 745
rect 6219 677 6253 693
rect 6219 659 6253 677
rect 6219 609 6253 621
rect 6219 587 6253 609
rect 6219 541 6253 549
rect 6219 515 6253 541
rect 6219 473 6253 477
rect 6219 443 6253 473
rect 6219 371 6253 405
rect 6677 1595 6711 1629
rect 6677 1527 6711 1557
rect 6677 1523 6711 1527
rect 6677 1459 6711 1485
rect 6677 1451 6711 1459
rect 6677 1391 6711 1413
rect 6677 1379 6711 1391
rect 6677 1323 6711 1341
rect 6677 1307 6711 1323
rect 6677 1255 6711 1269
rect 6677 1235 6711 1255
rect 6677 1187 6711 1197
rect 6677 1163 6711 1187
rect 6677 1119 6711 1125
rect 6677 1091 6711 1119
rect 6677 1051 6711 1053
rect 6677 1019 6711 1051
rect 6677 949 6711 981
rect 6677 947 6711 949
rect 6677 881 6711 909
rect 6677 875 6711 881
rect 6677 813 6711 837
rect 6677 803 6711 813
rect 6677 745 6711 765
rect 6677 731 6711 745
rect 6677 677 6711 693
rect 6677 659 6711 677
rect 6677 609 6711 621
rect 6677 587 6711 609
rect 6677 541 6711 549
rect 6677 515 6711 541
rect 6677 473 6711 477
rect 6677 443 6711 473
rect 6677 371 6711 405
rect 7135 1595 7169 1629
rect 7135 1527 7169 1557
rect 7135 1523 7169 1527
rect 7135 1459 7169 1485
rect 7135 1451 7169 1459
rect 7135 1391 7169 1413
rect 7135 1379 7169 1391
rect 7135 1323 7169 1341
rect 7135 1307 7169 1323
rect 7135 1255 7169 1269
rect 7135 1235 7169 1255
rect 7135 1187 7169 1197
rect 7135 1163 7169 1187
rect 7135 1119 7169 1125
rect 7135 1091 7169 1119
rect 7135 1051 7169 1053
rect 7135 1019 7169 1051
rect 7135 949 7169 981
rect 7135 947 7169 949
rect 7135 881 7169 909
rect 7135 875 7169 881
rect 7135 813 7169 837
rect 7135 803 7169 813
rect 7135 745 7169 765
rect 7135 731 7169 745
rect 7135 677 7169 693
rect 7135 659 7169 677
rect 7135 609 7169 621
rect 7135 587 7169 609
rect 7135 541 7169 549
rect 7135 515 7169 541
rect 7135 473 7169 477
rect 7135 443 7169 473
rect 7135 371 7169 405
rect 7593 1595 7627 1629
rect 7593 1527 7627 1557
rect 7593 1523 7627 1527
rect 7593 1459 7627 1485
rect 7593 1451 7627 1459
rect 7593 1391 7627 1413
rect 7593 1379 7627 1391
rect 7593 1323 7627 1341
rect 7593 1307 7627 1323
rect 7593 1255 7627 1269
rect 7593 1235 7627 1255
rect 7593 1187 7627 1197
rect 7593 1163 7627 1187
rect 7593 1119 7627 1125
rect 7593 1091 7627 1119
rect 7593 1051 7627 1053
rect 7593 1019 7627 1051
rect 7593 949 7627 981
rect 7593 947 7627 949
rect 7593 881 7627 909
rect 7593 875 7627 881
rect 7593 813 7627 837
rect 7593 803 7627 813
rect 7593 745 7627 765
rect 7593 731 7627 745
rect 7593 677 7627 693
rect 7593 659 7627 677
rect 7593 609 7627 621
rect 7593 587 7627 609
rect 7593 541 7627 549
rect 7593 515 7627 541
rect 7593 473 7627 477
rect 7593 443 7627 473
rect 7593 371 7627 405
rect 8051 1595 8085 1629
rect 8051 1527 8085 1557
rect 8051 1523 8085 1527
rect 8051 1459 8085 1485
rect 8051 1451 8085 1459
rect 8051 1391 8085 1413
rect 8051 1379 8085 1391
rect 8051 1323 8085 1341
rect 8051 1307 8085 1323
rect 8051 1255 8085 1269
rect 8051 1235 8085 1255
rect 8051 1187 8085 1197
rect 8051 1163 8085 1187
rect 8051 1119 8085 1125
rect 8051 1091 8085 1119
rect 8051 1051 8085 1053
rect 8051 1019 8085 1051
rect 8051 949 8085 981
rect 8051 947 8085 949
rect 8051 881 8085 909
rect 8051 875 8085 881
rect 8051 813 8085 837
rect 8051 803 8085 813
rect 8051 745 8085 765
rect 8051 731 8085 745
rect 8051 677 8085 693
rect 8051 659 8085 677
rect 8051 609 8085 621
rect 8051 587 8085 609
rect 8051 541 8085 549
rect 8051 515 8085 541
rect 8051 473 8085 477
rect 8051 443 8085 473
rect 8051 371 8085 405
rect 8509 1595 8543 1629
rect 8509 1527 8543 1557
rect 8509 1523 8543 1527
rect 8509 1459 8543 1485
rect 8509 1451 8543 1459
rect 8509 1391 8543 1413
rect 8509 1379 8543 1391
rect 8509 1323 8543 1341
rect 8509 1307 8543 1323
rect 8509 1255 8543 1269
rect 8509 1235 8543 1255
rect 8509 1187 8543 1197
rect 8509 1163 8543 1187
rect 8509 1119 8543 1125
rect 8509 1091 8543 1119
rect 8509 1051 8543 1053
rect 8509 1019 8543 1051
rect 8509 949 8543 981
rect 8509 947 8543 949
rect 8509 881 8543 909
rect 8509 875 8543 881
rect 8509 813 8543 837
rect 8509 803 8543 813
rect 8509 745 8543 765
rect 8509 731 8543 745
rect 8509 677 8543 693
rect 8509 659 8543 677
rect 8509 609 8543 621
rect 8509 587 8543 609
rect 8509 541 8543 549
rect 8509 515 8543 541
rect 8509 473 8543 477
rect 8509 443 8543 473
rect 8509 371 8543 405
rect 8967 1595 9001 1629
rect 8967 1527 9001 1557
rect 8967 1523 9001 1527
rect 8967 1459 9001 1485
rect 8967 1451 9001 1459
rect 8967 1391 9001 1413
rect 8967 1379 9001 1391
rect 8967 1323 9001 1341
rect 8967 1307 9001 1323
rect 8967 1255 9001 1269
rect 8967 1235 9001 1255
rect 8967 1187 9001 1197
rect 8967 1163 9001 1187
rect 8967 1119 9001 1125
rect 8967 1091 9001 1119
rect 8967 1051 9001 1053
rect 8967 1019 9001 1051
rect 8967 949 9001 981
rect 8967 947 9001 949
rect 8967 881 9001 909
rect 8967 875 9001 881
rect 8967 813 9001 837
rect 8967 803 9001 813
rect 8967 745 9001 765
rect 8967 731 9001 745
rect 8967 677 9001 693
rect 8967 659 9001 677
rect 8967 609 9001 621
rect 8967 587 9001 609
rect 8967 541 9001 549
rect 8967 515 9001 541
rect 8967 473 9001 477
rect 8967 443 9001 473
rect 8967 371 9001 405
rect 9425 1595 9459 1629
rect 9425 1527 9459 1557
rect 9425 1523 9459 1527
rect 9425 1459 9459 1485
rect 9425 1451 9459 1459
rect 9425 1391 9459 1413
rect 9425 1379 9459 1391
rect 9425 1323 9459 1341
rect 9425 1307 9459 1323
rect 9425 1255 9459 1269
rect 9425 1235 9459 1255
rect 9425 1187 9459 1197
rect 9425 1163 9459 1187
rect 9425 1119 9459 1125
rect 9425 1091 9459 1119
rect 9425 1051 9459 1053
rect 9425 1019 9459 1051
rect 9425 949 9459 981
rect 9425 947 9459 949
rect 9425 881 9459 909
rect 9425 875 9459 881
rect 9425 813 9459 837
rect 9425 803 9459 813
rect 9425 745 9459 765
rect 9425 731 9459 745
rect 9425 677 9459 693
rect 9425 659 9459 677
rect 9425 609 9459 621
rect 9425 587 9459 609
rect 9425 541 9459 549
rect 9425 515 9459 541
rect 9425 473 9459 477
rect 9425 443 9459 473
rect 9425 371 9459 405
rect 9883 1595 9917 1629
rect 9883 1527 9917 1557
rect 9883 1523 9917 1527
rect 9883 1459 9917 1485
rect 9883 1451 9917 1459
rect 9883 1391 9917 1413
rect 9883 1379 9917 1391
rect 9883 1323 9917 1341
rect 9883 1307 9917 1323
rect 9883 1255 9917 1269
rect 9883 1235 9917 1255
rect 9883 1187 9917 1197
rect 9883 1163 9917 1187
rect 9883 1119 9917 1125
rect 9883 1091 9917 1119
rect 9883 1051 9917 1053
rect 9883 1019 9917 1051
rect 9883 949 9917 981
rect 9883 947 9917 949
rect 9883 881 9917 909
rect 9883 875 9917 881
rect 9883 813 9917 837
rect 9883 803 9917 813
rect 9883 745 9917 765
rect 9883 731 9917 745
rect 9883 677 9917 693
rect 9883 659 9917 677
rect 9883 609 9917 621
rect 9883 587 9917 609
rect 9883 541 9917 549
rect 9883 515 9917 541
rect 9883 473 9917 477
rect 9883 443 9917 473
rect 9883 371 9917 405
rect 10341 1595 10375 1629
rect 10341 1527 10375 1557
rect 10341 1523 10375 1527
rect 10341 1459 10375 1485
rect 10341 1451 10375 1459
rect 10341 1391 10375 1413
rect 10341 1379 10375 1391
rect 10341 1323 10375 1341
rect 10341 1307 10375 1323
rect 10341 1255 10375 1269
rect 10341 1235 10375 1255
rect 10341 1187 10375 1197
rect 10341 1163 10375 1187
rect 10341 1119 10375 1125
rect 10341 1091 10375 1119
rect 10341 1051 10375 1053
rect 10341 1019 10375 1051
rect 10341 949 10375 981
rect 10341 947 10375 949
rect 10341 881 10375 909
rect 10341 875 10375 881
rect 10341 813 10375 837
rect 10341 803 10375 813
rect 10341 745 10375 765
rect 10341 731 10375 745
rect 10341 677 10375 693
rect 10341 659 10375 677
rect 10341 609 10375 621
rect 10341 587 10375 609
rect 10341 541 10375 549
rect 10341 515 10375 541
rect 10341 473 10375 477
rect 10341 443 10375 473
rect 10341 371 10375 405
rect 10799 1595 10833 1629
rect 10799 1527 10833 1557
rect 10799 1523 10833 1527
rect 10799 1459 10833 1485
rect 10799 1451 10833 1459
rect 10799 1391 10833 1413
rect 10799 1379 10833 1391
rect 10799 1323 10833 1341
rect 10799 1307 10833 1323
rect 10799 1255 10833 1269
rect 10799 1235 10833 1255
rect 10799 1187 10833 1197
rect 10799 1163 10833 1187
rect 10799 1119 10833 1125
rect 10799 1091 10833 1119
rect 10799 1051 10833 1053
rect 10799 1019 10833 1051
rect 10799 949 10833 981
rect 10799 947 10833 949
rect 10799 881 10833 909
rect 10799 875 10833 881
rect 10799 813 10833 837
rect 10799 803 10833 813
rect 10799 745 10833 765
rect 10799 731 10833 745
rect 10799 677 10833 693
rect 10799 659 10833 677
rect 10799 609 10833 621
rect 10799 587 10833 609
rect 10799 541 10833 549
rect 10799 515 10833 541
rect 10799 473 10833 477
rect 10799 443 10833 473
rect 10799 371 10833 405
rect 11257 1595 11291 1629
rect 11257 1527 11291 1557
rect 11257 1523 11291 1527
rect 11257 1459 11291 1485
rect 11257 1451 11291 1459
rect 11257 1391 11291 1413
rect 11257 1379 11291 1391
rect 11257 1323 11291 1341
rect 11257 1307 11291 1323
rect 11257 1255 11291 1269
rect 11257 1235 11291 1255
rect 11257 1187 11291 1197
rect 11257 1163 11291 1187
rect 11257 1119 11291 1125
rect 11257 1091 11291 1119
rect 11257 1051 11291 1053
rect 11257 1019 11291 1051
rect 11257 949 11291 981
rect 11257 947 11291 949
rect 11257 881 11291 909
rect 11257 875 11291 881
rect 11257 813 11291 837
rect 11257 803 11291 813
rect 11257 745 11291 765
rect 11257 731 11291 745
rect 11257 677 11291 693
rect 11257 659 11291 677
rect 11257 609 11291 621
rect 11257 587 11291 609
rect 11257 541 11291 549
rect 11257 515 11291 541
rect 11257 473 11291 477
rect 11257 443 11291 473
rect 11257 371 11291 405
rect 11715 1595 11749 1629
rect 11715 1527 11749 1557
rect 11715 1523 11749 1527
rect 11715 1459 11749 1485
rect 11715 1451 11749 1459
rect 11715 1391 11749 1413
rect 11715 1379 11749 1391
rect 11715 1323 11749 1341
rect 11715 1307 11749 1323
rect 11715 1255 11749 1269
rect 11715 1235 11749 1255
rect 11715 1187 11749 1197
rect 11715 1163 11749 1187
rect 11715 1119 11749 1125
rect 11715 1091 11749 1119
rect 11715 1051 11749 1053
rect 11715 1019 11749 1051
rect 11715 949 11749 981
rect 11715 947 11749 949
rect 11715 881 11749 909
rect 11715 875 11749 881
rect 11715 813 11749 837
rect 11715 803 11749 813
rect 11715 745 11749 765
rect 11715 731 11749 745
rect 11715 677 11749 693
rect 11715 659 11749 677
rect 11715 609 11749 621
rect 11715 587 11749 609
rect 11715 541 11749 549
rect 11715 515 11749 541
rect 11715 473 11749 477
rect 11715 443 11749 473
rect 11715 371 11749 405
rect 12173 1595 12207 1629
rect 12173 1527 12207 1557
rect 12173 1523 12207 1527
rect 12173 1459 12207 1485
rect 12173 1451 12207 1459
rect 12173 1391 12207 1413
rect 12173 1379 12207 1391
rect 12173 1323 12207 1341
rect 12173 1307 12207 1323
rect 12173 1255 12207 1269
rect 12173 1235 12207 1255
rect 12173 1187 12207 1197
rect 12173 1163 12207 1187
rect 12173 1119 12207 1125
rect 12173 1091 12207 1119
rect 12173 1051 12207 1053
rect 12173 1019 12207 1051
rect 12173 949 12207 981
rect 12173 947 12207 949
rect 12173 881 12207 909
rect 12173 875 12207 881
rect 12173 813 12207 837
rect 12173 803 12207 813
rect 12173 745 12207 765
rect 12173 731 12207 745
rect 12173 677 12207 693
rect 12173 659 12207 677
rect 12173 609 12207 621
rect 12173 587 12207 609
rect 12173 541 12207 549
rect 12173 515 12207 541
rect 12173 473 12207 477
rect 12173 443 12207 473
rect 12173 371 12207 405
rect 12631 1595 12665 1629
rect 12631 1527 12665 1557
rect 12631 1523 12665 1527
rect 12631 1459 12665 1485
rect 12631 1451 12665 1459
rect 12631 1391 12665 1413
rect 12631 1379 12665 1391
rect 12631 1323 12665 1341
rect 12631 1307 12665 1323
rect 12631 1255 12665 1269
rect 12631 1235 12665 1255
rect 12631 1187 12665 1197
rect 12631 1163 12665 1187
rect 12631 1119 12665 1125
rect 12631 1091 12665 1119
rect 12631 1051 12665 1053
rect 12631 1019 12665 1051
rect 12631 949 12665 981
rect 12631 947 12665 949
rect 12631 881 12665 909
rect 12631 875 12665 881
rect 12631 813 12665 837
rect 12631 803 12665 813
rect 12631 745 12665 765
rect 12631 731 12665 745
rect 12631 677 12665 693
rect 12631 659 12665 677
rect 12631 609 12665 621
rect 12631 587 12665 609
rect 12631 541 12665 549
rect 12631 515 12665 541
rect 12631 473 12665 477
rect 12631 443 12665 473
rect 12631 371 12665 405
rect 13089 1595 13123 1629
rect 13089 1527 13123 1557
rect 13089 1523 13123 1527
rect 13089 1459 13123 1485
rect 13089 1451 13123 1459
rect 13089 1391 13123 1413
rect 13089 1379 13123 1391
rect 13089 1323 13123 1341
rect 13089 1307 13123 1323
rect 13089 1255 13123 1269
rect 13089 1235 13123 1255
rect 13089 1187 13123 1197
rect 13089 1163 13123 1187
rect 13089 1119 13123 1125
rect 13089 1091 13123 1119
rect 13089 1051 13123 1053
rect 13089 1019 13123 1051
rect 13089 949 13123 981
rect 13089 947 13123 949
rect 13089 881 13123 909
rect 13089 875 13123 881
rect 13089 813 13123 837
rect 13089 803 13123 813
rect 13089 745 13123 765
rect 13089 731 13123 745
rect 13089 677 13123 693
rect 13089 659 13123 677
rect 13089 609 13123 621
rect 13089 587 13123 609
rect 13089 541 13123 549
rect 13089 515 13123 541
rect 13089 473 13123 477
rect 13089 443 13123 473
rect 13089 371 13123 405
rect 13547 1595 13581 1629
rect 13547 1527 13581 1557
rect 13547 1523 13581 1527
rect 13547 1459 13581 1485
rect 13547 1451 13581 1459
rect 13547 1391 13581 1413
rect 13547 1379 13581 1391
rect 13547 1323 13581 1341
rect 13547 1307 13581 1323
rect 13547 1255 13581 1269
rect 13547 1235 13581 1255
rect 13547 1187 13581 1197
rect 13547 1163 13581 1187
rect 13547 1119 13581 1125
rect 13547 1091 13581 1119
rect 13547 1051 13581 1053
rect 13547 1019 13581 1051
rect 13547 949 13581 981
rect 13547 947 13581 949
rect 13547 881 13581 909
rect 13547 875 13581 881
rect 13547 813 13581 837
rect 13547 803 13581 813
rect 13547 745 13581 765
rect 13547 731 13581 745
rect 13547 677 13581 693
rect 13547 659 13581 677
rect 13547 609 13581 621
rect 13547 587 13581 609
rect 13547 541 13581 549
rect 13547 515 13581 541
rect 13547 473 13581 477
rect 13547 443 13581 473
rect 13547 371 13581 405
rect 14005 1595 14039 1629
rect 14005 1527 14039 1557
rect 14005 1523 14039 1527
rect 14005 1459 14039 1485
rect 14005 1451 14039 1459
rect 14005 1391 14039 1413
rect 14005 1379 14039 1391
rect 14005 1323 14039 1341
rect 14005 1307 14039 1323
rect 14005 1255 14039 1269
rect 14005 1235 14039 1255
rect 14005 1187 14039 1197
rect 14005 1163 14039 1187
rect 14005 1119 14039 1125
rect 14005 1091 14039 1119
rect 14005 1051 14039 1053
rect 14005 1019 14039 1051
rect 14005 949 14039 981
rect 14005 947 14039 949
rect 14005 881 14039 909
rect 14005 875 14039 881
rect 14005 813 14039 837
rect 14005 803 14039 813
rect 14005 745 14039 765
rect 14005 731 14039 745
rect 14005 677 14039 693
rect 14005 659 14039 677
rect 14005 609 14039 621
rect 14005 587 14039 609
rect 14005 541 14039 549
rect 14005 515 14039 541
rect 14005 473 14039 477
rect 14005 443 14039 473
rect 14005 371 14039 405
rect 14463 1595 14497 1629
rect 14463 1527 14497 1557
rect 14463 1523 14497 1527
rect 14463 1459 14497 1485
rect 14463 1451 14497 1459
rect 14463 1391 14497 1413
rect 14463 1379 14497 1391
rect 14463 1323 14497 1341
rect 14463 1307 14497 1323
rect 14463 1255 14497 1269
rect 14463 1235 14497 1255
rect 14463 1187 14497 1197
rect 14463 1163 14497 1187
rect 14463 1119 14497 1125
rect 14463 1091 14497 1119
rect 14463 1051 14497 1053
rect 14463 1019 14497 1051
rect 14463 949 14497 981
rect 14463 947 14497 949
rect 14463 881 14497 909
rect 14463 875 14497 881
rect 14463 813 14497 837
rect 14463 803 14497 813
rect 14463 745 14497 765
rect 14463 731 14497 745
rect 14463 677 14497 693
rect 14463 659 14497 677
rect 14463 609 14497 621
rect 14463 587 14497 609
rect 14463 541 14497 549
rect 14463 515 14497 541
rect 14463 473 14497 477
rect 14463 443 14497 473
rect 14463 371 14497 405
rect 14921 1595 14955 1629
rect 14921 1527 14955 1557
rect 14921 1523 14955 1527
rect 14921 1459 14955 1485
rect 14921 1451 14955 1459
rect 14921 1391 14955 1413
rect 14921 1379 14955 1391
rect 14921 1323 14955 1341
rect 14921 1307 14955 1323
rect 14921 1255 14955 1269
rect 14921 1235 14955 1255
rect 14921 1187 14955 1197
rect 14921 1163 14955 1187
rect 14921 1119 14955 1125
rect 14921 1091 14955 1119
rect 14921 1051 14955 1053
rect 14921 1019 14955 1051
rect 14921 949 14955 981
rect 14921 947 14955 949
rect 14921 881 14955 909
rect 14921 875 14955 881
rect 14921 813 14955 837
rect 14921 803 14955 813
rect 14921 745 14955 765
rect 14921 731 14955 745
rect 14921 677 14955 693
rect 14921 659 14955 677
rect 14921 609 14955 621
rect 14921 587 14955 609
rect 14921 541 14955 549
rect 14921 515 14955 541
rect 14921 473 14955 477
rect 14921 443 14955 473
rect 14921 371 14955 405
rect 15379 1595 15413 1629
rect 15379 1527 15413 1557
rect 15379 1523 15413 1527
rect 15379 1459 15413 1485
rect 15379 1451 15413 1459
rect 15379 1391 15413 1413
rect 15379 1379 15413 1391
rect 15379 1323 15413 1341
rect 15379 1307 15413 1323
rect 15379 1255 15413 1269
rect 15379 1235 15413 1255
rect 15379 1187 15413 1197
rect 15379 1163 15413 1187
rect 15379 1119 15413 1125
rect 15379 1091 15413 1119
rect 15379 1051 15413 1053
rect 15379 1019 15413 1051
rect 15379 949 15413 981
rect 15379 947 15413 949
rect 15379 881 15413 909
rect 15379 875 15413 881
rect 15379 813 15413 837
rect 15379 803 15413 813
rect 15379 745 15413 765
rect 15379 731 15413 745
rect 15379 677 15413 693
rect 15379 659 15413 677
rect 15379 609 15413 621
rect 15379 587 15413 609
rect 15379 541 15413 549
rect 15379 515 15413 541
rect 15379 473 15413 477
rect 15379 443 15413 473
rect 15379 371 15413 405
rect 15837 1595 15871 1629
rect 15837 1527 15871 1557
rect 15837 1523 15871 1527
rect 15837 1459 15871 1485
rect 15837 1451 15871 1459
rect 15837 1391 15871 1413
rect 15837 1379 15871 1391
rect 15837 1323 15871 1341
rect 15837 1307 15871 1323
rect 15837 1255 15871 1269
rect 15837 1235 15871 1255
rect 15837 1187 15871 1197
rect 15837 1163 15871 1187
rect 15837 1119 15871 1125
rect 15837 1091 15871 1119
rect 15837 1051 15871 1053
rect 15837 1019 15871 1051
rect 15837 949 15871 981
rect 15837 947 15871 949
rect 15837 881 15871 909
rect 15837 875 15871 881
rect 15837 813 15871 837
rect 15837 803 15871 813
rect 15837 745 15871 765
rect 15837 731 15871 745
rect 15837 677 15871 693
rect 15837 659 15871 677
rect 15837 609 15871 621
rect 15837 587 15871 609
rect 15837 541 15871 549
rect 15837 515 15871 541
rect 15837 473 15871 477
rect 15837 443 15871 473
rect 15837 371 15871 405
rect 16295 1595 16329 1629
rect 16295 1527 16329 1557
rect 16295 1523 16329 1527
rect 16295 1459 16329 1485
rect 16295 1451 16329 1459
rect 16295 1391 16329 1413
rect 16295 1379 16329 1391
rect 16295 1323 16329 1341
rect 16295 1307 16329 1323
rect 16295 1255 16329 1269
rect 16295 1235 16329 1255
rect 16295 1187 16329 1197
rect 16295 1163 16329 1187
rect 16295 1119 16329 1125
rect 16295 1091 16329 1119
rect 16295 1051 16329 1053
rect 16295 1019 16329 1051
rect 16295 949 16329 981
rect 16295 947 16329 949
rect 16295 881 16329 909
rect 16295 875 16329 881
rect 16295 813 16329 837
rect 16295 803 16329 813
rect 16295 745 16329 765
rect 16295 731 16329 745
rect 16295 677 16329 693
rect 16295 659 16329 677
rect 16295 609 16329 621
rect 16295 587 16329 609
rect 16295 541 16329 549
rect 16295 515 16329 541
rect 16295 473 16329 477
rect 16295 443 16329 473
rect 16295 371 16329 405
rect 16753 1595 16787 1629
rect 16753 1527 16787 1557
rect 16753 1523 16787 1527
rect 16753 1459 16787 1485
rect 16753 1451 16787 1459
rect 16753 1391 16787 1413
rect 16753 1379 16787 1391
rect 16753 1323 16787 1341
rect 16753 1307 16787 1323
rect 16753 1255 16787 1269
rect 16753 1235 16787 1255
rect 16753 1187 16787 1197
rect 16753 1163 16787 1187
rect 16753 1119 16787 1125
rect 16753 1091 16787 1119
rect 16753 1051 16787 1053
rect 16753 1019 16787 1051
rect 16753 949 16787 981
rect 16753 947 16787 949
rect 16753 881 16787 909
rect 16753 875 16787 881
rect 16753 813 16787 837
rect 16753 803 16787 813
rect 16753 745 16787 765
rect 16753 731 16787 745
rect 16753 677 16787 693
rect 16753 659 16787 677
rect 16753 609 16787 621
rect 16753 587 16787 609
rect 16753 541 16787 549
rect 16753 515 16787 541
rect 16753 473 16787 477
rect 16753 443 16787 473
rect 16753 371 16787 405
rect 17211 1595 17245 1629
rect 17211 1527 17245 1557
rect 17211 1523 17245 1527
rect 17211 1459 17245 1485
rect 17211 1451 17245 1459
rect 17211 1391 17245 1413
rect 17211 1379 17245 1391
rect 17211 1323 17245 1341
rect 17211 1307 17245 1323
rect 17211 1255 17245 1269
rect 17211 1235 17245 1255
rect 17211 1187 17245 1197
rect 17211 1163 17245 1187
rect 17211 1119 17245 1125
rect 17211 1091 17245 1119
rect 17211 1051 17245 1053
rect 17211 1019 17245 1051
rect 17211 949 17245 981
rect 17211 947 17245 949
rect 17211 881 17245 909
rect 17211 875 17245 881
rect 17211 813 17245 837
rect 17211 803 17245 813
rect 17211 745 17245 765
rect 17211 731 17245 745
rect 17211 677 17245 693
rect 17211 659 17245 677
rect 17211 609 17245 621
rect 17211 587 17245 609
rect 17211 541 17245 549
rect 17211 515 17245 541
rect 17211 473 17245 477
rect 17211 443 17245 473
rect 17211 371 17245 405
rect 17669 1595 17703 1629
rect 17669 1527 17703 1557
rect 17669 1523 17703 1527
rect 17669 1459 17703 1485
rect 17669 1451 17703 1459
rect 17669 1391 17703 1413
rect 17669 1379 17703 1391
rect 17669 1323 17703 1341
rect 17669 1307 17703 1323
rect 17669 1255 17703 1269
rect 17669 1235 17703 1255
rect 17669 1187 17703 1197
rect 17669 1163 17703 1187
rect 17669 1119 17703 1125
rect 17669 1091 17703 1119
rect 17669 1051 17703 1053
rect 17669 1019 17703 1051
rect 17669 949 17703 981
rect 17669 947 17703 949
rect 17669 881 17703 909
rect 17669 875 17703 881
rect 17669 813 17703 837
rect 17669 803 17703 813
rect 17669 745 17703 765
rect 17669 731 17703 745
rect 17669 677 17703 693
rect 17669 659 17703 677
rect 17669 609 17703 621
rect 17669 587 17703 609
rect 17669 541 17703 549
rect 17669 515 17703 541
rect 17669 473 17703 477
rect 17669 443 17703 473
rect 17669 371 17703 405
rect 18127 1595 18161 1629
rect 18127 1527 18161 1557
rect 18127 1523 18161 1527
rect 18127 1459 18161 1485
rect 18127 1451 18161 1459
rect 18127 1391 18161 1413
rect 18127 1379 18161 1391
rect 18127 1323 18161 1341
rect 18127 1307 18161 1323
rect 18127 1255 18161 1269
rect 18127 1235 18161 1255
rect 18127 1187 18161 1197
rect 18127 1163 18161 1187
rect 18127 1119 18161 1125
rect 18127 1091 18161 1119
rect 18127 1051 18161 1053
rect 18127 1019 18161 1051
rect 18127 949 18161 981
rect 18127 947 18161 949
rect 18127 881 18161 909
rect 18127 875 18161 881
rect 18127 813 18161 837
rect 18127 803 18161 813
rect 18127 745 18161 765
rect 18127 731 18161 745
rect 18127 677 18161 693
rect 18127 659 18161 677
rect 18127 609 18161 621
rect 18127 587 18161 609
rect 18127 541 18161 549
rect 18127 515 18161 541
rect 18127 473 18161 477
rect 18127 443 18161 473
rect 18127 371 18161 405
rect 18585 1595 18619 1629
rect 18585 1527 18619 1557
rect 18585 1523 18619 1527
rect 18585 1459 18619 1485
rect 18585 1451 18619 1459
rect 18585 1391 18619 1413
rect 18585 1379 18619 1391
rect 18585 1323 18619 1341
rect 18585 1307 18619 1323
rect 18585 1255 18619 1269
rect 18585 1235 18619 1255
rect 18585 1187 18619 1197
rect 18585 1163 18619 1187
rect 18585 1119 18619 1125
rect 18585 1091 18619 1119
rect 18585 1051 18619 1053
rect 18585 1019 18619 1051
rect 18585 949 18619 981
rect 18585 947 18619 949
rect 18585 881 18619 909
rect 18585 875 18619 881
rect 18585 813 18619 837
rect 18585 803 18619 813
rect 18585 745 18619 765
rect 18585 731 18619 745
rect 18585 677 18619 693
rect 18585 659 18619 677
rect 18585 609 18619 621
rect 18585 587 18619 609
rect 18585 541 18619 549
rect 18585 515 18619 541
rect 18585 473 18619 477
rect 18585 443 18619 473
rect 18585 371 18619 405
rect 19043 1595 19077 1629
rect 19043 1527 19077 1557
rect 19043 1523 19077 1527
rect 19043 1459 19077 1485
rect 19043 1451 19077 1459
rect 19043 1391 19077 1413
rect 19043 1379 19077 1391
rect 19043 1323 19077 1341
rect 19043 1307 19077 1323
rect 19043 1255 19077 1269
rect 19043 1235 19077 1255
rect 19043 1187 19077 1197
rect 19043 1163 19077 1187
rect 19043 1119 19077 1125
rect 19043 1091 19077 1119
rect 19043 1051 19077 1053
rect 19043 1019 19077 1051
rect 19043 949 19077 981
rect 19043 947 19077 949
rect 19043 881 19077 909
rect 19043 875 19077 881
rect 19043 813 19077 837
rect 19043 803 19077 813
rect 19043 745 19077 765
rect 19043 731 19077 745
rect 19043 677 19077 693
rect 19043 659 19077 677
rect 19043 609 19077 621
rect 19043 587 19077 609
rect 19043 541 19077 549
rect 19043 515 19077 541
rect 19043 473 19077 477
rect 19043 443 19077 473
rect 19043 371 19077 405
rect 19501 1595 19535 1629
rect 19501 1527 19535 1557
rect 19501 1523 19535 1527
rect 19501 1459 19535 1485
rect 19501 1451 19535 1459
rect 19501 1391 19535 1413
rect 19501 1379 19535 1391
rect 19501 1323 19535 1341
rect 19501 1307 19535 1323
rect 19501 1255 19535 1269
rect 19501 1235 19535 1255
rect 19501 1187 19535 1197
rect 19501 1163 19535 1187
rect 19501 1119 19535 1125
rect 19501 1091 19535 1119
rect 19501 1051 19535 1053
rect 19501 1019 19535 1051
rect 19501 949 19535 981
rect 19501 947 19535 949
rect 19501 881 19535 909
rect 19501 875 19535 881
rect 19501 813 19535 837
rect 19501 803 19535 813
rect 19501 745 19535 765
rect 19501 731 19535 745
rect 19501 677 19535 693
rect 19501 659 19535 677
rect 19501 609 19535 621
rect 19501 587 19535 609
rect 19501 541 19535 549
rect 19501 515 19535 541
rect 19501 473 19535 477
rect 19501 443 19535 473
rect 19501 371 19535 405
rect 19959 1595 19993 1629
rect 19959 1527 19993 1557
rect 19959 1523 19993 1527
rect 19959 1459 19993 1485
rect 19959 1451 19993 1459
rect 19959 1391 19993 1413
rect 19959 1379 19993 1391
rect 19959 1323 19993 1341
rect 19959 1307 19993 1323
rect 19959 1255 19993 1269
rect 19959 1235 19993 1255
rect 19959 1187 19993 1197
rect 19959 1163 19993 1187
rect 19959 1119 19993 1125
rect 19959 1091 19993 1119
rect 19959 1051 19993 1053
rect 19959 1019 19993 1051
rect 19959 949 19993 981
rect 19959 947 19993 949
rect 19959 881 19993 909
rect 19959 875 19993 881
rect 19959 813 19993 837
rect 19959 803 19993 813
rect 19959 745 19993 765
rect 19959 731 19993 745
rect 19959 677 19993 693
rect 19959 659 19993 677
rect 19959 609 19993 621
rect 19959 587 19993 609
rect 19959 541 19993 549
rect 19959 515 19993 541
rect 19959 473 19993 477
rect 19959 443 19993 473
rect 19959 371 19993 405
rect 20417 1595 20451 1629
rect 20417 1527 20451 1557
rect 20417 1523 20451 1527
rect 20417 1459 20451 1485
rect 20417 1451 20451 1459
rect 20417 1391 20451 1413
rect 20417 1379 20451 1391
rect 20417 1323 20451 1341
rect 20417 1307 20451 1323
rect 20417 1255 20451 1269
rect 20417 1235 20451 1255
rect 20417 1187 20451 1197
rect 20417 1163 20451 1187
rect 20417 1119 20451 1125
rect 20417 1091 20451 1119
rect 20417 1051 20451 1053
rect 20417 1019 20451 1051
rect 20417 949 20451 981
rect 20417 947 20451 949
rect 20417 881 20451 909
rect 20417 875 20451 881
rect 20417 813 20451 837
rect 20417 803 20451 813
rect 20417 745 20451 765
rect 20417 731 20451 745
rect 20417 677 20451 693
rect 20417 659 20451 677
rect 20417 609 20451 621
rect 20417 587 20451 609
rect 20417 541 20451 549
rect 20417 515 20451 541
rect 20417 473 20451 477
rect 20417 443 20451 473
rect 20417 371 20451 405
rect 20875 1595 20909 1629
rect 20875 1527 20909 1557
rect 20875 1523 20909 1527
rect 20875 1459 20909 1485
rect 20875 1451 20909 1459
rect 20875 1391 20909 1413
rect 20875 1379 20909 1391
rect 20875 1323 20909 1341
rect 20875 1307 20909 1323
rect 20875 1255 20909 1269
rect 20875 1235 20909 1255
rect 20875 1187 20909 1197
rect 20875 1163 20909 1187
rect 20875 1119 20909 1125
rect 20875 1091 20909 1119
rect 20875 1051 20909 1053
rect 20875 1019 20909 1051
rect 20875 949 20909 981
rect 20875 947 20909 949
rect 20875 881 20909 909
rect 20875 875 20909 881
rect 20875 813 20909 837
rect 20875 803 20909 813
rect 20875 745 20909 765
rect 20875 731 20909 745
rect 20875 677 20909 693
rect 20875 659 20909 677
rect 20875 609 20909 621
rect 20875 587 20909 609
rect 20875 541 20909 549
rect 20875 515 20909 541
rect 20875 473 20909 477
rect 20875 443 20909 473
rect 20875 371 20909 405
rect 21333 1595 21367 1629
rect 21333 1527 21367 1557
rect 21333 1523 21367 1527
rect 21333 1459 21367 1485
rect 21333 1451 21367 1459
rect 21333 1391 21367 1413
rect 21333 1379 21367 1391
rect 21333 1323 21367 1341
rect 21333 1307 21367 1323
rect 21333 1255 21367 1269
rect 21333 1235 21367 1255
rect 21333 1187 21367 1197
rect 21333 1163 21367 1187
rect 21333 1119 21367 1125
rect 21333 1091 21367 1119
rect 21333 1051 21367 1053
rect 21333 1019 21367 1051
rect 21333 949 21367 981
rect 21333 947 21367 949
rect 21333 881 21367 909
rect 21333 875 21367 881
rect 21333 813 21367 837
rect 21333 803 21367 813
rect 21333 745 21367 765
rect 21333 731 21367 745
rect 21333 677 21367 693
rect 21333 659 21367 677
rect 21333 609 21367 621
rect 21333 587 21367 609
rect 21333 541 21367 549
rect 21333 515 21367 541
rect 21333 473 21367 477
rect 21333 443 21367 473
rect 21333 371 21367 405
rect 21791 1595 21825 1629
rect 21791 1527 21825 1557
rect 21791 1523 21825 1527
rect 21791 1459 21825 1485
rect 21791 1451 21825 1459
rect 21791 1391 21825 1413
rect 21791 1379 21825 1391
rect 21791 1323 21825 1341
rect 21791 1307 21825 1323
rect 21791 1255 21825 1269
rect 21791 1235 21825 1255
rect 21791 1187 21825 1197
rect 21791 1163 21825 1187
rect 21791 1119 21825 1125
rect 21791 1091 21825 1119
rect 21791 1051 21825 1053
rect 21791 1019 21825 1051
rect 21791 949 21825 981
rect 21791 947 21825 949
rect 21791 881 21825 909
rect 21791 875 21825 881
rect 21791 813 21825 837
rect 21791 803 21825 813
rect 21791 745 21825 765
rect 21791 731 21825 745
rect 21791 677 21825 693
rect 21791 659 21825 677
rect 21791 609 21825 621
rect 21791 587 21825 609
rect 21791 541 21825 549
rect 21791 515 21825 541
rect 21791 473 21825 477
rect 21791 443 21825 473
rect 21791 371 21825 405
rect 22249 1595 22283 1629
rect 22249 1527 22283 1557
rect 22249 1523 22283 1527
rect 22249 1459 22283 1485
rect 22249 1451 22283 1459
rect 22249 1391 22283 1413
rect 22249 1379 22283 1391
rect 22249 1323 22283 1341
rect 22249 1307 22283 1323
rect 22249 1255 22283 1269
rect 22249 1235 22283 1255
rect 22249 1187 22283 1197
rect 22249 1163 22283 1187
rect 22249 1119 22283 1125
rect 22249 1091 22283 1119
rect 22249 1051 22283 1053
rect 22249 1019 22283 1051
rect 22249 949 22283 981
rect 22249 947 22283 949
rect 22249 881 22283 909
rect 22249 875 22283 881
rect 22249 813 22283 837
rect 22249 803 22283 813
rect 22249 745 22283 765
rect 22249 731 22283 745
rect 22249 677 22283 693
rect 22249 659 22283 677
rect 22249 609 22283 621
rect 22249 587 22283 609
rect 22249 541 22283 549
rect 22249 515 22283 541
rect 22249 473 22283 477
rect 22249 443 22283 473
rect 22249 371 22283 405
rect 22707 1595 22741 1629
rect 22707 1527 22741 1557
rect 22707 1523 22741 1527
rect 22707 1459 22741 1485
rect 22707 1451 22741 1459
rect 22707 1391 22741 1413
rect 22707 1379 22741 1391
rect 22707 1323 22741 1341
rect 22707 1307 22741 1323
rect 22707 1255 22741 1269
rect 22707 1235 22741 1255
rect 22707 1187 22741 1197
rect 22707 1163 22741 1187
rect 22707 1119 22741 1125
rect 22707 1091 22741 1119
rect 22707 1051 22741 1053
rect 22707 1019 22741 1051
rect 22707 949 22741 981
rect 22707 947 22741 949
rect 22707 881 22741 909
rect 22707 875 22741 881
rect 22707 813 22741 837
rect 22707 803 22741 813
rect 22707 745 22741 765
rect 22707 731 22741 745
rect 22707 677 22741 693
rect 22707 659 22741 677
rect 22707 609 22741 621
rect 22707 587 22741 609
rect 22707 541 22741 549
rect 22707 515 22741 541
rect 22707 473 22741 477
rect 22707 443 22741 473
rect 22707 371 22741 405
rect 23165 1595 23199 1629
rect 23165 1527 23199 1557
rect 23165 1523 23199 1527
rect 23165 1459 23199 1485
rect 23165 1451 23199 1459
rect 23165 1391 23199 1413
rect 23165 1379 23199 1391
rect 23165 1323 23199 1341
rect 23165 1307 23199 1323
rect 23165 1255 23199 1269
rect 23165 1235 23199 1255
rect 23165 1187 23199 1197
rect 23165 1163 23199 1187
rect 23165 1119 23199 1125
rect 23165 1091 23199 1119
rect 23165 1051 23199 1053
rect 23165 1019 23199 1051
rect 23165 949 23199 981
rect 23165 947 23199 949
rect 23165 881 23199 909
rect 23165 875 23199 881
rect 23165 813 23199 837
rect 23165 803 23199 813
rect 23165 745 23199 765
rect 23165 731 23199 745
rect 23165 677 23199 693
rect 23165 659 23199 677
rect 23165 609 23199 621
rect 23165 587 23199 609
rect 23165 541 23199 549
rect 23165 515 23199 541
rect 23165 473 23199 477
rect 23165 443 23199 473
rect 23165 371 23199 405
rect 23623 1595 23657 1629
rect 23623 1527 23657 1557
rect 23623 1523 23657 1527
rect 23623 1459 23657 1485
rect 23623 1451 23657 1459
rect 23623 1391 23657 1413
rect 23623 1379 23657 1391
rect 23623 1323 23657 1341
rect 23623 1307 23657 1323
rect 23623 1255 23657 1269
rect 23623 1235 23657 1255
rect 23623 1187 23657 1197
rect 23623 1163 23657 1187
rect 23623 1119 23657 1125
rect 23623 1091 23657 1119
rect 23623 1051 23657 1053
rect 23623 1019 23657 1051
rect 23623 949 23657 981
rect 23623 947 23657 949
rect 23623 881 23657 909
rect 23623 875 23657 881
rect 23623 813 23657 837
rect 23623 803 23657 813
rect 23623 745 23657 765
rect 23623 731 23657 745
rect 23623 677 23657 693
rect 23623 659 23657 677
rect 23623 609 23657 621
rect 23623 587 23657 609
rect 23623 541 23657 549
rect 23623 515 23657 541
rect 23623 473 23657 477
rect 23623 443 23657 473
rect 23623 371 23657 405
rect 24081 1595 24115 1629
rect 24081 1527 24115 1557
rect 24081 1523 24115 1527
rect 24081 1459 24115 1485
rect 24081 1451 24115 1459
rect 24081 1391 24115 1413
rect 24081 1379 24115 1391
rect 24081 1323 24115 1341
rect 24081 1307 24115 1323
rect 24081 1255 24115 1269
rect 24081 1235 24115 1255
rect 24081 1187 24115 1197
rect 24081 1163 24115 1187
rect 24081 1119 24115 1125
rect 24081 1091 24115 1119
rect 24081 1051 24115 1053
rect 24081 1019 24115 1051
rect 24081 949 24115 981
rect 24081 947 24115 949
rect 24081 881 24115 909
rect 24081 875 24115 881
rect 24081 813 24115 837
rect 24081 803 24115 813
rect 24081 745 24115 765
rect 24081 731 24115 745
rect 24081 677 24115 693
rect 24081 659 24115 677
rect 24081 609 24115 621
rect 24081 587 24115 609
rect 24081 541 24115 549
rect 24081 515 24115 541
rect 24081 473 24115 477
rect 24081 443 24115 473
rect 24081 371 24115 405
rect 24539 1595 24573 1629
rect 24539 1527 24573 1557
rect 24539 1523 24573 1527
rect 24539 1459 24573 1485
rect 24539 1451 24573 1459
rect 24539 1391 24573 1413
rect 24539 1379 24573 1391
rect 24539 1323 24573 1341
rect 24539 1307 24573 1323
rect 24539 1255 24573 1269
rect 24539 1235 24573 1255
rect 24539 1187 24573 1197
rect 24539 1163 24573 1187
rect 24539 1119 24573 1125
rect 24539 1091 24573 1119
rect 24539 1051 24573 1053
rect 24539 1019 24573 1051
rect 24539 949 24573 981
rect 24539 947 24573 949
rect 24539 881 24573 909
rect 24539 875 24573 881
rect 24539 813 24573 837
rect 24539 803 24573 813
rect 24539 745 24573 765
rect 24539 731 24573 745
rect 24539 677 24573 693
rect 24539 659 24573 677
rect 24539 609 24573 621
rect 24539 587 24573 609
rect 24539 541 24573 549
rect 24539 515 24573 541
rect 24539 473 24573 477
rect 24539 443 24573 473
rect 24539 371 24573 405
rect 24997 1595 25031 1629
rect 24997 1527 25031 1557
rect 24997 1523 25031 1527
rect 24997 1459 25031 1485
rect 24997 1451 25031 1459
rect 24997 1391 25031 1413
rect 24997 1379 25031 1391
rect 24997 1323 25031 1341
rect 24997 1307 25031 1323
rect 24997 1255 25031 1269
rect 24997 1235 25031 1255
rect 24997 1187 25031 1197
rect 24997 1163 25031 1187
rect 24997 1119 25031 1125
rect 24997 1091 25031 1119
rect 24997 1051 25031 1053
rect 24997 1019 25031 1051
rect 24997 949 25031 981
rect 24997 947 25031 949
rect 24997 881 25031 909
rect 24997 875 25031 881
rect 24997 813 25031 837
rect 24997 803 25031 813
rect 24997 745 25031 765
rect 24997 731 25031 745
rect 24997 677 25031 693
rect 24997 659 25031 677
rect 24997 609 25031 621
rect 24997 587 25031 609
rect 24997 541 25031 549
rect 24997 515 25031 541
rect 24997 473 25031 477
rect 24997 443 25031 473
rect 24997 371 25031 405
rect 25455 1595 25489 1629
rect 25455 1527 25489 1557
rect 25455 1523 25489 1527
rect 25455 1459 25489 1485
rect 25455 1451 25489 1459
rect 25455 1391 25489 1413
rect 25455 1379 25489 1391
rect 25455 1323 25489 1341
rect 25455 1307 25489 1323
rect 25455 1255 25489 1269
rect 25455 1235 25489 1255
rect 25455 1187 25489 1197
rect 25455 1163 25489 1187
rect 25455 1119 25489 1125
rect 25455 1091 25489 1119
rect 25455 1051 25489 1053
rect 25455 1019 25489 1051
rect 25455 949 25489 981
rect 25455 947 25489 949
rect 25455 881 25489 909
rect 25455 875 25489 881
rect 25455 813 25489 837
rect 25455 803 25489 813
rect 25455 745 25489 765
rect 25455 731 25489 745
rect 25455 677 25489 693
rect 25455 659 25489 677
rect 25455 609 25489 621
rect 25455 587 25489 609
rect 25455 541 25489 549
rect 25455 515 25489 541
rect 25455 473 25489 477
rect 25455 443 25489 473
rect 25455 371 25489 405
rect 25913 1595 25947 1629
rect 25913 1527 25947 1557
rect 25913 1523 25947 1527
rect 25913 1459 25947 1485
rect 25913 1451 25947 1459
rect 25913 1391 25947 1413
rect 25913 1379 25947 1391
rect 25913 1323 25947 1341
rect 25913 1307 25947 1323
rect 25913 1255 25947 1269
rect 25913 1235 25947 1255
rect 25913 1187 25947 1197
rect 25913 1163 25947 1187
rect 25913 1119 25947 1125
rect 25913 1091 25947 1119
rect 25913 1051 25947 1053
rect 25913 1019 25947 1051
rect 25913 949 25947 981
rect 25913 947 25947 949
rect 25913 881 25947 909
rect 25913 875 25947 881
rect 25913 813 25947 837
rect 25913 803 25947 813
rect 25913 745 25947 765
rect 25913 731 25947 745
rect 25913 677 25947 693
rect 25913 659 25947 677
rect 25913 609 25947 621
rect 25913 587 25947 609
rect 25913 541 25947 549
rect 25913 515 25947 541
rect 25913 473 25947 477
rect 25913 443 25947 473
rect 25913 371 25947 405
rect 26371 1595 26405 1629
rect 26371 1527 26405 1557
rect 26371 1523 26405 1527
rect 26371 1459 26405 1485
rect 26371 1451 26405 1459
rect 26371 1391 26405 1413
rect 26371 1379 26405 1391
rect 26371 1323 26405 1341
rect 26371 1307 26405 1323
rect 26371 1255 26405 1269
rect 26371 1235 26405 1255
rect 26371 1187 26405 1197
rect 26371 1163 26405 1187
rect 26371 1119 26405 1125
rect 26371 1091 26405 1119
rect 26371 1051 26405 1053
rect 26371 1019 26405 1051
rect 26371 949 26405 981
rect 26371 947 26405 949
rect 26371 881 26405 909
rect 26371 875 26405 881
rect 26371 813 26405 837
rect 26371 803 26405 813
rect 26371 745 26405 765
rect 26371 731 26405 745
rect 26371 677 26405 693
rect 26371 659 26405 677
rect 26371 609 26405 621
rect 26371 587 26405 609
rect 26371 541 26405 549
rect 26371 515 26405 541
rect 26371 473 26405 477
rect 26371 443 26405 473
rect 26371 371 26405 405
rect 26829 1595 26863 1629
rect 26829 1527 26863 1557
rect 26829 1523 26863 1527
rect 26829 1459 26863 1485
rect 26829 1451 26863 1459
rect 26829 1391 26863 1413
rect 26829 1379 26863 1391
rect 26829 1323 26863 1341
rect 26829 1307 26863 1323
rect 26829 1255 26863 1269
rect 26829 1235 26863 1255
rect 26829 1187 26863 1197
rect 26829 1163 26863 1187
rect 26829 1119 26863 1125
rect 26829 1091 26863 1119
rect 26829 1051 26863 1053
rect 26829 1019 26863 1051
rect 26829 949 26863 981
rect 26829 947 26863 949
rect 26829 881 26863 909
rect 26829 875 26863 881
rect 26829 813 26863 837
rect 26829 803 26863 813
rect 26829 745 26863 765
rect 26829 731 26863 745
rect 26829 677 26863 693
rect 26829 659 26863 677
rect 26829 609 26863 621
rect 26829 587 26863 609
rect 26829 541 26863 549
rect 26829 515 26863 541
rect 26829 473 26863 477
rect 26829 443 26863 473
rect 26829 371 26863 405
rect 27287 1595 27321 1629
rect 27287 1527 27321 1557
rect 27287 1523 27321 1527
rect 27287 1459 27321 1485
rect 27287 1451 27321 1459
rect 27287 1391 27321 1413
rect 27287 1379 27321 1391
rect 27287 1323 27321 1341
rect 27287 1307 27321 1323
rect 27287 1255 27321 1269
rect 27287 1235 27321 1255
rect 27287 1187 27321 1197
rect 27287 1163 27321 1187
rect 27287 1119 27321 1125
rect 27287 1091 27321 1119
rect 27287 1051 27321 1053
rect 27287 1019 27321 1051
rect 27287 949 27321 981
rect 27287 947 27321 949
rect 27287 881 27321 909
rect 27287 875 27321 881
rect 27287 813 27321 837
rect 27287 803 27321 813
rect 27287 745 27321 765
rect 27287 731 27321 745
rect 27287 677 27321 693
rect 27287 659 27321 677
rect 27287 609 27321 621
rect 27287 587 27321 609
rect 27287 541 27321 549
rect 27287 515 27321 541
rect 27287 473 27321 477
rect 27287 443 27321 473
rect 27287 371 27321 405
rect 27745 1595 27779 1629
rect 27745 1527 27779 1557
rect 27745 1523 27779 1527
rect 27745 1459 27779 1485
rect 27745 1451 27779 1459
rect 27745 1391 27779 1413
rect 27745 1379 27779 1391
rect 27745 1323 27779 1341
rect 27745 1307 27779 1323
rect 27745 1255 27779 1269
rect 27745 1235 27779 1255
rect 27745 1187 27779 1197
rect 27745 1163 27779 1187
rect 27745 1119 27779 1125
rect 27745 1091 27779 1119
rect 27745 1051 27779 1053
rect 27745 1019 27779 1051
rect 27745 949 27779 981
rect 27745 947 27779 949
rect 27745 881 27779 909
rect 27745 875 27779 881
rect 27745 813 27779 837
rect 27745 803 27779 813
rect 27745 745 27779 765
rect 27745 731 27779 745
rect 27745 677 27779 693
rect 27745 659 27779 677
rect 27745 609 27779 621
rect 27745 587 27779 609
rect 27745 541 27779 549
rect 27745 515 27779 541
rect 27745 473 27779 477
rect 27745 443 27779 473
rect 27745 371 27779 405
rect 401 -17 435 17
rect 801 -17 835 17
rect 1201 -17 1235 17
rect 1601 -17 1635 17
rect 2001 -17 2035 17
rect 2401 -17 2435 17
rect 2801 -17 2835 17
rect 3201 -17 3235 17
rect 3601 -17 3635 17
rect 4001 -17 4035 17
rect 4401 -17 4435 17
rect 4801 -17 4835 17
rect 5201 -17 5235 17
rect 5601 -17 5635 17
rect 6001 -17 6035 17
rect 6401 -17 6435 17
rect 6801 -17 6835 17
rect 7201 -17 7235 17
rect 7601 -17 7635 17
rect 8001 -17 8035 17
rect 8401 -17 8435 17
rect 8801 -17 8835 17
rect 9201 -17 9235 17
rect 9601 -17 9635 17
rect 10001 -17 10035 17
rect 10401 -17 10435 17
rect 10801 -17 10835 17
rect 11201 -17 11235 17
rect 11601 -17 11635 17
rect 12001 -17 12035 17
rect 12401 -17 12435 17
rect 12801 -17 12835 17
rect 13201 -17 13235 17
rect 13601 -17 13635 17
rect 14001 -17 14035 17
rect 14401 -17 14435 17
rect 14801 -17 14835 17
rect 15201 -17 15235 17
rect 15601 -17 15635 17
rect 16001 -17 16035 17
rect 16401 -17 16435 17
rect 16801 -17 16835 17
rect 17201 -17 17235 17
rect 17601 -17 17635 17
rect 18001 -17 18035 17
rect 18401 -17 18435 17
rect 18801 -17 18835 17
rect 19201 -17 19235 17
rect 19601 -17 19635 17
rect 20001 -17 20035 17
rect 20401 -17 20435 17
rect 20801 -17 20835 17
rect 21201 -17 21235 17
rect 21601 -17 21635 17
rect 22001 -17 22035 17
rect 22401 -17 22435 17
rect 22801 -17 22835 17
rect 23201 -17 23235 17
rect 23601 -17 23635 17
rect 24001 -17 24035 17
rect 24401 -17 24435 17
rect 24801 -17 24835 17
rect 25201 -17 25235 17
rect 25601 -17 25635 17
rect 26001 -17 26035 17
rect 26401 -17 26435 17
rect 26801 -17 26835 17
rect 27201 -17 27235 17
rect 27601 -17 27635 17
<< metal1 >>
rect 120 1897 27826 1940
rect 120 1863 401 1897
rect 435 1863 801 1897
rect 835 1863 1201 1897
rect 1235 1863 1601 1897
rect 1635 1863 2001 1897
rect 2035 1863 2401 1897
rect 2435 1863 2801 1897
rect 2835 1863 3201 1897
rect 3235 1863 3601 1897
rect 3635 1863 4001 1897
rect 4035 1863 4401 1897
rect 4435 1863 4801 1897
rect 4835 1863 5201 1897
rect 5235 1863 5601 1897
rect 5635 1863 6001 1897
rect 6035 1863 6401 1897
rect 6435 1863 6801 1897
rect 6835 1863 7201 1897
rect 7235 1863 7601 1897
rect 7635 1863 8001 1897
rect 8035 1863 8401 1897
rect 8435 1863 8801 1897
rect 8835 1863 9201 1897
rect 9235 1863 9601 1897
rect 9635 1863 10001 1897
rect 10035 1863 10401 1897
rect 10435 1863 10801 1897
rect 10835 1863 11201 1897
rect 11235 1863 11601 1897
rect 11635 1863 12001 1897
rect 12035 1863 12401 1897
rect 12435 1863 12801 1897
rect 12835 1863 13201 1897
rect 13235 1863 13601 1897
rect 13635 1863 14001 1897
rect 14035 1863 14401 1897
rect 14435 1863 14801 1897
rect 14835 1863 15201 1897
rect 15235 1863 15601 1897
rect 15635 1863 16001 1897
rect 16035 1863 16401 1897
rect 16435 1863 16801 1897
rect 16835 1863 17201 1897
rect 17235 1863 17601 1897
rect 17635 1863 18001 1897
rect 18035 1863 18401 1897
rect 18435 1863 18801 1897
rect 18835 1863 19201 1897
rect 19235 1863 19601 1897
rect 19635 1863 20001 1897
rect 20035 1863 20401 1897
rect 20435 1863 20801 1897
rect 20835 1863 21201 1897
rect 21235 1863 21601 1897
rect 21635 1863 22001 1897
rect 22035 1863 22401 1897
rect 22435 1863 22801 1897
rect 22835 1863 23201 1897
rect 23235 1863 23601 1897
rect 23635 1863 24001 1897
rect 24035 1863 24401 1897
rect 24435 1863 24801 1897
rect 24835 1863 25201 1897
rect 25235 1863 25601 1897
rect 25635 1863 26001 1897
rect 26035 1863 26401 1897
rect 26435 1863 26801 1897
rect 26835 1863 27201 1897
rect 27235 1863 27601 1897
rect 27635 1863 27826 1897
rect 120 1820 27826 1863
rect 259 1629 305 1645
rect 259 1595 265 1629
rect 299 1595 305 1629
rect 259 1557 305 1595
rect 259 1523 265 1557
rect 299 1523 305 1557
rect 259 1485 305 1523
rect 259 1451 265 1485
rect 299 1451 305 1485
rect 259 1413 305 1451
rect 259 1379 265 1413
rect 299 1379 305 1413
rect 259 1341 305 1379
rect 259 1307 265 1341
rect 299 1307 305 1341
rect 259 1269 305 1307
rect 259 1235 265 1269
rect 299 1235 305 1269
rect 259 1197 305 1235
rect 259 1163 265 1197
rect 299 1163 305 1197
rect 259 1125 305 1163
rect 259 1091 265 1125
rect 299 1091 305 1125
rect 259 1053 305 1091
rect 259 1019 265 1053
rect 299 1019 305 1053
rect 259 981 305 1019
rect 259 947 265 981
rect 299 947 305 981
rect 259 909 305 947
rect 259 875 265 909
rect 299 875 305 909
rect 259 837 305 875
rect 259 803 265 837
rect 299 803 305 837
rect 259 765 305 803
rect 259 731 265 765
rect 299 731 305 765
rect 259 693 305 731
rect 259 659 265 693
rect 299 659 305 693
rect 259 621 305 659
rect 259 587 265 621
rect 299 587 305 621
rect 259 549 305 587
rect 259 515 265 549
rect 299 515 305 549
rect 259 477 305 515
rect 259 443 265 477
rect 299 443 305 477
rect 259 405 305 443
rect 259 371 265 405
rect 299 371 305 405
rect 259 355 305 371
rect 717 1629 763 1645
rect 717 1595 723 1629
rect 757 1595 763 1629
rect 717 1557 763 1595
rect 717 1523 723 1557
rect 757 1523 763 1557
rect 717 1485 763 1523
rect 717 1451 723 1485
rect 757 1451 763 1485
rect 717 1413 763 1451
rect 717 1379 723 1413
rect 757 1379 763 1413
rect 717 1341 763 1379
rect 717 1307 723 1341
rect 757 1307 763 1341
rect 717 1269 763 1307
rect 717 1235 723 1269
rect 757 1235 763 1269
rect 717 1197 763 1235
rect 717 1163 723 1197
rect 757 1163 763 1197
rect 717 1125 763 1163
rect 717 1091 723 1125
rect 757 1091 763 1125
rect 717 1053 763 1091
rect 717 1019 723 1053
rect 757 1019 763 1053
rect 717 981 763 1019
rect 717 947 723 981
rect 757 947 763 981
rect 717 909 763 947
rect 717 875 723 909
rect 757 875 763 909
rect 717 837 763 875
rect 717 803 723 837
rect 757 803 763 837
rect 717 765 763 803
rect 717 731 723 765
rect 757 731 763 765
rect 717 693 763 731
rect 717 659 723 693
rect 757 659 763 693
rect 717 621 763 659
rect 717 587 723 621
rect 757 587 763 621
rect 717 549 763 587
rect 717 515 723 549
rect 757 515 763 549
rect 717 477 763 515
rect 717 443 723 477
rect 757 443 763 477
rect 717 405 763 443
rect 717 371 723 405
rect 757 371 763 405
rect 717 355 763 371
rect 1175 1629 1221 1645
rect 1175 1595 1181 1629
rect 1215 1595 1221 1629
rect 1175 1557 1221 1595
rect 1175 1523 1181 1557
rect 1215 1523 1221 1557
rect 1175 1485 1221 1523
rect 1175 1451 1181 1485
rect 1215 1451 1221 1485
rect 1175 1413 1221 1451
rect 1175 1379 1181 1413
rect 1215 1379 1221 1413
rect 1175 1341 1221 1379
rect 1175 1307 1181 1341
rect 1215 1307 1221 1341
rect 1175 1269 1221 1307
rect 1175 1235 1181 1269
rect 1215 1235 1221 1269
rect 1175 1197 1221 1235
rect 1175 1163 1181 1197
rect 1215 1163 1221 1197
rect 1175 1125 1221 1163
rect 1175 1091 1181 1125
rect 1215 1091 1221 1125
rect 1175 1053 1221 1091
rect 1175 1019 1181 1053
rect 1215 1019 1221 1053
rect 1175 981 1221 1019
rect 1175 947 1181 981
rect 1215 947 1221 981
rect 1175 909 1221 947
rect 1175 875 1181 909
rect 1215 875 1221 909
rect 1175 837 1221 875
rect 1175 803 1181 837
rect 1215 803 1221 837
rect 1175 765 1221 803
rect 1175 731 1181 765
rect 1215 731 1221 765
rect 1175 693 1221 731
rect 1175 659 1181 693
rect 1215 659 1221 693
rect 1175 621 1221 659
rect 1175 587 1181 621
rect 1215 587 1221 621
rect 1175 549 1221 587
rect 1175 515 1181 549
rect 1215 515 1221 549
rect 1175 477 1221 515
rect 1175 443 1181 477
rect 1215 443 1221 477
rect 1175 405 1221 443
rect 1175 371 1181 405
rect 1215 371 1221 405
rect 1175 355 1221 371
rect 1633 1629 1679 1645
rect 1633 1595 1639 1629
rect 1673 1595 1679 1629
rect 1633 1557 1679 1595
rect 1633 1523 1639 1557
rect 1673 1523 1679 1557
rect 1633 1485 1679 1523
rect 1633 1451 1639 1485
rect 1673 1451 1679 1485
rect 1633 1413 1679 1451
rect 1633 1379 1639 1413
rect 1673 1379 1679 1413
rect 1633 1341 1679 1379
rect 1633 1307 1639 1341
rect 1673 1307 1679 1341
rect 1633 1269 1679 1307
rect 1633 1235 1639 1269
rect 1673 1235 1679 1269
rect 1633 1197 1679 1235
rect 1633 1163 1639 1197
rect 1673 1163 1679 1197
rect 1633 1125 1679 1163
rect 1633 1091 1639 1125
rect 1673 1091 1679 1125
rect 1633 1053 1679 1091
rect 1633 1019 1639 1053
rect 1673 1019 1679 1053
rect 1633 981 1679 1019
rect 1633 947 1639 981
rect 1673 947 1679 981
rect 1633 909 1679 947
rect 1633 875 1639 909
rect 1673 875 1679 909
rect 1633 837 1679 875
rect 1633 803 1639 837
rect 1673 803 1679 837
rect 1633 765 1679 803
rect 1633 731 1639 765
rect 1673 731 1679 765
rect 1633 693 1679 731
rect 1633 659 1639 693
rect 1673 659 1679 693
rect 1633 621 1679 659
rect 1633 587 1639 621
rect 1673 587 1679 621
rect 1633 549 1679 587
rect 1633 515 1639 549
rect 1673 515 1679 549
rect 1633 477 1679 515
rect 1633 443 1639 477
rect 1673 443 1679 477
rect 1633 405 1679 443
rect 1633 371 1639 405
rect 1673 371 1679 405
rect 1633 355 1679 371
rect 2091 1629 2137 1645
rect 2091 1595 2097 1629
rect 2131 1595 2137 1629
rect 2091 1557 2137 1595
rect 2091 1523 2097 1557
rect 2131 1523 2137 1557
rect 2091 1485 2137 1523
rect 2091 1451 2097 1485
rect 2131 1451 2137 1485
rect 2091 1413 2137 1451
rect 2091 1379 2097 1413
rect 2131 1379 2137 1413
rect 2091 1341 2137 1379
rect 2091 1307 2097 1341
rect 2131 1307 2137 1341
rect 2091 1269 2137 1307
rect 2091 1235 2097 1269
rect 2131 1235 2137 1269
rect 2091 1197 2137 1235
rect 2091 1163 2097 1197
rect 2131 1163 2137 1197
rect 2091 1125 2137 1163
rect 2091 1091 2097 1125
rect 2131 1091 2137 1125
rect 2091 1053 2137 1091
rect 2091 1019 2097 1053
rect 2131 1019 2137 1053
rect 2091 981 2137 1019
rect 2091 947 2097 981
rect 2131 947 2137 981
rect 2091 909 2137 947
rect 2091 875 2097 909
rect 2131 875 2137 909
rect 2091 837 2137 875
rect 2091 803 2097 837
rect 2131 803 2137 837
rect 2091 765 2137 803
rect 2091 731 2097 765
rect 2131 731 2137 765
rect 2091 693 2137 731
rect 2091 659 2097 693
rect 2131 659 2137 693
rect 2091 621 2137 659
rect 2091 587 2097 621
rect 2131 587 2137 621
rect 2091 549 2137 587
rect 2091 515 2097 549
rect 2131 515 2137 549
rect 2091 477 2137 515
rect 2091 443 2097 477
rect 2131 443 2137 477
rect 2091 405 2137 443
rect 2091 371 2097 405
rect 2131 371 2137 405
rect 2091 355 2137 371
rect 2549 1629 2595 1645
rect 2549 1595 2555 1629
rect 2589 1595 2595 1629
rect 2549 1557 2595 1595
rect 2549 1523 2555 1557
rect 2589 1523 2595 1557
rect 2549 1485 2595 1523
rect 2549 1451 2555 1485
rect 2589 1451 2595 1485
rect 2549 1413 2595 1451
rect 2549 1379 2555 1413
rect 2589 1379 2595 1413
rect 2549 1341 2595 1379
rect 2549 1307 2555 1341
rect 2589 1307 2595 1341
rect 2549 1269 2595 1307
rect 2549 1235 2555 1269
rect 2589 1235 2595 1269
rect 2549 1197 2595 1235
rect 2549 1163 2555 1197
rect 2589 1163 2595 1197
rect 2549 1125 2595 1163
rect 2549 1091 2555 1125
rect 2589 1091 2595 1125
rect 2549 1053 2595 1091
rect 2549 1019 2555 1053
rect 2589 1019 2595 1053
rect 2549 981 2595 1019
rect 2549 947 2555 981
rect 2589 947 2595 981
rect 2549 909 2595 947
rect 2549 875 2555 909
rect 2589 875 2595 909
rect 2549 837 2595 875
rect 2549 803 2555 837
rect 2589 803 2595 837
rect 2549 765 2595 803
rect 2549 731 2555 765
rect 2589 731 2595 765
rect 2549 693 2595 731
rect 2549 659 2555 693
rect 2589 659 2595 693
rect 2549 621 2595 659
rect 2549 587 2555 621
rect 2589 587 2595 621
rect 2549 549 2595 587
rect 2549 515 2555 549
rect 2589 515 2595 549
rect 2549 477 2595 515
rect 2549 443 2555 477
rect 2589 443 2595 477
rect 2549 405 2595 443
rect 2549 371 2555 405
rect 2589 371 2595 405
rect 2549 355 2595 371
rect 3007 1629 3053 1645
rect 3007 1595 3013 1629
rect 3047 1595 3053 1629
rect 3007 1557 3053 1595
rect 3007 1523 3013 1557
rect 3047 1523 3053 1557
rect 3007 1485 3053 1523
rect 3007 1451 3013 1485
rect 3047 1451 3053 1485
rect 3007 1413 3053 1451
rect 3007 1379 3013 1413
rect 3047 1379 3053 1413
rect 3007 1341 3053 1379
rect 3007 1307 3013 1341
rect 3047 1307 3053 1341
rect 3007 1269 3053 1307
rect 3007 1235 3013 1269
rect 3047 1235 3053 1269
rect 3007 1197 3053 1235
rect 3007 1163 3013 1197
rect 3047 1163 3053 1197
rect 3007 1125 3053 1163
rect 3007 1091 3013 1125
rect 3047 1091 3053 1125
rect 3007 1053 3053 1091
rect 3007 1019 3013 1053
rect 3047 1019 3053 1053
rect 3007 981 3053 1019
rect 3007 947 3013 981
rect 3047 947 3053 981
rect 3007 909 3053 947
rect 3007 875 3013 909
rect 3047 875 3053 909
rect 3007 837 3053 875
rect 3007 803 3013 837
rect 3047 803 3053 837
rect 3007 765 3053 803
rect 3007 731 3013 765
rect 3047 731 3053 765
rect 3007 693 3053 731
rect 3007 659 3013 693
rect 3047 659 3053 693
rect 3007 621 3053 659
rect 3007 587 3013 621
rect 3047 587 3053 621
rect 3007 549 3053 587
rect 3007 515 3013 549
rect 3047 515 3053 549
rect 3007 477 3053 515
rect 3007 443 3013 477
rect 3047 443 3053 477
rect 3007 405 3053 443
rect 3007 371 3013 405
rect 3047 371 3053 405
rect 3007 355 3053 371
rect 3465 1629 3511 1645
rect 3465 1595 3471 1629
rect 3505 1595 3511 1629
rect 3465 1557 3511 1595
rect 3465 1523 3471 1557
rect 3505 1523 3511 1557
rect 3465 1485 3511 1523
rect 3465 1451 3471 1485
rect 3505 1451 3511 1485
rect 3465 1413 3511 1451
rect 3465 1379 3471 1413
rect 3505 1379 3511 1413
rect 3465 1341 3511 1379
rect 3465 1307 3471 1341
rect 3505 1307 3511 1341
rect 3465 1269 3511 1307
rect 3465 1235 3471 1269
rect 3505 1235 3511 1269
rect 3465 1197 3511 1235
rect 3465 1163 3471 1197
rect 3505 1163 3511 1197
rect 3465 1125 3511 1163
rect 3465 1091 3471 1125
rect 3505 1091 3511 1125
rect 3465 1053 3511 1091
rect 3465 1019 3471 1053
rect 3505 1019 3511 1053
rect 3465 981 3511 1019
rect 3465 947 3471 981
rect 3505 947 3511 981
rect 3465 909 3511 947
rect 3465 875 3471 909
rect 3505 875 3511 909
rect 3465 837 3511 875
rect 3465 803 3471 837
rect 3505 803 3511 837
rect 3465 765 3511 803
rect 3465 731 3471 765
rect 3505 731 3511 765
rect 3465 693 3511 731
rect 3465 659 3471 693
rect 3505 659 3511 693
rect 3465 621 3511 659
rect 3465 587 3471 621
rect 3505 587 3511 621
rect 3465 549 3511 587
rect 3465 515 3471 549
rect 3505 515 3511 549
rect 3465 477 3511 515
rect 3465 443 3471 477
rect 3505 443 3511 477
rect 3465 405 3511 443
rect 3465 371 3471 405
rect 3505 371 3511 405
rect 3465 355 3511 371
rect 3923 1629 3969 1645
rect 3923 1595 3929 1629
rect 3963 1595 3969 1629
rect 3923 1557 3969 1595
rect 3923 1523 3929 1557
rect 3963 1523 3969 1557
rect 3923 1485 3969 1523
rect 3923 1451 3929 1485
rect 3963 1451 3969 1485
rect 3923 1413 3969 1451
rect 3923 1379 3929 1413
rect 3963 1379 3969 1413
rect 3923 1341 3969 1379
rect 3923 1307 3929 1341
rect 3963 1307 3969 1341
rect 3923 1269 3969 1307
rect 3923 1235 3929 1269
rect 3963 1235 3969 1269
rect 3923 1197 3969 1235
rect 3923 1163 3929 1197
rect 3963 1163 3969 1197
rect 3923 1125 3969 1163
rect 3923 1091 3929 1125
rect 3963 1091 3969 1125
rect 3923 1053 3969 1091
rect 3923 1019 3929 1053
rect 3963 1019 3969 1053
rect 3923 981 3969 1019
rect 3923 947 3929 981
rect 3963 947 3969 981
rect 3923 909 3969 947
rect 3923 875 3929 909
rect 3963 875 3969 909
rect 3923 837 3969 875
rect 3923 803 3929 837
rect 3963 803 3969 837
rect 3923 765 3969 803
rect 3923 731 3929 765
rect 3963 731 3969 765
rect 3923 693 3969 731
rect 3923 659 3929 693
rect 3963 659 3969 693
rect 3923 621 3969 659
rect 3923 587 3929 621
rect 3963 587 3969 621
rect 3923 549 3969 587
rect 3923 515 3929 549
rect 3963 515 3969 549
rect 3923 477 3969 515
rect 3923 443 3929 477
rect 3963 443 3969 477
rect 3923 405 3969 443
rect 3923 371 3929 405
rect 3963 371 3969 405
rect 3923 355 3969 371
rect 4381 1629 4427 1645
rect 4381 1595 4387 1629
rect 4421 1595 4427 1629
rect 4381 1557 4427 1595
rect 4381 1523 4387 1557
rect 4421 1523 4427 1557
rect 4381 1485 4427 1523
rect 4381 1451 4387 1485
rect 4421 1451 4427 1485
rect 4381 1413 4427 1451
rect 4381 1379 4387 1413
rect 4421 1379 4427 1413
rect 4381 1341 4427 1379
rect 4381 1307 4387 1341
rect 4421 1307 4427 1341
rect 4381 1269 4427 1307
rect 4381 1235 4387 1269
rect 4421 1235 4427 1269
rect 4381 1197 4427 1235
rect 4381 1163 4387 1197
rect 4421 1163 4427 1197
rect 4381 1125 4427 1163
rect 4381 1091 4387 1125
rect 4421 1091 4427 1125
rect 4381 1053 4427 1091
rect 4381 1019 4387 1053
rect 4421 1019 4427 1053
rect 4381 981 4427 1019
rect 4381 947 4387 981
rect 4421 947 4427 981
rect 4381 909 4427 947
rect 4381 875 4387 909
rect 4421 875 4427 909
rect 4381 837 4427 875
rect 4381 803 4387 837
rect 4421 803 4427 837
rect 4381 765 4427 803
rect 4381 731 4387 765
rect 4421 731 4427 765
rect 4381 693 4427 731
rect 4381 659 4387 693
rect 4421 659 4427 693
rect 4381 621 4427 659
rect 4381 587 4387 621
rect 4421 587 4427 621
rect 4381 549 4427 587
rect 4381 515 4387 549
rect 4421 515 4427 549
rect 4381 477 4427 515
rect 4381 443 4387 477
rect 4421 443 4427 477
rect 4381 405 4427 443
rect 4381 371 4387 405
rect 4421 371 4427 405
rect 4381 355 4427 371
rect 4839 1629 4885 1645
rect 4839 1595 4845 1629
rect 4879 1595 4885 1629
rect 4839 1557 4885 1595
rect 4839 1523 4845 1557
rect 4879 1523 4885 1557
rect 4839 1485 4885 1523
rect 4839 1451 4845 1485
rect 4879 1451 4885 1485
rect 4839 1413 4885 1451
rect 4839 1379 4845 1413
rect 4879 1379 4885 1413
rect 4839 1341 4885 1379
rect 4839 1307 4845 1341
rect 4879 1307 4885 1341
rect 4839 1269 4885 1307
rect 4839 1235 4845 1269
rect 4879 1235 4885 1269
rect 4839 1197 4885 1235
rect 4839 1163 4845 1197
rect 4879 1163 4885 1197
rect 4839 1125 4885 1163
rect 4839 1091 4845 1125
rect 4879 1091 4885 1125
rect 4839 1053 4885 1091
rect 4839 1019 4845 1053
rect 4879 1019 4885 1053
rect 4839 981 4885 1019
rect 4839 947 4845 981
rect 4879 947 4885 981
rect 4839 909 4885 947
rect 4839 875 4845 909
rect 4879 875 4885 909
rect 4839 837 4885 875
rect 4839 803 4845 837
rect 4879 803 4885 837
rect 4839 765 4885 803
rect 4839 731 4845 765
rect 4879 731 4885 765
rect 4839 693 4885 731
rect 4839 659 4845 693
rect 4879 659 4885 693
rect 4839 621 4885 659
rect 4839 587 4845 621
rect 4879 587 4885 621
rect 4839 549 4885 587
rect 4839 515 4845 549
rect 4879 515 4885 549
rect 4839 477 4885 515
rect 4839 443 4845 477
rect 4879 443 4885 477
rect 4839 405 4885 443
rect 4839 371 4845 405
rect 4879 371 4885 405
rect 4839 355 4885 371
rect 5297 1629 5343 1645
rect 5297 1595 5303 1629
rect 5337 1595 5343 1629
rect 5297 1557 5343 1595
rect 5297 1523 5303 1557
rect 5337 1523 5343 1557
rect 5297 1485 5343 1523
rect 5297 1451 5303 1485
rect 5337 1451 5343 1485
rect 5297 1413 5343 1451
rect 5297 1379 5303 1413
rect 5337 1379 5343 1413
rect 5297 1341 5343 1379
rect 5297 1307 5303 1341
rect 5337 1307 5343 1341
rect 5297 1269 5343 1307
rect 5297 1235 5303 1269
rect 5337 1235 5343 1269
rect 5297 1197 5343 1235
rect 5297 1163 5303 1197
rect 5337 1163 5343 1197
rect 5297 1125 5343 1163
rect 5297 1091 5303 1125
rect 5337 1091 5343 1125
rect 5297 1053 5343 1091
rect 5297 1019 5303 1053
rect 5337 1019 5343 1053
rect 5297 981 5343 1019
rect 5297 947 5303 981
rect 5337 947 5343 981
rect 5297 909 5343 947
rect 5297 875 5303 909
rect 5337 875 5343 909
rect 5297 837 5343 875
rect 5297 803 5303 837
rect 5337 803 5343 837
rect 5297 765 5343 803
rect 5297 731 5303 765
rect 5337 731 5343 765
rect 5297 693 5343 731
rect 5297 659 5303 693
rect 5337 659 5343 693
rect 5297 621 5343 659
rect 5297 587 5303 621
rect 5337 587 5343 621
rect 5297 549 5343 587
rect 5297 515 5303 549
rect 5337 515 5343 549
rect 5297 477 5343 515
rect 5297 443 5303 477
rect 5337 443 5343 477
rect 5297 405 5343 443
rect 5297 371 5303 405
rect 5337 371 5343 405
rect 5297 355 5343 371
rect 5755 1629 5801 1645
rect 5755 1595 5761 1629
rect 5795 1595 5801 1629
rect 5755 1557 5801 1595
rect 5755 1523 5761 1557
rect 5795 1523 5801 1557
rect 5755 1485 5801 1523
rect 5755 1451 5761 1485
rect 5795 1451 5801 1485
rect 5755 1413 5801 1451
rect 5755 1379 5761 1413
rect 5795 1379 5801 1413
rect 5755 1341 5801 1379
rect 5755 1307 5761 1341
rect 5795 1307 5801 1341
rect 5755 1269 5801 1307
rect 5755 1235 5761 1269
rect 5795 1235 5801 1269
rect 5755 1197 5801 1235
rect 5755 1163 5761 1197
rect 5795 1163 5801 1197
rect 5755 1125 5801 1163
rect 5755 1091 5761 1125
rect 5795 1091 5801 1125
rect 5755 1053 5801 1091
rect 5755 1019 5761 1053
rect 5795 1019 5801 1053
rect 5755 981 5801 1019
rect 5755 947 5761 981
rect 5795 947 5801 981
rect 5755 909 5801 947
rect 5755 875 5761 909
rect 5795 875 5801 909
rect 5755 837 5801 875
rect 5755 803 5761 837
rect 5795 803 5801 837
rect 5755 765 5801 803
rect 5755 731 5761 765
rect 5795 731 5801 765
rect 5755 693 5801 731
rect 5755 659 5761 693
rect 5795 659 5801 693
rect 5755 621 5801 659
rect 5755 587 5761 621
rect 5795 587 5801 621
rect 5755 549 5801 587
rect 5755 515 5761 549
rect 5795 515 5801 549
rect 5755 477 5801 515
rect 5755 443 5761 477
rect 5795 443 5801 477
rect 5755 405 5801 443
rect 5755 371 5761 405
rect 5795 371 5801 405
rect 5755 355 5801 371
rect 6213 1629 6259 1645
rect 6213 1595 6219 1629
rect 6253 1595 6259 1629
rect 6213 1557 6259 1595
rect 6213 1523 6219 1557
rect 6253 1523 6259 1557
rect 6213 1485 6259 1523
rect 6213 1451 6219 1485
rect 6253 1451 6259 1485
rect 6213 1413 6259 1451
rect 6213 1379 6219 1413
rect 6253 1379 6259 1413
rect 6213 1341 6259 1379
rect 6213 1307 6219 1341
rect 6253 1307 6259 1341
rect 6213 1269 6259 1307
rect 6213 1235 6219 1269
rect 6253 1235 6259 1269
rect 6213 1197 6259 1235
rect 6213 1163 6219 1197
rect 6253 1163 6259 1197
rect 6213 1125 6259 1163
rect 6213 1091 6219 1125
rect 6253 1091 6259 1125
rect 6213 1053 6259 1091
rect 6213 1019 6219 1053
rect 6253 1019 6259 1053
rect 6213 981 6259 1019
rect 6213 947 6219 981
rect 6253 947 6259 981
rect 6213 909 6259 947
rect 6213 875 6219 909
rect 6253 875 6259 909
rect 6213 837 6259 875
rect 6213 803 6219 837
rect 6253 803 6259 837
rect 6213 765 6259 803
rect 6213 731 6219 765
rect 6253 731 6259 765
rect 6213 693 6259 731
rect 6213 659 6219 693
rect 6253 659 6259 693
rect 6213 621 6259 659
rect 6213 587 6219 621
rect 6253 587 6259 621
rect 6213 549 6259 587
rect 6213 515 6219 549
rect 6253 515 6259 549
rect 6213 477 6259 515
rect 6213 443 6219 477
rect 6253 443 6259 477
rect 6213 405 6259 443
rect 6213 371 6219 405
rect 6253 371 6259 405
rect 6213 355 6259 371
rect 6671 1629 6717 1645
rect 6671 1595 6677 1629
rect 6711 1595 6717 1629
rect 6671 1557 6717 1595
rect 6671 1523 6677 1557
rect 6711 1523 6717 1557
rect 6671 1485 6717 1523
rect 6671 1451 6677 1485
rect 6711 1451 6717 1485
rect 6671 1413 6717 1451
rect 6671 1379 6677 1413
rect 6711 1379 6717 1413
rect 6671 1341 6717 1379
rect 6671 1307 6677 1341
rect 6711 1307 6717 1341
rect 6671 1269 6717 1307
rect 6671 1235 6677 1269
rect 6711 1235 6717 1269
rect 6671 1197 6717 1235
rect 6671 1163 6677 1197
rect 6711 1163 6717 1197
rect 6671 1125 6717 1163
rect 6671 1091 6677 1125
rect 6711 1091 6717 1125
rect 6671 1053 6717 1091
rect 6671 1019 6677 1053
rect 6711 1019 6717 1053
rect 6671 981 6717 1019
rect 6671 947 6677 981
rect 6711 947 6717 981
rect 6671 909 6717 947
rect 6671 875 6677 909
rect 6711 875 6717 909
rect 6671 837 6717 875
rect 6671 803 6677 837
rect 6711 803 6717 837
rect 6671 765 6717 803
rect 6671 731 6677 765
rect 6711 731 6717 765
rect 6671 693 6717 731
rect 6671 659 6677 693
rect 6711 659 6717 693
rect 6671 621 6717 659
rect 6671 587 6677 621
rect 6711 587 6717 621
rect 6671 549 6717 587
rect 6671 515 6677 549
rect 6711 515 6717 549
rect 6671 477 6717 515
rect 6671 443 6677 477
rect 6711 443 6717 477
rect 6671 405 6717 443
rect 6671 371 6677 405
rect 6711 371 6717 405
rect 6671 355 6717 371
rect 7129 1629 7175 1645
rect 7129 1595 7135 1629
rect 7169 1595 7175 1629
rect 7129 1557 7175 1595
rect 7129 1523 7135 1557
rect 7169 1523 7175 1557
rect 7129 1485 7175 1523
rect 7129 1451 7135 1485
rect 7169 1451 7175 1485
rect 7129 1413 7175 1451
rect 7129 1379 7135 1413
rect 7169 1379 7175 1413
rect 7129 1341 7175 1379
rect 7129 1307 7135 1341
rect 7169 1307 7175 1341
rect 7129 1269 7175 1307
rect 7129 1235 7135 1269
rect 7169 1235 7175 1269
rect 7129 1197 7175 1235
rect 7129 1163 7135 1197
rect 7169 1163 7175 1197
rect 7129 1125 7175 1163
rect 7129 1091 7135 1125
rect 7169 1091 7175 1125
rect 7129 1053 7175 1091
rect 7129 1019 7135 1053
rect 7169 1019 7175 1053
rect 7129 981 7175 1019
rect 7129 947 7135 981
rect 7169 947 7175 981
rect 7129 909 7175 947
rect 7129 875 7135 909
rect 7169 875 7175 909
rect 7129 837 7175 875
rect 7129 803 7135 837
rect 7169 803 7175 837
rect 7129 765 7175 803
rect 7129 731 7135 765
rect 7169 731 7175 765
rect 7129 693 7175 731
rect 7129 659 7135 693
rect 7169 659 7175 693
rect 7129 621 7175 659
rect 7129 587 7135 621
rect 7169 587 7175 621
rect 7129 549 7175 587
rect 7129 515 7135 549
rect 7169 515 7175 549
rect 7129 477 7175 515
rect 7129 443 7135 477
rect 7169 443 7175 477
rect 7129 405 7175 443
rect 7129 371 7135 405
rect 7169 371 7175 405
rect 7129 355 7175 371
rect 7587 1629 7633 1645
rect 7587 1595 7593 1629
rect 7627 1595 7633 1629
rect 7587 1557 7633 1595
rect 7587 1523 7593 1557
rect 7627 1523 7633 1557
rect 7587 1485 7633 1523
rect 7587 1451 7593 1485
rect 7627 1451 7633 1485
rect 7587 1413 7633 1451
rect 7587 1379 7593 1413
rect 7627 1379 7633 1413
rect 7587 1341 7633 1379
rect 7587 1307 7593 1341
rect 7627 1307 7633 1341
rect 7587 1269 7633 1307
rect 7587 1235 7593 1269
rect 7627 1235 7633 1269
rect 7587 1197 7633 1235
rect 7587 1163 7593 1197
rect 7627 1163 7633 1197
rect 7587 1125 7633 1163
rect 7587 1091 7593 1125
rect 7627 1091 7633 1125
rect 7587 1053 7633 1091
rect 7587 1019 7593 1053
rect 7627 1019 7633 1053
rect 7587 981 7633 1019
rect 7587 947 7593 981
rect 7627 947 7633 981
rect 7587 909 7633 947
rect 7587 875 7593 909
rect 7627 875 7633 909
rect 7587 837 7633 875
rect 7587 803 7593 837
rect 7627 803 7633 837
rect 7587 765 7633 803
rect 7587 731 7593 765
rect 7627 731 7633 765
rect 7587 693 7633 731
rect 7587 659 7593 693
rect 7627 659 7633 693
rect 7587 621 7633 659
rect 7587 587 7593 621
rect 7627 587 7633 621
rect 7587 549 7633 587
rect 7587 515 7593 549
rect 7627 515 7633 549
rect 7587 477 7633 515
rect 7587 443 7593 477
rect 7627 443 7633 477
rect 7587 405 7633 443
rect 7587 371 7593 405
rect 7627 371 7633 405
rect 7587 355 7633 371
rect 8045 1629 8091 1645
rect 8045 1595 8051 1629
rect 8085 1595 8091 1629
rect 8045 1557 8091 1595
rect 8045 1523 8051 1557
rect 8085 1523 8091 1557
rect 8045 1485 8091 1523
rect 8045 1451 8051 1485
rect 8085 1451 8091 1485
rect 8045 1413 8091 1451
rect 8045 1379 8051 1413
rect 8085 1379 8091 1413
rect 8045 1341 8091 1379
rect 8045 1307 8051 1341
rect 8085 1307 8091 1341
rect 8045 1269 8091 1307
rect 8045 1235 8051 1269
rect 8085 1235 8091 1269
rect 8045 1197 8091 1235
rect 8045 1163 8051 1197
rect 8085 1163 8091 1197
rect 8045 1125 8091 1163
rect 8045 1091 8051 1125
rect 8085 1091 8091 1125
rect 8045 1053 8091 1091
rect 8045 1019 8051 1053
rect 8085 1019 8091 1053
rect 8045 981 8091 1019
rect 8045 947 8051 981
rect 8085 947 8091 981
rect 8045 909 8091 947
rect 8045 875 8051 909
rect 8085 875 8091 909
rect 8045 837 8091 875
rect 8045 803 8051 837
rect 8085 803 8091 837
rect 8045 765 8091 803
rect 8045 731 8051 765
rect 8085 731 8091 765
rect 8045 693 8091 731
rect 8045 659 8051 693
rect 8085 659 8091 693
rect 8045 621 8091 659
rect 8045 587 8051 621
rect 8085 587 8091 621
rect 8045 549 8091 587
rect 8045 515 8051 549
rect 8085 515 8091 549
rect 8045 477 8091 515
rect 8045 443 8051 477
rect 8085 443 8091 477
rect 8045 405 8091 443
rect 8045 371 8051 405
rect 8085 371 8091 405
rect 8045 355 8091 371
rect 8503 1629 8549 1645
rect 8503 1595 8509 1629
rect 8543 1595 8549 1629
rect 8503 1557 8549 1595
rect 8503 1523 8509 1557
rect 8543 1523 8549 1557
rect 8503 1485 8549 1523
rect 8503 1451 8509 1485
rect 8543 1451 8549 1485
rect 8503 1413 8549 1451
rect 8503 1379 8509 1413
rect 8543 1379 8549 1413
rect 8503 1341 8549 1379
rect 8503 1307 8509 1341
rect 8543 1307 8549 1341
rect 8503 1269 8549 1307
rect 8503 1235 8509 1269
rect 8543 1235 8549 1269
rect 8503 1197 8549 1235
rect 8503 1163 8509 1197
rect 8543 1163 8549 1197
rect 8503 1125 8549 1163
rect 8503 1091 8509 1125
rect 8543 1091 8549 1125
rect 8503 1053 8549 1091
rect 8503 1019 8509 1053
rect 8543 1019 8549 1053
rect 8503 981 8549 1019
rect 8503 947 8509 981
rect 8543 947 8549 981
rect 8503 909 8549 947
rect 8503 875 8509 909
rect 8543 875 8549 909
rect 8503 837 8549 875
rect 8503 803 8509 837
rect 8543 803 8549 837
rect 8503 765 8549 803
rect 8503 731 8509 765
rect 8543 731 8549 765
rect 8503 693 8549 731
rect 8503 659 8509 693
rect 8543 659 8549 693
rect 8503 621 8549 659
rect 8503 587 8509 621
rect 8543 587 8549 621
rect 8503 549 8549 587
rect 8503 515 8509 549
rect 8543 515 8549 549
rect 8503 477 8549 515
rect 8503 443 8509 477
rect 8543 443 8549 477
rect 8503 405 8549 443
rect 8503 371 8509 405
rect 8543 371 8549 405
rect 8503 355 8549 371
rect 8961 1629 9007 1645
rect 8961 1595 8967 1629
rect 9001 1595 9007 1629
rect 8961 1557 9007 1595
rect 8961 1523 8967 1557
rect 9001 1523 9007 1557
rect 8961 1485 9007 1523
rect 8961 1451 8967 1485
rect 9001 1451 9007 1485
rect 8961 1413 9007 1451
rect 8961 1379 8967 1413
rect 9001 1379 9007 1413
rect 8961 1341 9007 1379
rect 8961 1307 8967 1341
rect 9001 1307 9007 1341
rect 8961 1269 9007 1307
rect 8961 1235 8967 1269
rect 9001 1235 9007 1269
rect 8961 1197 9007 1235
rect 8961 1163 8967 1197
rect 9001 1163 9007 1197
rect 8961 1125 9007 1163
rect 8961 1091 8967 1125
rect 9001 1091 9007 1125
rect 8961 1053 9007 1091
rect 8961 1019 8967 1053
rect 9001 1019 9007 1053
rect 8961 981 9007 1019
rect 8961 947 8967 981
rect 9001 947 9007 981
rect 8961 909 9007 947
rect 8961 875 8967 909
rect 9001 875 9007 909
rect 8961 837 9007 875
rect 8961 803 8967 837
rect 9001 803 9007 837
rect 8961 765 9007 803
rect 8961 731 8967 765
rect 9001 731 9007 765
rect 8961 693 9007 731
rect 8961 659 8967 693
rect 9001 659 9007 693
rect 8961 621 9007 659
rect 8961 587 8967 621
rect 9001 587 9007 621
rect 8961 549 9007 587
rect 8961 515 8967 549
rect 9001 515 9007 549
rect 8961 477 9007 515
rect 8961 443 8967 477
rect 9001 443 9007 477
rect 8961 405 9007 443
rect 8961 371 8967 405
rect 9001 371 9007 405
rect 8961 355 9007 371
rect 9419 1629 9465 1645
rect 9419 1595 9425 1629
rect 9459 1595 9465 1629
rect 9419 1557 9465 1595
rect 9419 1523 9425 1557
rect 9459 1523 9465 1557
rect 9419 1485 9465 1523
rect 9419 1451 9425 1485
rect 9459 1451 9465 1485
rect 9419 1413 9465 1451
rect 9419 1379 9425 1413
rect 9459 1379 9465 1413
rect 9419 1341 9465 1379
rect 9419 1307 9425 1341
rect 9459 1307 9465 1341
rect 9419 1269 9465 1307
rect 9419 1235 9425 1269
rect 9459 1235 9465 1269
rect 9419 1197 9465 1235
rect 9419 1163 9425 1197
rect 9459 1163 9465 1197
rect 9419 1125 9465 1163
rect 9419 1091 9425 1125
rect 9459 1091 9465 1125
rect 9419 1053 9465 1091
rect 9419 1019 9425 1053
rect 9459 1019 9465 1053
rect 9419 981 9465 1019
rect 9419 947 9425 981
rect 9459 947 9465 981
rect 9419 909 9465 947
rect 9419 875 9425 909
rect 9459 875 9465 909
rect 9419 837 9465 875
rect 9419 803 9425 837
rect 9459 803 9465 837
rect 9419 765 9465 803
rect 9419 731 9425 765
rect 9459 731 9465 765
rect 9419 693 9465 731
rect 9419 659 9425 693
rect 9459 659 9465 693
rect 9419 621 9465 659
rect 9419 587 9425 621
rect 9459 587 9465 621
rect 9419 549 9465 587
rect 9419 515 9425 549
rect 9459 515 9465 549
rect 9419 477 9465 515
rect 9419 443 9425 477
rect 9459 443 9465 477
rect 9419 405 9465 443
rect 9419 371 9425 405
rect 9459 371 9465 405
rect 9419 355 9465 371
rect 9877 1629 9923 1645
rect 9877 1595 9883 1629
rect 9917 1595 9923 1629
rect 9877 1557 9923 1595
rect 9877 1523 9883 1557
rect 9917 1523 9923 1557
rect 9877 1485 9923 1523
rect 9877 1451 9883 1485
rect 9917 1451 9923 1485
rect 9877 1413 9923 1451
rect 9877 1379 9883 1413
rect 9917 1379 9923 1413
rect 9877 1341 9923 1379
rect 9877 1307 9883 1341
rect 9917 1307 9923 1341
rect 9877 1269 9923 1307
rect 9877 1235 9883 1269
rect 9917 1235 9923 1269
rect 9877 1197 9923 1235
rect 9877 1163 9883 1197
rect 9917 1163 9923 1197
rect 9877 1125 9923 1163
rect 9877 1091 9883 1125
rect 9917 1091 9923 1125
rect 9877 1053 9923 1091
rect 9877 1019 9883 1053
rect 9917 1019 9923 1053
rect 9877 981 9923 1019
rect 9877 947 9883 981
rect 9917 947 9923 981
rect 9877 909 9923 947
rect 9877 875 9883 909
rect 9917 875 9923 909
rect 9877 837 9923 875
rect 9877 803 9883 837
rect 9917 803 9923 837
rect 9877 765 9923 803
rect 9877 731 9883 765
rect 9917 731 9923 765
rect 9877 693 9923 731
rect 9877 659 9883 693
rect 9917 659 9923 693
rect 9877 621 9923 659
rect 9877 587 9883 621
rect 9917 587 9923 621
rect 9877 549 9923 587
rect 9877 515 9883 549
rect 9917 515 9923 549
rect 9877 477 9923 515
rect 9877 443 9883 477
rect 9917 443 9923 477
rect 9877 405 9923 443
rect 9877 371 9883 405
rect 9917 371 9923 405
rect 9877 355 9923 371
rect 10335 1629 10381 1645
rect 10335 1595 10341 1629
rect 10375 1595 10381 1629
rect 10335 1557 10381 1595
rect 10335 1523 10341 1557
rect 10375 1523 10381 1557
rect 10335 1485 10381 1523
rect 10335 1451 10341 1485
rect 10375 1451 10381 1485
rect 10335 1413 10381 1451
rect 10335 1379 10341 1413
rect 10375 1379 10381 1413
rect 10335 1341 10381 1379
rect 10335 1307 10341 1341
rect 10375 1307 10381 1341
rect 10335 1269 10381 1307
rect 10335 1235 10341 1269
rect 10375 1235 10381 1269
rect 10335 1197 10381 1235
rect 10335 1163 10341 1197
rect 10375 1163 10381 1197
rect 10335 1125 10381 1163
rect 10335 1091 10341 1125
rect 10375 1091 10381 1125
rect 10335 1053 10381 1091
rect 10335 1019 10341 1053
rect 10375 1019 10381 1053
rect 10335 981 10381 1019
rect 10335 947 10341 981
rect 10375 947 10381 981
rect 10335 909 10381 947
rect 10335 875 10341 909
rect 10375 875 10381 909
rect 10335 837 10381 875
rect 10335 803 10341 837
rect 10375 803 10381 837
rect 10335 765 10381 803
rect 10335 731 10341 765
rect 10375 731 10381 765
rect 10335 693 10381 731
rect 10335 659 10341 693
rect 10375 659 10381 693
rect 10335 621 10381 659
rect 10335 587 10341 621
rect 10375 587 10381 621
rect 10335 549 10381 587
rect 10335 515 10341 549
rect 10375 515 10381 549
rect 10335 477 10381 515
rect 10335 443 10341 477
rect 10375 443 10381 477
rect 10335 405 10381 443
rect 10335 371 10341 405
rect 10375 371 10381 405
rect 10335 355 10381 371
rect 10793 1629 10839 1645
rect 10793 1595 10799 1629
rect 10833 1595 10839 1629
rect 10793 1557 10839 1595
rect 10793 1523 10799 1557
rect 10833 1523 10839 1557
rect 10793 1485 10839 1523
rect 10793 1451 10799 1485
rect 10833 1451 10839 1485
rect 10793 1413 10839 1451
rect 10793 1379 10799 1413
rect 10833 1379 10839 1413
rect 10793 1341 10839 1379
rect 10793 1307 10799 1341
rect 10833 1307 10839 1341
rect 10793 1269 10839 1307
rect 10793 1235 10799 1269
rect 10833 1235 10839 1269
rect 10793 1197 10839 1235
rect 10793 1163 10799 1197
rect 10833 1163 10839 1197
rect 10793 1125 10839 1163
rect 10793 1091 10799 1125
rect 10833 1091 10839 1125
rect 10793 1053 10839 1091
rect 10793 1019 10799 1053
rect 10833 1019 10839 1053
rect 10793 981 10839 1019
rect 10793 947 10799 981
rect 10833 947 10839 981
rect 10793 909 10839 947
rect 10793 875 10799 909
rect 10833 875 10839 909
rect 10793 837 10839 875
rect 10793 803 10799 837
rect 10833 803 10839 837
rect 10793 765 10839 803
rect 10793 731 10799 765
rect 10833 731 10839 765
rect 10793 693 10839 731
rect 10793 659 10799 693
rect 10833 659 10839 693
rect 10793 621 10839 659
rect 10793 587 10799 621
rect 10833 587 10839 621
rect 10793 549 10839 587
rect 10793 515 10799 549
rect 10833 515 10839 549
rect 10793 477 10839 515
rect 10793 443 10799 477
rect 10833 443 10839 477
rect 10793 405 10839 443
rect 10793 371 10799 405
rect 10833 371 10839 405
rect 10793 355 10839 371
rect 11251 1629 11297 1645
rect 11251 1595 11257 1629
rect 11291 1595 11297 1629
rect 11251 1557 11297 1595
rect 11251 1523 11257 1557
rect 11291 1523 11297 1557
rect 11251 1485 11297 1523
rect 11251 1451 11257 1485
rect 11291 1451 11297 1485
rect 11251 1413 11297 1451
rect 11251 1379 11257 1413
rect 11291 1379 11297 1413
rect 11251 1341 11297 1379
rect 11251 1307 11257 1341
rect 11291 1307 11297 1341
rect 11251 1269 11297 1307
rect 11251 1235 11257 1269
rect 11291 1235 11297 1269
rect 11251 1197 11297 1235
rect 11251 1163 11257 1197
rect 11291 1163 11297 1197
rect 11251 1125 11297 1163
rect 11251 1091 11257 1125
rect 11291 1091 11297 1125
rect 11251 1053 11297 1091
rect 11251 1019 11257 1053
rect 11291 1019 11297 1053
rect 11251 981 11297 1019
rect 11251 947 11257 981
rect 11291 947 11297 981
rect 11251 909 11297 947
rect 11251 875 11257 909
rect 11291 875 11297 909
rect 11251 837 11297 875
rect 11251 803 11257 837
rect 11291 803 11297 837
rect 11251 765 11297 803
rect 11251 731 11257 765
rect 11291 731 11297 765
rect 11251 693 11297 731
rect 11251 659 11257 693
rect 11291 659 11297 693
rect 11251 621 11297 659
rect 11251 587 11257 621
rect 11291 587 11297 621
rect 11251 549 11297 587
rect 11251 515 11257 549
rect 11291 515 11297 549
rect 11251 477 11297 515
rect 11251 443 11257 477
rect 11291 443 11297 477
rect 11251 405 11297 443
rect 11251 371 11257 405
rect 11291 371 11297 405
rect 11251 355 11297 371
rect 11709 1629 11755 1645
rect 11709 1595 11715 1629
rect 11749 1595 11755 1629
rect 11709 1557 11755 1595
rect 11709 1523 11715 1557
rect 11749 1523 11755 1557
rect 11709 1485 11755 1523
rect 11709 1451 11715 1485
rect 11749 1451 11755 1485
rect 11709 1413 11755 1451
rect 11709 1379 11715 1413
rect 11749 1379 11755 1413
rect 11709 1341 11755 1379
rect 11709 1307 11715 1341
rect 11749 1307 11755 1341
rect 11709 1269 11755 1307
rect 11709 1235 11715 1269
rect 11749 1235 11755 1269
rect 11709 1197 11755 1235
rect 11709 1163 11715 1197
rect 11749 1163 11755 1197
rect 11709 1125 11755 1163
rect 11709 1091 11715 1125
rect 11749 1091 11755 1125
rect 11709 1053 11755 1091
rect 11709 1019 11715 1053
rect 11749 1019 11755 1053
rect 11709 981 11755 1019
rect 11709 947 11715 981
rect 11749 947 11755 981
rect 11709 909 11755 947
rect 11709 875 11715 909
rect 11749 875 11755 909
rect 11709 837 11755 875
rect 11709 803 11715 837
rect 11749 803 11755 837
rect 11709 765 11755 803
rect 11709 731 11715 765
rect 11749 731 11755 765
rect 11709 693 11755 731
rect 11709 659 11715 693
rect 11749 659 11755 693
rect 11709 621 11755 659
rect 11709 587 11715 621
rect 11749 587 11755 621
rect 11709 549 11755 587
rect 11709 515 11715 549
rect 11749 515 11755 549
rect 11709 477 11755 515
rect 11709 443 11715 477
rect 11749 443 11755 477
rect 11709 405 11755 443
rect 11709 371 11715 405
rect 11749 371 11755 405
rect 11709 355 11755 371
rect 12167 1629 12213 1645
rect 12167 1595 12173 1629
rect 12207 1595 12213 1629
rect 12167 1557 12213 1595
rect 12167 1523 12173 1557
rect 12207 1523 12213 1557
rect 12167 1485 12213 1523
rect 12167 1451 12173 1485
rect 12207 1451 12213 1485
rect 12167 1413 12213 1451
rect 12167 1379 12173 1413
rect 12207 1379 12213 1413
rect 12167 1341 12213 1379
rect 12167 1307 12173 1341
rect 12207 1307 12213 1341
rect 12167 1269 12213 1307
rect 12167 1235 12173 1269
rect 12207 1235 12213 1269
rect 12167 1197 12213 1235
rect 12167 1163 12173 1197
rect 12207 1163 12213 1197
rect 12167 1125 12213 1163
rect 12167 1091 12173 1125
rect 12207 1091 12213 1125
rect 12167 1053 12213 1091
rect 12167 1019 12173 1053
rect 12207 1019 12213 1053
rect 12167 981 12213 1019
rect 12167 947 12173 981
rect 12207 947 12213 981
rect 12167 909 12213 947
rect 12167 875 12173 909
rect 12207 875 12213 909
rect 12167 837 12213 875
rect 12167 803 12173 837
rect 12207 803 12213 837
rect 12167 765 12213 803
rect 12167 731 12173 765
rect 12207 731 12213 765
rect 12167 693 12213 731
rect 12167 659 12173 693
rect 12207 659 12213 693
rect 12167 621 12213 659
rect 12167 587 12173 621
rect 12207 587 12213 621
rect 12167 549 12213 587
rect 12167 515 12173 549
rect 12207 515 12213 549
rect 12167 477 12213 515
rect 12167 443 12173 477
rect 12207 443 12213 477
rect 12167 405 12213 443
rect 12167 371 12173 405
rect 12207 371 12213 405
rect 12167 355 12213 371
rect 12625 1629 12671 1645
rect 12625 1595 12631 1629
rect 12665 1595 12671 1629
rect 12625 1557 12671 1595
rect 12625 1523 12631 1557
rect 12665 1523 12671 1557
rect 12625 1485 12671 1523
rect 12625 1451 12631 1485
rect 12665 1451 12671 1485
rect 12625 1413 12671 1451
rect 12625 1379 12631 1413
rect 12665 1379 12671 1413
rect 12625 1341 12671 1379
rect 12625 1307 12631 1341
rect 12665 1307 12671 1341
rect 12625 1269 12671 1307
rect 12625 1235 12631 1269
rect 12665 1235 12671 1269
rect 12625 1197 12671 1235
rect 12625 1163 12631 1197
rect 12665 1163 12671 1197
rect 12625 1125 12671 1163
rect 12625 1091 12631 1125
rect 12665 1091 12671 1125
rect 12625 1053 12671 1091
rect 12625 1019 12631 1053
rect 12665 1019 12671 1053
rect 12625 981 12671 1019
rect 12625 947 12631 981
rect 12665 947 12671 981
rect 12625 909 12671 947
rect 12625 875 12631 909
rect 12665 875 12671 909
rect 12625 837 12671 875
rect 12625 803 12631 837
rect 12665 803 12671 837
rect 12625 765 12671 803
rect 12625 731 12631 765
rect 12665 731 12671 765
rect 12625 693 12671 731
rect 12625 659 12631 693
rect 12665 659 12671 693
rect 12625 621 12671 659
rect 12625 587 12631 621
rect 12665 587 12671 621
rect 12625 549 12671 587
rect 12625 515 12631 549
rect 12665 515 12671 549
rect 12625 477 12671 515
rect 12625 443 12631 477
rect 12665 443 12671 477
rect 12625 405 12671 443
rect 12625 371 12631 405
rect 12665 371 12671 405
rect 12625 355 12671 371
rect 13083 1629 13129 1645
rect 13083 1595 13089 1629
rect 13123 1595 13129 1629
rect 13083 1557 13129 1595
rect 13083 1523 13089 1557
rect 13123 1523 13129 1557
rect 13083 1485 13129 1523
rect 13083 1451 13089 1485
rect 13123 1451 13129 1485
rect 13083 1413 13129 1451
rect 13083 1379 13089 1413
rect 13123 1379 13129 1413
rect 13083 1341 13129 1379
rect 13083 1307 13089 1341
rect 13123 1307 13129 1341
rect 13083 1269 13129 1307
rect 13083 1235 13089 1269
rect 13123 1235 13129 1269
rect 13083 1197 13129 1235
rect 13083 1163 13089 1197
rect 13123 1163 13129 1197
rect 13083 1125 13129 1163
rect 13083 1091 13089 1125
rect 13123 1091 13129 1125
rect 13083 1053 13129 1091
rect 13083 1019 13089 1053
rect 13123 1019 13129 1053
rect 13083 981 13129 1019
rect 13083 947 13089 981
rect 13123 947 13129 981
rect 13083 909 13129 947
rect 13083 875 13089 909
rect 13123 875 13129 909
rect 13083 837 13129 875
rect 13083 803 13089 837
rect 13123 803 13129 837
rect 13083 765 13129 803
rect 13083 731 13089 765
rect 13123 731 13129 765
rect 13083 693 13129 731
rect 13083 659 13089 693
rect 13123 659 13129 693
rect 13083 621 13129 659
rect 13083 587 13089 621
rect 13123 587 13129 621
rect 13083 549 13129 587
rect 13083 515 13089 549
rect 13123 515 13129 549
rect 13083 477 13129 515
rect 13083 443 13089 477
rect 13123 443 13129 477
rect 13083 405 13129 443
rect 13083 371 13089 405
rect 13123 371 13129 405
rect 13083 355 13129 371
rect 13541 1629 13587 1645
rect 13541 1595 13547 1629
rect 13581 1595 13587 1629
rect 13541 1557 13587 1595
rect 13541 1523 13547 1557
rect 13581 1523 13587 1557
rect 13541 1485 13587 1523
rect 13541 1451 13547 1485
rect 13581 1451 13587 1485
rect 13541 1413 13587 1451
rect 13541 1379 13547 1413
rect 13581 1379 13587 1413
rect 13541 1341 13587 1379
rect 13541 1307 13547 1341
rect 13581 1307 13587 1341
rect 13541 1269 13587 1307
rect 13541 1235 13547 1269
rect 13581 1235 13587 1269
rect 13541 1197 13587 1235
rect 13541 1163 13547 1197
rect 13581 1163 13587 1197
rect 13541 1125 13587 1163
rect 13541 1091 13547 1125
rect 13581 1091 13587 1125
rect 13541 1053 13587 1091
rect 13541 1019 13547 1053
rect 13581 1019 13587 1053
rect 13541 981 13587 1019
rect 13541 947 13547 981
rect 13581 947 13587 981
rect 13541 909 13587 947
rect 13541 875 13547 909
rect 13581 875 13587 909
rect 13541 837 13587 875
rect 13541 803 13547 837
rect 13581 803 13587 837
rect 13541 765 13587 803
rect 13541 731 13547 765
rect 13581 731 13587 765
rect 13541 693 13587 731
rect 13541 659 13547 693
rect 13581 659 13587 693
rect 13541 621 13587 659
rect 13541 587 13547 621
rect 13581 587 13587 621
rect 13541 549 13587 587
rect 13541 515 13547 549
rect 13581 515 13587 549
rect 13541 477 13587 515
rect 13541 443 13547 477
rect 13581 443 13587 477
rect 13541 405 13587 443
rect 13541 371 13547 405
rect 13581 371 13587 405
rect 13541 355 13587 371
rect 13999 1629 14045 1645
rect 13999 1595 14005 1629
rect 14039 1595 14045 1629
rect 13999 1557 14045 1595
rect 13999 1523 14005 1557
rect 14039 1523 14045 1557
rect 13999 1485 14045 1523
rect 13999 1451 14005 1485
rect 14039 1451 14045 1485
rect 13999 1413 14045 1451
rect 13999 1379 14005 1413
rect 14039 1379 14045 1413
rect 13999 1341 14045 1379
rect 13999 1307 14005 1341
rect 14039 1307 14045 1341
rect 13999 1269 14045 1307
rect 13999 1235 14005 1269
rect 14039 1235 14045 1269
rect 13999 1197 14045 1235
rect 13999 1163 14005 1197
rect 14039 1163 14045 1197
rect 13999 1125 14045 1163
rect 13999 1091 14005 1125
rect 14039 1091 14045 1125
rect 13999 1053 14045 1091
rect 13999 1019 14005 1053
rect 14039 1019 14045 1053
rect 13999 981 14045 1019
rect 13999 947 14005 981
rect 14039 947 14045 981
rect 13999 909 14045 947
rect 13999 875 14005 909
rect 14039 875 14045 909
rect 13999 837 14045 875
rect 13999 803 14005 837
rect 14039 803 14045 837
rect 13999 765 14045 803
rect 13999 731 14005 765
rect 14039 731 14045 765
rect 13999 693 14045 731
rect 13999 659 14005 693
rect 14039 659 14045 693
rect 13999 621 14045 659
rect 13999 587 14005 621
rect 14039 587 14045 621
rect 13999 549 14045 587
rect 13999 515 14005 549
rect 14039 515 14045 549
rect 13999 477 14045 515
rect 13999 443 14005 477
rect 14039 443 14045 477
rect 13999 405 14045 443
rect 13999 371 14005 405
rect 14039 371 14045 405
rect 13999 355 14045 371
rect 14457 1629 14503 1645
rect 14457 1595 14463 1629
rect 14497 1595 14503 1629
rect 14457 1557 14503 1595
rect 14457 1523 14463 1557
rect 14497 1523 14503 1557
rect 14457 1485 14503 1523
rect 14457 1451 14463 1485
rect 14497 1451 14503 1485
rect 14457 1413 14503 1451
rect 14457 1379 14463 1413
rect 14497 1379 14503 1413
rect 14457 1341 14503 1379
rect 14457 1307 14463 1341
rect 14497 1307 14503 1341
rect 14457 1269 14503 1307
rect 14457 1235 14463 1269
rect 14497 1235 14503 1269
rect 14457 1197 14503 1235
rect 14457 1163 14463 1197
rect 14497 1163 14503 1197
rect 14457 1125 14503 1163
rect 14457 1091 14463 1125
rect 14497 1091 14503 1125
rect 14457 1053 14503 1091
rect 14457 1019 14463 1053
rect 14497 1019 14503 1053
rect 14457 981 14503 1019
rect 14457 947 14463 981
rect 14497 947 14503 981
rect 14457 909 14503 947
rect 14457 875 14463 909
rect 14497 875 14503 909
rect 14457 837 14503 875
rect 14457 803 14463 837
rect 14497 803 14503 837
rect 14457 765 14503 803
rect 14457 731 14463 765
rect 14497 731 14503 765
rect 14457 693 14503 731
rect 14457 659 14463 693
rect 14497 659 14503 693
rect 14457 621 14503 659
rect 14457 587 14463 621
rect 14497 587 14503 621
rect 14457 549 14503 587
rect 14457 515 14463 549
rect 14497 515 14503 549
rect 14457 477 14503 515
rect 14457 443 14463 477
rect 14497 443 14503 477
rect 14457 405 14503 443
rect 14457 371 14463 405
rect 14497 371 14503 405
rect 14457 355 14503 371
rect 14915 1629 14961 1645
rect 14915 1595 14921 1629
rect 14955 1595 14961 1629
rect 14915 1557 14961 1595
rect 14915 1523 14921 1557
rect 14955 1523 14961 1557
rect 14915 1485 14961 1523
rect 14915 1451 14921 1485
rect 14955 1451 14961 1485
rect 14915 1413 14961 1451
rect 14915 1379 14921 1413
rect 14955 1379 14961 1413
rect 14915 1341 14961 1379
rect 14915 1307 14921 1341
rect 14955 1307 14961 1341
rect 14915 1269 14961 1307
rect 14915 1235 14921 1269
rect 14955 1235 14961 1269
rect 14915 1197 14961 1235
rect 14915 1163 14921 1197
rect 14955 1163 14961 1197
rect 14915 1125 14961 1163
rect 14915 1091 14921 1125
rect 14955 1091 14961 1125
rect 14915 1053 14961 1091
rect 14915 1019 14921 1053
rect 14955 1019 14961 1053
rect 14915 981 14961 1019
rect 14915 947 14921 981
rect 14955 947 14961 981
rect 14915 909 14961 947
rect 14915 875 14921 909
rect 14955 875 14961 909
rect 14915 837 14961 875
rect 14915 803 14921 837
rect 14955 803 14961 837
rect 14915 765 14961 803
rect 14915 731 14921 765
rect 14955 731 14961 765
rect 14915 693 14961 731
rect 14915 659 14921 693
rect 14955 659 14961 693
rect 14915 621 14961 659
rect 14915 587 14921 621
rect 14955 587 14961 621
rect 14915 549 14961 587
rect 14915 515 14921 549
rect 14955 515 14961 549
rect 14915 477 14961 515
rect 14915 443 14921 477
rect 14955 443 14961 477
rect 14915 405 14961 443
rect 14915 371 14921 405
rect 14955 371 14961 405
rect 14915 355 14961 371
rect 15373 1629 15419 1645
rect 15373 1595 15379 1629
rect 15413 1595 15419 1629
rect 15373 1557 15419 1595
rect 15373 1523 15379 1557
rect 15413 1523 15419 1557
rect 15373 1485 15419 1523
rect 15373 1451 15379 1485
rect 15413 1451 15419 1485
rect 15373 1413 15419 1451
rect 15373 1379 15379 1413
rect 15413 1379 15419 1413
rect 15373 1341 15419 1379
rect 15373 1307 15379 1341
rect 15413 1307 15419 1341
rect 15373 1269 15419 1307
rect 15373 1235 15379 1269
rect 15413 1235 15419 1269
rect 15373 1197 15419 1235
rect 15373 1163 15379 1197
rect 15413 1163 15419 1197
rect 15373 1125 15419 1163
rect 15373 1091 15379 1125
rect 15413 1091 15419 1125
rect 15373 1053 15419 1091
rect 15373 1019 15379 1053
rect 15413 1019 15419 1053
rect 15373 981 15419 1019
rect 15373 947 15379 981
rect 15413 947 15419 981
rect 15373 909 15419 947
rect 15373 875 15379 909
rect 15413 875 15419 909
rect 15373 837 15419 875
rect 15373 803 15379 837
rect 15413 803 15419 837
rect 15373 765 15419 803
rect 15373 731 15379 765
rect 15413 731 15419 765
rect 15373 693 15419 731
rect 15373 659 15379 693
rect 15413 659 15419 693
rect 15373 621 15419 659
rect 15373 587 15379 621
rect 15413 587 15419 621
rect 15373 549 15419 587
rect 15373 515 15379 549
rect 15413 515 15419 549
rect 15373 477 15419 515
rect 15373 443 15379 477
rect 15413 443 15419 477
rect 15373 405 15419 443
rect 15373 371 15379 405
rect 15413 371 15419 405
rect 15373 355 15419 371
rect 15831 1629 15877 1645
rect 15831 1595 15837 1629
rect 15871 1595 15877 1629
rect 15831 1557 15877 1595
rect 15831 1523 15837 1557
rect 15871 1523 15877 1557
rect 15831 1485 15877 1523
rect 15831 1451 15837 1485
rect 15871 1451 15877 1485
rect 15831 1413 15877 1451
rect 15831 1379 15837 1413
rect 15871 1379 15877 1413
rect 15831 1341 15877 1379
rect 15831 1307 15837 1341
rect 15871 1307 15877 1341
rect 15831 1269 15877 1307
rect 15831 1235 15837 1269
rect 15871 1235 15877 1269
rect 15831 1197 15877 1235
rect 15831 1163 15837 1197
rect 15871 1163 15877 1197
rect 15831 1125 15877 1163
rect 15831 1091 15837 1125
rect 15871 1091 15877 1125
rect 15831 1053 15877 1091
rect 15831 1019 15837 1053
rect 15871 1019 15877 1053
rect 15831 981 15877 1019
rect 15831 947 15837 981
rect 15871 947 15877 981
rect 15831 909 15877 947
rect 15831 875 15837 909
rect 15871 875 15877 909
rect 15831 837 15877 875
rect 15831 803 15837 837
rect 15871 803 15877 837
rect 15831 765 15877 803
rect 15831 731 15837 765
rect 15871 731 15877 765
rect 15831 693 15877 731
rect 15831 659 15837 693
rect 15871 659 15877 693
rect 15831 621 15877 659
rect 15831 587 15837 621
rect 15871 587 15877 621
rect 15831 549 15877 587
rect 15831 515 15837 549
rect 15871 515 15877 549
rect 15831 477 15877 515
rect 15831 443 15837 477
rect 15871 443 15877 477
rect 15831 405 15877 443
rect 15831 371 15837 405
rect 15871 371 15877 405
rect 15831 355 15877 371
rect 16289 1629 16335 1645
rect 16289 1595 16295 1629
rect 16329 1595 16335 1629
rect 16289 1557 16335 1595
rect 16289 1523 16295 1557
rect 16329 1523 16335 1557
rect 16289 1485 16335 1523
rect 16289 1451 16295 1485
rect 16329 1451 16335 1485
rect 16289 1413 16335 1451
rect 16289 1379 16295 1413
rect 16329 1379 16335 1413
rect 16289 1341 16335 1379
rect 16289 1307 16295 1341
rect 16329 1307 16335 1341
rect 16289 1269 16335 1307
rect 16289 1235 16295 1269
rect 16329 1235 16335 1269
rect 16289 1197 16335 1235
rect 16289 1163 16295 1197
rect 16329 1163 16335 1197
rect 16289 1125 16335 1163
rect 16289 1091 16295 1125
rect 16329 1091 16335 1125
rect 16289 1053 16335 1091
rect 16289 1019 16295 1053
rect 16329 1019 16335 1053
rect 16289 981 16335 1019
rect 16289 947 16295 981
rect 16329 947 16335 981
rect 16289 909 16335 947
rect 16289 875 16295 909
rect 16329 875 16335 909
rect 16289 837 16335 875
rect 16289 803 16295 837
rect 16329 803 16335 837
rect 16289 765 16335 803
rect 16289 731 16295 765
rect 16329 731 16335 765
rect 16289 693 16335 731
rect 16289 659 16295 693
rect 16329 659 16335 693
rect 16289 621 16335 659
rect 16289 587 16295 621
rect 16329 587 16335 621
rect 16289 549 16335 587
rect 16289 515 16295 549
rect 16329 515 16335 549
rect 16289 477 16335 515
rect 16289 443 16295 477
rect 16329 443 16335 477
rect 16289 405 16335 443
rect 16289 371 16295 405
rect 16329 371 16335 405
rect 16289 355 16335 371
rect 16747 1629 16793 1645
rect 16747 1595 16753 1629
rect 16787 1595 16793 1629
rect 16747 1557 16793 1595
rect 16747 1523 16753 1557
rect 16787 1523 16793 1557
rect 16747 1485 16793 1523
rect 16747 1451 16753 1485
rect 16787 1451 16793 1485
rect 16747 1413 16793 1451
rect 16747 1379 16753 1413
rect 16787 1379 16793 1413
rect 16747 1341 16793 1379
rect 16747 1307 16753 1341
rect 16787 1307 16793 1341
rect 16747 1269 16793 1307
rect 16747 1235 16753 1269
rect 16787 1235 16793 1269
rect 16747 1197 16793 1235
rect 16747 1163 16753 1197
rect 16787 1163 16793 1197
rect 16747 1125 16793 1163
rect 16747 1091 16753 1125
rect 16787 1091 16793 1125
rect 16747 1053 16793 1091
rect 16747 1019 16753 1053
rect 16787 1019 16793 1053
rect 16747 981 16793 1019
rect 16747 947 16753 981
rect 16787 947 16793 981
rect 16747 909 16793 947
rect 16747 875 16753 909
rect 16787 875 16793 909
rect 16747 837 16793 875
rect 16747 803 16753 837
rect 16787 803 16793 837
rect 16747 765 16793 803
rect 16747 731 16753 765
rect 16787 731 16793 765
rect 16747 693 16793 731
rect 16747 659 16753 693
rect 16787 659 16793 693
rect 16747 621 16793 659
rect 16747 587 16753 621
rect 16787 587 16793 621
rect 16747 549 16793 587
rect 16747 515 16753 549
rect 16787 515 16793 549
rect 16747 477 16793 515
rect 16747 443 16753 477
rect 16787 443 16793 477
rect 16747 405 16793 443
rect 16747 371 16753 405
rect 16787 371 16793 405
rect 16747 355 16793 371
rect 17205 1629 17251 1645
rect 17205 1595 17211 1629
rect 17245 1595 17251 1629
rect 17205 1557 17251 1595
rect 17205 1523 17211 1557
rect 17245 1523 17251 1557
rect 17205 1485 17251 1523
rect 17205 1451 17211 1485
rect 17245 1451 17251 1485
rect 17205 1413 17251 1451
rect 17205 1379 17211 1413
rect 17245 1379 17251 1413
rect 17205 1341 17251 1379
rect 17205 1307 17211 1341
rect 17245 1307 17251 1341
rect 17205 1269 17251 1307
rect 17205 1235 17211 1269
rect 17245 1235 17251 1269
rect 17205 1197 17251 1235
rect 17205 1163 17211 1197
rect 17245 1163 17251 1197
rect 17205 1125 17251 1163
rect 17205 1091 17211 1125
rect 17245 1091 17251 1125
rect 17205 1053 17251 1091
rect 17205 1019 17211 1053
rect 17245 1019 17251 1053
rect 17205 981 17251 1019
rect 17205 947 17211 981
rect 17245 947 17251 981
rect 17205 909 17251 947
rect 17205 875 17211 909
rect 17245 875 17251 909
rect 17205 837 17251 875
rect 17205 803 17211 837
rect 17245 803 17251 837
rect 17205 765 17251 803
rect 17205 731 17211 765
rect 17245 731 17251 765
rect 17205 693 17251 731
rect 17205 659 17211 693
rect 17245 659 17251 693
rect 17205 621 17251 659
rect 17205 587 17211 621
rect 17245 587 17251 621
rect 17205 549 17251 587
rect 17205 515 17211 549
rect 17245 515 17251 549
rect 17205 477 17251 515
rect 17205 443 17211 477
rect 17245 443 17251 477
rect 17205 405 17251 443
rect 17205 371 17211 405
rect 17245 371 17251 405
rect 17205 355 17251 371
rect 17663 1629 17709 1645
rect 17663 1595 17669 1629
rect 17703 1595 17709 1629
rect 17663 1557 17709 1595
rect 17663 1523 17669 1557
rect 17703 1523 17709 1557
rect 17663 1485 17709 1523
rect 17663 1451 17669 1485
rect 17703 1451 17709 1485
rect 17663 1413 17709 1451
rect 17663 1379 17669 1413
rect 17703 1379 17709 1413
rect 17663 1341 17709 1379
rect 17663 1307 17669 1341
rect 17703 1307 17709 1341
rect 17663 1269 17709 1307
rect 17663 1235 17669 1269
rect 17703 1235 17709 1269
rect 17663 1197 17709 1235
rect 17663 1163 17669 1197
rect 17703 1163 17709 1197
rect 17663 1125 17709 1163
rect 17663 1091 17669 1125
rect 17703 1091 17709 1125
rect 17663 1053 17709 1091
rect 17663 1019 17669 1053
rect 17703 1019 17709 1053
rect 17663 981 17709 1019
rect 17663 947 17669 981
rect 17703 947 17709 981
rect 17663 909 17709 947
rect 17663 875 17669 909
rect 17703 875 17709 909
rect 17663 837 17709 875
rect 17663 803 17669 837
rect 17703 803 17709 837
rect 17663 765 17709 803
rect 17663 731 17669 765
rect 17703 731 17709 765
rect 17663 693 17709 731
rect 17663 659 17669 693
rect 17703 659 17709 693
rect 17663 621 17709 659
rect 17663 587 17669 621
rect 17703 587 17709 621
rect 17663 549 17709 587
rect 17663 515 17669 549
rect 17703 515 17709 549
rect 17663 477 17709 515
rect 17663 443 17669 477
rect 17703 443 17709 477
rect 17663 405 17709 443
rect 17663 371 17669 405
rect 17703 371 17709 405
rect 17663 355 17709 371
rect 18121 1629 18167 1645
rect 18121 1595 18127 1629
rect 18161 1595 18167 1629
rect 18121 1557 18167 1595
rect 18121 1523 18127 1557
rect 18161 1523 18167 1557
rect 18121 1485 18167 1523
rect 18121 1451 18127 1485
rect 18161 1451 18167 1485
rect 18121 1413 18167 1451
rect 18121 1379 18127 1413
rect 18161 1379 18167 1413
rect 18121 1341 18167 1379
rect 18121 1307 18127 1341
rect 18161 1307 18167 1341
rect 18121 1269 18167 1307
rect 18121 1235 18127 1269
rect 18161 1235 18167 1269
rect 18121 1197 18167 1235
rect 18121 1163 18127 1197
rect 18161 1163 18167 1197
rect 18121 1125 18167 1163
rect 18121 1091 18127 1125
rect 18161 1091 18167 1125
rect 18121 1053 18167 1091
rect 18121 1019 18127 1053
rect 18161 1019 18167 1053
rect 18121 981 18167 1019
rect 18121 947 18127 981
rect 18161 947 18167 981
rect 18121 909 18167 947
rect 18121 875 18127 909
rect 18161 875 18167 909
rect 18121 837 18167 875
rect 18121 803 18127 837
rect 18161 803 18167 837
rect 18121 765 18167 803
rect 18121 731 18127 765
rect 18161 731 18167 765
rect 18121 693 18167 731
rect 18121 659 18127 693
rect 18161 659 18167 693
rect 18121 621 18167 659
rect 18121 587 18127 621
rect 18161 587 18167 621
rect 18121 549 18167 587
rect 18121 515 18127 549
rect 18161 515 18167 549
rect 18121 477 18167 515
rect 18121 443 18127 477
rect 18161 443 18167 477
rect 18121 405 18167 443
rect 18121 371 18127 405
rect 18161 371 18167 405
rect 18121 355 18167 371
rect 18579 1629 18625 1645
rect 18579 1595 18585 1629
rect 18619 1595 18625 1629
rect 18579 1557 18625 1595
rect 18579 1523 18585 1557
rect 18619 1523 18625 1557
rect 18579 1485 18625 1523
rect 18579 1451 18585 1485
rect 18619 1451 18625 1485
rect 18579 1413 18625 1451
rect 18579 1379 18585 1413
rect 18619 1379 18625 1413
rect 18579 1341 18625 1379
rect 18579 1307 18585 1341
rect 18619 1307 18625 1341
rect 18579 1269 18625 1307
rect 18579 1235 18585 1269
rect 18619 1235 18625 1269
rect 18579 1197 18625 1235
rect 18579 1163 18585 1197
rect 18619 1163 18625 1197
rect 18579 1125 18625 1163
rect 18579 1091 18585 1125
rect 18619 1091 18625 1125
rect 18579 1053 18625 1091
rect 18579 1019 18585 1053
rect 18619 1019 18625 1053
rect 18579 981 18625 1019
rect 18579 947 18585 981
rect 18619 947 18625 981
rect 18579 909 18625 947
rect 18579 875 18585 909
rect 18619 875 18625 909
rect 18579 837 18625 875
rect 18579 803 18585 837
rect 18619 803 18625 837
rect 18579 765 18625 803
rect 18579 731 18585 765
rect 18619 731 18625 765
rect 18579 693 18625 731
rect 18579 659 18585 693
rect 18619 659 18625 693
rect 18579 621 18625 659
rect 18579 587 18585 621
rect 18619 587 18625 621
rect 18579 549 18625 587
rect 18579 515 18585 549
rect 18619 515 18625 549
rect 18579 477 18625 515
rect 18579 443 18585 477
rect 18619 443 18625 477
rect 18579 405 18625 443
rect 18579 371 18585 405
rect 18619 371 18625 405
rect 18579 355 18625 371
rect 19037 1629 19083 1645
rect 19037 1595 19043 1629
rect 19077 1595 19083 1629
rect 19037 1557 19083 1595
rect 19037 1523 19043 1557
rect 19077 1523 19083 1557
rect 19037 1485 19083 1523
rect 19037 1451 19043 1485
rect 19077 1451 19083 1485
rect 19037 1413 19083 1451
rect 19037 1379 19043 1413
rect 19077 1379 19083 1413
rect 19037 1341 19083 1379
rect 19037 1307 19043 1341
rect 19077 1307 19083 1341
rect 19037 1269 19083 1307
rect 19037 1235 19043 1269
rect 19077 1235 19083 1269
rect 19037 1197 19083 1235
rect 19037 1163 19043 1197
rect 19077 1163 19083 1197
rect 19037 1125 19083 1163
rect 19037 1091 19043 1125
rect 19077 1091 19083 1125
rect 19037 1053 19083 1091
rect 19037 1019 19043 1053
rect 19077 1019 19083 1053
rect 19037 981 19083 1019
rect 19037 947 19043 981
rect 19077 947 19083 981
rect 19037 909 19083 947
rect 19037 875 19043 909
rect 19077 875 19083 909
rect 19037 837 19083 875
rect 19037 803 19043 837
rect 19077 803 19083 837
rect 19037 765 19083 803
rect 19037 731 19043 765
rect 19077 731 19083 765
rect 19037 693 19083 731
rect 19037 659 19043 693
rect 19077 659 19083 693
rect 19037 621 19083 659
rect 19037 587 19043 621
rect 19077 587 19083 621
rect 19037 549 19083 587
rect 19037 515 19043 549
rect 19077 515 19083 549
rect 19037 477 19083 515
rect 19037 443 19043 477
rect 19077 443 19083 477
rect 19037 405 19083 443
rect 19037 371 19043 405
rect 19077 371 19083 405
rect 19037 355 19083 371
rect 19495 1629 19541 1645
rect 19495 1595 19501 1629
rect 19535 1595 19541 1629
rect 19495 1557 19541 1595
rect 19495 1523 19501 1557
rect 19535 1523 19541 1557
rect 19495 1485 19541 1523
rect 19495 1451 19501 1485
rect 19535 1451 19541 1485
rect 19495 1413 19541 1451
rect 19495 1379 19501 1413
rect 19535 1379 19541 1413
rect 19495 1341 19541 1379
rect 19495 1307 19501 1341
rect 19535 1307 19541 1341
rect 19495 1269 19541 1307
rect 19495 1235 19501 1269
rect 19535 1235 19541 1269
rect 19495 1197 19541 1235
rect 19495 1163 19501 1197
rect 19535 1163 19541 1197
rect 19495 1125 19541 1163
rect 19495 1091 19501 1125
rect 19535 1091 19541 1125
rect 19495 1053 19541 1091
rect 19495 1019 19501 1053
rect 19535 1019 19541 1053
rect 19495 981 19541 1019
rect 19495 947 19501 981
rect 19535 947 19541 981
rect 19495 909 19541 947
rect 19495 875 19501 909
rect 19535 875 19541 909
rect 19495 837 19541 875
rect 19495 803 19501 837
rect 19535 803 19541 837
rect 19495 765 19541 803
rect 19495 731 19501 765
rect 19535 731 19541 765
rect 19495 693 19541 731
rect 19495 659 19501 693
rect 19535 659 19541 693
rect 19495 621 19541 659
rect 19495 587 19501 621
rect 19535 587 19541 621
rect 19495 549 19541 587
rect 19495 515 19501 549
rect 19535 515 19541 549
rect 19495 477 19541 515
rect 19495 443 19501 477
rect 19535 443 19541 477
rect 19495 405 19541 443
rect 19495 371 19501 405
rect 19535 371 19541 405
rect 19495 355 19541 371
rect 19953 1629 19999 1645
rect 19953 1595 19959 1629
rect 19993 1595 19999 1629
rect 19953 1557 19999 1595
rect 19953 1523 19959 1557
rect 19993 1523 19999 1557
rect 19953 1485 19999 1523
rect 19953 1451 19959 1485
rect 19993 1451 19999 1485
rect 19953 1413 19999 1451
rect 19953 1379 19959 1413
rect 19993 1379 19999 1413
rect 19953 1341 19999 1379
rect 19953 1307 19959 1341
rect 19993 1307 19999 1341
rect 19953 1269 19999 1307
rect 19953 1235 19959 1269
rect 19993 1235 19999 1269
rect 19953 1197 19999 1235
rect 19953 1163 19959 1197
rect 19993 1163 19999 1197
rect 19953 1125 19999 1163
rect 19953 1091 19959 1125
rect 19993 1091 19999 1125
rect 19953 1053 19999 1091
rect 19953 1019 19959 1053
rect 19993 1019 19999 1053
rect 19953 981 19999 1019
rect 19953 947 19959 981
rect 19993 947 19999 981
rect 19953 909 19999 947
rect 19953 875 19959 909
rect 19993 875 19999 909
rect 19953 837 19999 875
rect 19953 803 19959 837
rect 19993 803 19999 837
rect 19953 765 19999 803
rect 19953 731 19959 765
rect 19993 731 19999 765
rect 19953 693 19999 731
rect 19953 659 19959 693
rect 19993 659 19999 693
rect 19953 621 19999 659
rect 19953 587 19959 621
rect 19993 587 19999 621
rect 19953 549 19999 587
rect 19953 515 19959 549
rect 19993 515 19999 549
rect 19953 477 19999 515
rect 19953 443 19959 477
rect 19993 443 19999 477
rect 19953 405 19999 443
rect 19953 371 19959 405
rect 19993 371 19999 405
rect 19953 355 19999 371
rect 20411 1629 20457 1645
rect 20411 1595 20417 1629
rect 20451 1595 20457 1629
rect 20411 1557 20457 1595
rect 20411 1523 20417 1557
rect 20451 1523 20457 1557
rect 20411 1485 20457 1523
rect 20411 1451 20417 1485
rect 20451 1451 20457 1485
rect 20411 1413 20457 1451
rect 20411 1379 20417 1413
rect 20451 1379 20457 1413
rect 20411 1341 20457 1379
rect 20411 1307 20417 1341
rect 20451 1307 20457 1341
rect 20411 1269 20457 1307
rect 20411 1235 20417 1269
rect 20451 1235 20457 1269
rect 20411 1197 20457 1235
rect 20411 1163 20417 1197
rect 20451 1163 20457 1197
rect 20411 1125 20457 1163
rect 20411 1091 20417 1125
rect 20451 1091 20457 1125
rect 20411 1053 20457 1091
rect 20411 1019 20417 1053
rect 20451 1019 20457 1053
rect 20411 981 20457 1019
rect 20411 947 20417 981
rect 20451 947 20457 981
rect 20411 909 20457 947
rect 20411 875 20417 909
rect 20451 875 20457 909
rect 20411 837 20457 875
rect 20411 803 20417 837
rect 20451 803 20457 837
rect 20411 765 20457 803
rect 20411 731 20417 765
rect 20451 731 20457 765
rect 20411 693 20457 731
rect 20411 659 20417 693
rect 20451 659 20457 693
rect 20411 621 20457 659
rect 20411 587 20417 621
rect 20451 587 20457 621
rect 20411 549 20457 587
rect 20411 515 20417 549
rect 20451 515 20457 549
rect 20411 477 20457 515
rect 20411 443 20417 477
rect 20451 443 20457 477
rect 20411 405 20457 443
rect 20411 371 20417 405
rect 20451 371 20457 405
rect 20411 355 20457 371
rect 20869 1629 20915 1645
rect 20869 1595 20875 1629
rect 20909 1595 20915 1629
rect 20869 1557 20915 1595
rect 20869 1523 20875 1557
rect 20909 1523 20915 1557
rect 20869 1485 20915 1523
rect 20869 1451 20875 1485
rect 20909 1451 20915 1485
rect 20869 1413 20915 1451
rect 20869 1379 20875 1413
rect 20909 1379 20915 1413
rect 20869 1341 20915 1379
rect 20869 1307 20875 1341
rect 20909 1307 20915 1341
rect 20869 1269 20915 1307
rect 20869 1235 20875 1269
rect 20909 1235 20915 1269
rect 20869 1197 20915 1235
rect 20869 1163 20875 1197
rect 20909 1163 20915 1197
rect 20869 1125 20915 1163
rect 20869 1091 20875 1125
rect 20909 1091 20915 1125
rect 20869 1053 20915 1091
rect 20869 1019 20875 1053
rect 20909 1019 20915 1053
rect 20869 981 20915 1019
rect 20869 947 20875 981
rect 20909 947 20915 981
rect 20869 909 20915 947
rect 20869 875 20875 909
rect 20909 875 20915 909
rect 20869 837 20915 875
rect 20869 803 20875 837
rect 20909 803 20915 837
rect 20869 765 20915 803
rect 20869 731 20875 765
rect 20909 731 20915 765
rect 20869 693 20915 731
rect 20869 659 20875 693
rect 20909 659 20915 693
rect 20869 621 20915 659
rect 20869 587 20875 621
rect 20909 587 20915 621
rect 20869 549 20915 587
rect 20869 515 20875 549
rect 20909 515 20915 549
rect 20869 477 20915 515
rect 20869 443 20875 477
rect 20909 443 20915 477
rect 20869 405 20915 443
rect 20869 371 20875 405
rect 20909 371 20915 405
rect 20869 355 20915 371
rect 21327 1629 21373 1645
rect 21327 1595 21333 1629
rect 21367 1595 21373 1629
rect 21327 1557 21373 1595
rect 21327 1523 21333 1557
rect 21367 1523 21373 1557
rect 21327 1485 21373 1523
rect 21327 1451 21333 1485
rect 21367 1451 21373 1485
rect 21327 1413 21373 1451
rect 21327 1379 21333 1413
rect 21367 1379 21373 1413
rect 21327 1341 21373 1379
rect 21327 1307 21333 1341
rect 21367 1307 21373 1341
rect 21327 1269 21373 1307
rect 21327 1235 21333 1269
rect 21367 1235 21373 1269
rect 21327 1197 21373 1235
rect 21327 1163 21333 1197
rect 21367 1163 21373 1197
rect 21327 1125 21373 1163
rect 21327 1091 21333 1125
rect 21367 1091 21373 1125
rect 21327 1053 21373 1091
rect 21327 1019 21333 1053
rect 21367 1019 21373 1053
rect 21327 981 21373 1019
rect 21327 947 21333 981
rect 21367 947 21373 981
rect 21327 909 21373 947
rect 21327 875 21333 909
rect 21367 875 21373 909
rect 21327 837 21373 875
rect 21327 803 21333 837
rect 21367 803 21373 837
rect 21327 765 21373 803
rect 21327 731 21333 765
rect 21367 731 21373 765
rect 21327 693 21373 731
rect 21327 659 21333 693
rect 21367 659 21373 693
rect 21327 621 21373 659
rect 21327 587 21333 621
rect 21367 587 21373 621
rect 21327 549 21373 587
rect 21327 515 21333 549
rect 21367 515 21373 549
rect 21327 477 21373 515
rect 21327 443 21333 477
rect 21367 443 21373 477
rect 21327 405 21373 443
rect 21327 371 21333 405
rect 21367 371 21373 405
rect 21327 355 21373 371
rect 21785 1629 21831 1645
rect 21785 1595 21791 1629
rect 21825 1595 21831 1629
rect 21785 1557 21831 1595
rect 21785 1523 21791 1557
rect 21825 1523 21831 1557
rect 21785 1485 21831 1523
rect 21785 1451 21791 1485
rect 21825 1451 21831 1485
rect 21785 1413 21831 1451
rect 21785 1379 21791 1413
rect 21825 1379 21831 1413
rect 21785 1341 21831 1379
rect 21785 1307 21791 1341
rect 21825 1307 21831 1341
rect 21785 1269 21831 1307
rect 21785 1235 21791 1269
rect 21825 1235 21831 1269
rect 21785 1197 21831 1235
rect 21785 1163 21791 1197
rect 21825 1163 21831 1197
rect 21785 1125 21831 1163
rect 21785 1091 21791 1125
rect 21825 1091 21831 1125
rect 21785 1053 21831 1091
rect 21785 1019 21791 1053
rect 21825 1019 21831 1053
rect 21785 981 21831 1019
rect 21785 947 21791 981
rect 21825 947 21831 981
rect 21785 909 21831 947
rect 21785 875 21791 909
rect 21825 875 21831 909
rect 21785 837 21831 875
rect 21785 803 21791 837
rect 21825 803 21831 837
rect 21785 765 21831 803
rect 21785 731 21791 765
rect 21825 731 21831 765
rect 21785 693 21831 731
rect 21785 659 21791 693
rect 21825 659 21831 693
rect 21785 621 21831 659
rect 21785 587 21791 621
rect 21825 587 21831 621
rect 21785 549 21831 587
rect 21785 515 21791 549
rect 21825 515 21831 549
rect 21785 477 21831 515
rect 21785 443 21791 477
rect 21825 443 21831 477
rect 21785 405 21831 443
rect 21785 371 21791 405
rect 21825 371 21831 405
rect 21785 355 21831 371
rect 22243 1629 22289 1645
rect 22243 1595 22249 1629
rect 22283 1595 22289 1629
rect 22243 1557 22289 1595
rect 22243 1523 22249 1557
rect 22283 1523 22289 1557
rect 22243 1485 22289 1523
rect 22243 1451 22249 1485
rect 22283 1451 22289 1485
rect 22243 1413 22289 1451
rect 22243 1379 22249 1413
rect 22283 1379 22289 1413
rect 22243 1341 22289 1379
rect 22243 1307 22249 1341
rect 22283 1307 22289 1341
rect 22243 1269 22289 1307
rect 22243 1235 22249 1269
rect 22283 1235 22289 1269
rect 22243 1197 22289 1235
rect 22243 1163 22249 1197
rect 22283 1163 22289 1197
rect 22243 1125 22289 1163
rect 22243 1091 22249 1125
rect 22283 1091 22289 1125
rect 22243 1053 22289 1091
rect 22243 1019 22249 1053
rect 22283 1019 22289 1053
rect 22243 981 22289 1019
rect 22243 947 22249 981
rect 22283 947 22289 981
rect 22243 909 22289 947
rect 22243 875 22249 909
rect 22283 875 22289 909
rect 22243 837 22289 875
rect 22243 803 22249 837
rect 22283 803 22289 837
rect 22243 765 22289 803
rect 22243 731 22249 765
rect 22283 731 22289 765
rect 22243 693 22289 731
rect 22243 659 22249 693
rect 22283 659 22289 693
rect 22243 621 22289 659
rect 22243 587 22249 621
rect 22283 587 22289 621
rect 22243 549 22289 587
rect 22243 515 22249 549
rect 22283 515 22289 549
rect 22243 477 22289 515
rect 22243 443 22249 477
rect 22283 443 22289 477
rect 22243 405 22289 443
rect 22243 371 22249 405
rect 22283 371 22289 405
rect 22243 355 22289 371
rect 22701 1629 22747 1645
rect 22701 1595 22707 1629
rect 22741 1595 22747 1629
rect 22701 1557 22747 1595
rect 22701 1523 22707 1557
rect 22741 1523 22747 1557
rect 22701 1485 22747 1523
rect 22701 1451 22707 1485
rect 22741 1451 22747 1485
rect 22701 1413 22747 1451
rect 22701 1379 22707 1413
rect 22741 1379 22747 1413
rect 22701 1341 22747 1379
rect 22701 1307 22707 1341
rect 22741 1307 22747 1341
rect 22701 1269 22747 1307
rect 22701 1235 22707 1269
rect 22741 1235 22747 1269
rect 22701 1197 22747 1235
rect 22701 1163 22707 1197
rect 22741 1163 22747 1197
rect 22701 1125 22747 1163
rect 22701 1091 22707 1125
rect 22741 1091 22747 1125
rect 22701 1053 22747 1091
rect 22701 1019 22707 1053
rect 22741 1019 22747 1053
rect 22701 981 22747 1019
rect 22701 947 22707 981
rect 22741 947 22747 981
rect 22701 909 22747 947
rect 22701 875 22707 909
rect 22741 875 22747 909
rect 22701 837 22747 875
rect 22701 803 22707 837
rect 22741 803 22747 837
rect 22701 765 22747 803
rect 22701 731 22707 765
rect 22741 731 22747 765
rect 22701 693 22747 731
rect 22701 659 22707 693
rect 22741 659 22747 693
rect 22701 621 22747 659
rect 22701 587 22707 621
rect 22741 587 22747 621
rect 22701 549 22747 587
rect 22701 515 22707 549
rect 22741 515 22747 549
rect 22701 477 22747 515
rect 22701 443 22707 477
rect 22741 443 22747 477
rect 22701 405 22747 443
rect 22701 371 22707 405
rect 22741 371 22747 405
rect 22701 355 22747 371
rect 23159 1629 23205 1645
rect 23159 1595 23165 1629
rect 23199 1595 23205 1629
rect 23159 1557 23205 1595
rect 23159 1523 23165 1557
rect 23199 1523 23205 1557
rect 23159 1485 23205 1523
rect 23159 1451 23165 1485
rect 23199 1451 23205 1485
rect 23159 1413 23205 1451
rect 23159 1379 23165 1413
rect 23199 1379 23205 1413
rect 23159 1341 23205 1379
rect 23159 1307 23165 1341
rect 23199 1307 23205 1341
rect 23159 1269 23205 1307
rect 23159 1235 23165 1269
rect 23199 1235 23205 1269
rect 23159 1197 23205 1235
rect 23159 1163 23165 1197
rect 23199 1163 23205 1197
rect 23159 1125 23205 1163
rect 23159 1091 23165 1125
rect 23199 1091 23205 1125
rect 23159 1053 23205 1091
rect 23159 1019 23165 1053
rect 23199 1019 23205 1053
rect 23159 981 23205 1019
rect 23159 947 23165 981
rect 23199 947 23205 981
rect 23159 909 23205 947
rect 23159 875 23165 909
rect 23199 875 23205 909
rect 23159 837 23205 875
rect 23159 803 23165 837
rect 23199 803 23205 837
rect 23159 765 23205 803
rect 23159 731 23165 765
rect 23199 731 23205 765
rect 23159 693 23205 731
rect 23159 659 23165 693
rect 23199 659 23205 693
rect 23159 621 23205 659
rect 23159 587 23165 621
rect 23199 587 23205 621
rect 23159 549 23205 587
rect 23159 515 23165 549
rect 23199 515 23205 549
rect 23159 477 23205 515
rect 23159 443 23165 477
rect 23199 443 23205 477
rect 23159 405 23205 443
rect 23159 371 23165 405
rect 23199 371 23205 405
rect 23159 355 23205 371
rect 23617 1629 23663 1645
rect 23617 1595 23623 1629
rect 23657 1595 23663 1629
rect 23617 1557 23663 1595
rect 23617 1523 23623 1557
rect 23657 1523 23663 1557
rect 23617 1485 23663 1523
rect 23617 1451 23623 1485
rect 23657 1451 23663 1485
rect 23617 1413 23663 1451
rect 23617 1379 23623 1413
rect 23657 1379 23663 1413
rect 23617 1341 23663 1379
rect 23617 1307 23623 1341
rect 23657 1307 23663 1341
rect 23617 1269 23663 1307
rect 23617 1235 23623 1269
rect 23657 1235 23663 1269
rect 23617 1197 23663 1235
rect 23617 1163 23623 1197
rect 23657 1163 23663 1197
rect 23617 1125 23663 1163
rect 23617 1091 23623 1125
rect 23657 1091 23663 1125
rect 23617 1053 23663 1091
rect 23617 1019 23623 1053
rect 23657 1019 23663 1053
rect 23617 981 23663 1019
rect 23617 947 23623 981
rect 23657 947 23663 981
rect 23617 909 23663 947
rect 23617 875 23623 909
rect 23657 875 23663 909
rect 23617 837 23663 875
rect 23617 803 23623 837
rect 23657 803 23663 837
rect 23617 765 23663 803
rect 23617 731 23623 765
rect 23657 731 23663 765
rect 23617 693 23663 731
rect 23617 659 23623 693
rect 23657 659 23663 693
rect 23617 621 23663 659
rect 23617 587 23623 621
rect 23657 587 23663 621
rect 23617 549 23663 587
rect 23617 515 23623 549
rect 23657 515 23663 549
rect 23617 477 23663 515
rect 23617 443 23623 477
rect 23657 443 23663 477
rect 23617 405 23663 443
rect 23617 371 23623 405
rect 23657 371 23663 405
rect 23617 355 23663 371
rect 24075 1629 24121 1645
rect 24075 1595 24081 1629
rect 24115 1595 24121 1629
rect 24075 1557 24121 1595
rect 24075 1523 24081 1557
rect 24115 1523 24121 1557
rect 24075 1485 24121 1523
rect 24075 1451 24081 1485
rect 24115 1451 24121 1485
rect 24075 1413 24121 1451
rect 24075 1379 24081 1413
rect 24115 1379 24121 1413
rect 24075 1341 24121 1379
rect 24075 1307 24081 1341
rect 24115 1307 24121 1341
rect 24075 1269 24121 1307
rect 24075 1235 24081 1269
rect 24115 1235 24121 1269
rect 24075 1197 24121 1235
rect 24075 1163 24081 1197
rect 24115 1163 24121 1197
rect 24075 1125 24121 1163
rect 24075 1091 24081 1125
rect 24115 1091 24121 1125
rect 24075 1053 24121 1091
rect 24075 1019 24081 1053
rect 24115 1019 24121 1053
rect 24075 981 24121 1019
rect 24075 947 24081 981
rect 24115 947 24121 981
rect 24075 909 24121 947
rect 24075 875 24081 909
rect 24115 875 24121 909
rect 24075 837 24121 875
rect 24075 803 24081 837
rect 24115 803 24121 837
rect 24075 765 24121 803
rect 24075 731 24081 765
rect 24115 731 24121 765
rect 24075 693 24121 731
rect 24075 659 24081 693
rect 24115 659 24121 693
rect 24075 621 24121 659
rect 24075 587 24081 621
rect 24115 587 24121 621
rect 24075 549 24121 587
rect 24075 515 24081 549
rect 24115 515 24121 549
rect 24075 477 24121 515
rect 24075 443 24081 477
rect 24115 443 24121 477
rect 24075 405 24121 443
rect 24075 371 24081 405
rect 24115 371 24121 405
rect 24075 355 24121 371
rect 24533 1629 24579 1645
rect 24533 1595 24539 1629
rect 24573 1595 24579 1629
rect 24533 1557 24579 1595
rect 24533 1523 24539 1557
rect 24573 1523 24579 1557
rect 24533 1485 24579 1523
rect 24533 1451 24539 1485
rect 24573 1451 24579 1485
rect 24533 1413 24579 1451
rect 24533 1379 24539 1413
rect 24573 1379 24579 1413
rect 24533 1341 24579 1379
rect 24533 1307 24539 1341
rect 24573 1307 24579 1341
rect 24533 1269 24579 1307
rect 24533 1235 24539 1269
rect 24573 1235 24579 1269
rect 24533 1197 24579 1235
rect 24533 1163 24539 1197
rect 24573 1163 24579 1197
rect 24533 1125 24579 1163
rect 24533 1091 24539 1125
rect 24573 1091 24579 1125
rect 24533 1053 24579 1091
rect 24533 1019 24539 1053
rect 24573 1019 24579 1053
rect 24533 981 24579 1019
rect 24533 947 24539 981
rect 24573 947 24579 981
rect 24533 909 24579 947
rect 24533 875 24539 909
rect 24573 875 24579 909
rect 24533 837 24579 875
rect 24533 803 24539 837
rect 24573 803 24579 837
rect 24533 765 24579 803
rect 24533 731 24539 765
rect 24573 731 24579 765
rect 24533 693 24579 731
rect 24533 659 24539 693
rect 24573 659 24579 693
rect 24533 621 24579 659
rect 24533 587 24539 621
rect 24573 587 24579 621
rect 24533 549 24579 587
rect 24533 515 24539 549
rect 24573 515 24579 549
rect 24533 477 24579 515
rect 24533 443 24539 477
rect 24573 443 24579 477
rect 24533 405 24579 443
rect 24533 371 24539 405
rect 24573 371 24579 405
rect 24533 355 24579 371
rect 24991 1629 25037 1645
rect 24991 1595 24997 1629
rect 25031 1595 25037 1629
rect 24991 1557 25037 1595
rect 24991 1523 24997 1557
rect 25031 1523 25037 1557
rect 24991 1485 25037 1523
rect 24991 1451 24997 1485
rect 25031 1451 25037 1485
rect 24991 1413 25037 1451
rect 24991 1379 24997 1413
rect 25031 1379 25037 1413
rect 24991 1341 25037 1379
rect 24991 1307 24997 1341
rect 25031 1307 25037 1341
rect 24991 1269 25037 1307
rect 24991 1235 24997 1269
rect 25031 1235 25037 1269
rect 24991 1197 25037 1235
rect 24991 1163 24997 1197
rect 25031 1163 25037 1197
rect 24991 1125 25037 1163
rect 24991 1091 24997 1125
rect 25031 1091 25037 1125
rect 24991 1053 25037 1091
rect 24991 1019 24997 1053
rect 25031 1019 25037 1053
rect 24991 981 25037 1019
rect 24991 947 24997 981
rect 25031 947 25037 981
rect 24991 909 25037 947
rect 24991 875 24997 909
rect 25031 875 25037 909
rect 24991 837 25037 875
rect 24991 803 24997 837
rect 25031 803 25037 837
rect 24991 765 25037 803
rect 24991 731 24997 765
rect 25031 731 25037 765
rect 24991 693 25037 731
rect 24991 659 24997 693
rect 25031 659 25037 693
rect 24991 621 25037 659
rect 24991 587 24997 621
rect 25031 587 25037 621
rect 24991 549 25037 587
rect 24991 515 24997 549
rect 25031 515 25037 549
rect 24991 477 25037 515
rect 24991 443 24997 477
rect 25031 443 25037 477
rect 24991 405 25037 443
rect 24991 371 24997 405
rect 25031 371 25037 405
rect 24991 355 25037 371
rect 25449 1629 25495 1645
rect 25449 1595 25455 1629
rect 25489 1595 25495 1629
rect 25449 1557 25495 1595
rect 25449 1523 25455 1557
rect 25489 1523 25495 1557
rect 25449 1485 25495 1523
rect 25449 1451 25455 1485
rect 25489 1451 25495 1485
rect 25449 1413 25495 1451
rect 25449 1379 25455 1413
rect 25489 1379 25495 1413
rect 25449 1341 25495 1379
rect 25449 1307 25455 1341
rect 25489 1307 25495 1341
rect 25449 1269 25495 1307
rect 25449 1235 25455 1269
rect 25489 1235 25495 1269
rect 25449 1197 25495 1235
rect 25449 1163 25455 1197
rect 25489 1163 25495 1197
rect 25449 1125 25495 1163
rect 25449 1091 25455 1125
rect 25489 1091 25495 1125
rect 25449 1053 25495 1091
rect 25449 1019 25455 1053
rect 25489 1019 25495 1053
rect 25449 981 25495 1019
rect 25449 947 25455 981
rect 25489 947 25495 981
rect 25449 909 25495 947
rect 25449 875 25455 909
rect 25489 875 25495 909
rect 25449 837 25495 875
rect 25449 803 25455 837
rect 25489 803 25495 837
rect 25449 765 25495 803
rect 25449 731 25455 765
rect 25489 731 25495 765
rect 25449 693 25495 731
rect 25449 659 25455 693
rect 25489 659 25495 693
rect 25449 621 25495 659
rect 25449 587 25455 621
rect 25489 587 25495 621
rect 25449 549 25495 587
rect 25449 515 25455 549
rect 25489 515 25495 549
rect 25449 477 25495 515
rect 25449 443 25455 477
rect 25489 443 25495 477
rect 25449 405 25495 443
rect 25449 371 25455 405
rect 25489 371 25495 405
rect 25449 355 25495 371
rect 25907 1629 25953 1645
rect 25907 1595 25913 1629
rect 25947 1595 25953 1629
rect 25907 1557 25953 1595
rect 25907 1523 25913 1557
rect 25947 1523 25953 1557
rect 25907 1485 25953 1523
rect 25907 1451 25913 1485
rect 25947 1451 25953 1485
rect 25907 1413 25953 1451
rect 25907 1379 25913 1413
rect 25947 1379 25953 1413
rect 25907 1341 25953 1379
rect 25907 1307 25913 1341
rect 25947 1307 25953 1341
rect 25907 1269 25953 1307
rect 25907 1235 25913 1269
rect 25947 1235 25953 1269
rect 25907 1197 25953 1235
rect 25907 1163 25913 1197
rect 25947 1163 25953 1197
rect 25907 1125 25953 1163
rect 25907 1091 25913 1125
rect 25947 1091 25953 1125
rect 25907 1053 25953 1091
rect 25907 1019 25913 1053
rect 25947 1019 25953 1053
rect 25907 981 25953 1019
rect 25907 947 25913 981
rect 25947 947 25953 981
rect 25907 909 25953 947
rect 25907 875 25913 909
rect 25947 875 25953 909
rect 25907 837 25953 875
rect 25907 803 25913 837
rect 25947 803 25953 837
rect 25907 765 25953 803
rect 25907 731 25913 765
rect 25947 731 25953 765
rect 25907 693 25953 731
rect 25907 659 25913 693
rect 25947 659 25953 693
rect 25907 621 25953 659
rect 25907 587 25913 621
rect 25947 587 25953 621
rect 25907 549 25953 587
rect 25907 515 25913 549
rect 25947 515 25953 549
rect 25907 477 25953 515
rect 25907 443 25913 477
rect 25947 443 25953 477
rect 25907 405 25953 443
rect 25907 371 25913 405
rect 25947 371 25953 405
rect 25907 355 25953 371
rect 26365 1629 26411 1645
rect 26365 1595 26371 1629
rect 26405 1595 26411 1629
rect 26365 1557 26411 1595
rect 26365 1523 26371 1557
rect 26405 1523 26411 1557
rect 26365 1485 26411 1523
rect 26365 1451 26371 1485
rect 26405 1451 26411 1485
rect 26365 1413 26411 1451
rect 26365 1379 26371 1413
rect 26405 1379 26411 1413
rect 26365 1341 26411 1379
rect 26365 1307 26371 1341
rect 26405 1307 26411 1341
rect 26365 1269 26411 1307
rect 26365 1235 26371 1269
rect 26405 1235 26411 1269
rect 26365 1197 26411 1235
rect 26365 1163 26371 1197
rect 26405 1163 26411 1197
rect 26365 1125 26411 1163
rect 26365 1091 26371 1125
rect 26405 1091 26411 1125
rect 26365 1053 26411 1091
rect 26365 1019 26371 1053
rect 26405 1019 26411 1053
rect 26365 981 26411 1019
rect 26365 947 26371 981
rect 26405 947 26411 981
rect 26365 909 26411 947
rect 26365 875 26371 909
rect 26405 875 26411 909
rect 26365 837 26411 875
rect 26365 803 26371 837
rect 26405 803 26411 837
rect 26365 765 26411 803
rect 26365 731 26371 765
rect 26405 731 26411 765
rect 26365 693 26411 731
rect 26365 659 26371 693
rect 26405 659 26411 693
rect 26365 621 26411 659
rect 26365 587 26371 621
rect 26405 587 26411 621
rect 26365 549 26411 587
rect 26365 515 26371 549
rect 26405 515 26411 549
rect 26365 477 26411 515
rect 26365 443 26371 477
rect 26405 443 26411 477
rect 26365 405 26411 443
rect 26365 371 26371 405
rect 26405 371 26411 405
rect 26365 355 26411 371
rect 26823 1629 26869 1645
rect 26823 1595 26829 1629
rect 26863 1595 26869 1629
rect 26823 1557 26869 1595
rect 26823 1523 26829 1557
rect 26863 1523 26869 1557
rect 26823 1485 26869 1523
rect 26823 1451 26829 1485
rect 26863 1451 26869 1485
rect 26823 1413 26869 1451
rect 26823 1379 26829 1413
rect 26863 1379 26869 1413
rect 26823 1341 26869 1379
rect 26823 1307 26829 1341
rect 26863 1307 26869 1341
rect 26823 1269 26869 1307
rect 26823 1235 26829 1269
rect 26863 1235 26869 1269
rect 26823 1197 26869 1235
rect 26823 1163 26829 1197
rect 26863 1163 26869 1197
rect 26823 1125 26869 1163
rect 26823 1091 26829 1125
rect 26863 1091 26869 1125
rect 26823 1053 26869 1091
rect 26823 1019 26829 1053
rect 26863 1019 26869 1053
rect 26823 981 26869 1019
rect 26823 947 26829 981
rect 26863 947 26869 981
rect 26823 909 26869 947
rect 26823 875 26829 909
rect 26863 875 26869 909
rect 26823 837 26869 875
rect 26823 803 26829 837
rect 26863 803 26869 837
rect 26823 765 26869 803
rect 26823 731 26829 765
rect 26863 731 26869 765
rect 26823 693 26869 731
rect 26823 659 26829 693
rect 26863 659 26869 693
rect 26823 621 26869 659
rect 26823 587 26829 621
rect 26863 587 26869 621
rect 26823 549 26869 587
rect 26823 515 26829 549
rect 26863 515 26869 549
rect 26823 477 26869 515
rect 26823 443 26829 477
rect 26863 443 26869 477
rect 26823 405 26869 443
rect 26823 371 26829 405
rect 26863 371 26869 405
rect 26823 355 26869 371
rect 27281 1629 27327 1645
rect 27281 1595 27287 1629
rect 27321 1595 27327 1629
rect 27281 1557 27327 1595
rect 27281 1523 27287 1557
rect 27321 1523 27327 1557
rect 27281 1485 27327 1523
rect 27281 1451 27287 1485
rect 27321 1451 27327 1485
rect 27281 1413 27327 1451
rect 27281 1379 27287 1413
rect 27321 1379 27327 1413
rect 27281 1341 27327 1379
rect 27281 1307 27287 1341
rect 27321 1307 27327 1341
rect 27281 1269 27327 1307
rect 27281 1235 27287 1269
rect 27321 1235 27327 1269
rect 27281 1197 27327 1235
rect 27281 1163 27287 1197
rect 27321 1163 27327 1197
rect 27281 1125 27327 1163
rect 27281 1091 27287 1125
rect 27321 1091 27327 1125
rect 27281 1053 27327 1091
rect 27281 1019 27287 1053
rect 27321 1019 27327 1053
rect 27281 981 27327 1019
rect 27281 947 27287 981
rect 27321 947 27327 981
rect 27281 909 27327 947
rect 27281 875 27287 909
rect 27321 875 27327 909
rect 27281 837 27327 875
rect 27281 803 27287 837
rect 27321 803 27327 837
rect 27281 765 27327 803
rect 27281 731 27287 765
rect 27321 731 27327 765
rect 27281 693 27327 731
rect 27281 659 27287 693
rect 27321 659 27327 693
rect 27281 621 27327 659
rect 27281 587 27287 621
rect 27321 587 27327 621
rect 27281 549 27327 587
rect 27281 515 27287 549
rect 27321 515 27327 549
rect 27281 477 27327 515
rect 27281 443 27287 477
rect 27321 443 27327 477
rect 27281 405 27327 443
rect 27281 371 27287 405
rect 27321 371 27327 405
rect 27281 355 27327 371
rect 27739 1629 27785 1645
rect 27739 1595 27745 1629
rect 27779 1595 27785 1629
rect 27739 1557 27785 1595
rect 27739 1523 27745 1557
rect 27779 1523 27785 1557
rect 27739 1485 27785 1523
rect 27739 1451 27745 1485
rect 27779 1451 27785 1485
rect 27739 1413 27785 1451
rect 27739 1379 27745 1413
rect 27779 1379 27785 1413
rect 27739 1341 27785 1379
rect 27739 1307 27745 1341
rect 27779 1307 27785 1341
rect 27739 1269 27785 1307
rect 27739 1235 27745 1269
rect 27779 1235 27785 1269
rect 27739 1197 27785 1235
rect 27739 1163 27745 1197
rect 27779 1163 27785 1197
rect 27739 1125 27785 1163
rect 27739 1091 27745 1125
rect 27779 1091 27785 1125
rect 27739 1053 27785 1091
rect 27739 1019 27745 1053
rect 27779 1019 27785 1053
rect 27739 981 27785 1019
rect 27739 947 27745 981
rect 27779 947 27785 981
rect 27739 909 27785 947
rect 27739 875 27745 909
rect 27779 875 27785 909
rect 27739 837 27785 875
rect 27739 803 27745 837
rect 27779 803 27785 837
rect 27739 765 27785 803
rect 27739 731 27745 765
rect 27779 731 27785 765
rect 27739 693 27785 731
rect 27739 659 27745 693
rect 27779 659 27785 693
rect 27739 621 27785 659
rect 27739 587 27745 621
rect 27779 587 27785 621
rect 27739 549 27785 587
rect 27739 515 27745 549
rect 27779 515 27785 549
rect 27739 477 27785 515
rect 27739 443 27745 477
rect 27779 443 27785 477
rect 27739 405 27785 443
rect 27739 371 27745 405
rect 27779 371 27785 405
rect 27739 355 27785 371
rect 120 17 27826 60
rect 120 -17 401 17
rect 435 -17 801 17
rect 835 -17 1201 17
rect 1235 -17 1601 17
rect 1635 -17 2001 17
rect 2035 -17 2401 17
rect 2435 -17 2801 17
rect 2835 -17 3201 17
rect 3235 -17 3601 17
rect 3635 -17 4001 17
rect 4035 -17 4401 17
rect 4435 -17 4801 17
rect 4835 -17 5201 17
rect 5235 -17 5601 17
rect 5635 -17 6001 17
rect 6035 -17 6401 17
rect 6435 -17 6801 17
rect 6835 -17 7201 17
rect 7235 -17 7601 17
rect 7635 -17 8001 17
rect 8035 -17 8401 17
rect 8435 -17 8801 17
rect 8835 -17 9201 17
rect 9235 -17 9601 17
rect 9635 -17 10001 17
rect 10035 -17 10401 17
rect 10435 -17 10801 17
rect 10835 -17 11201 17
rect 11235 -17 11601 17
rect 11635 -17 12001 17
rect 12035 -17 12401 17
rect 12435 -17 12801 17
rect 12835 -17 13201 17
rect 13235 -17 13601 17
rect 13635 -17 14001 17
rect 14035 -17 14401 17
rect 14435 -17 14801 17
rect 14835 -17 15201 17
rect 15235 -17 15601 17
rect 15635 -17 16001 17
rect 16035 -17 16401 17
rect 16435 -17 16801 17
rect 16835 -17 17201 17
rect 17235 -17 17601 17
rect 17635 -17 18001 17
rect 18035 -17 18401 17
rect 18435 -17 18801 17
rect 18835 -17 19201 17
rect 19235 -17 19601 17
rect 19635 -17 20001 17
rect 20035 -17 20401 17
rect 20435 -17 20801 17
rect 20835 -17 21201 17
rect 21235 -17 21601 17
rect 21635 -17 22001 17
rect 22035 -17 22401 17
rect 22435 -17 22801 17
rect 22835 -17 23201 17
rect 23235 -17 23601 17
rect 23635 -17 24001 17
rect 24035 -17 24401 17
rect 24435 -17 24801 17
rect 24835 -17 25201 17
rect 25235 -17 25601 17
rect 25635 -17 26001 17
rect 26035 -17 26401 17
rect 26435 -17 26801 17
rect 26835 -17 27201 17
rect 27235 -17 27601 17
rect 27635 -17 27826 17
rect 120 -60 27826 -17
<< labels >>
flabel locali s 27766 104 27826 164 1 FreeSans 1250 0 0 0 GATE
port 1 nsew
flabel locali s 27766 1690 27826 1730 1 FreeSans 1250 0 0 0 SOURCE
port 2 nsew
flabel locali s 27766 210 27826 270 1 FreeSans 1250 0 0 0 DRAIN
port 3 nsew
flabel nwell s 120 1850 180 1910 1 FreeSans 1250 0 0 0 VPWR
port 4 nsew
flabel metal1 s 120 -30 278 30 1 FreeSans 1250 0 0 0 VGND
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 27947 1880
<< end >>
