magic
tech sky130A
timestamp 1655323538
<< metal4 >>
rect -500 459 500 500
rect -500 -459 -459 459
rect 459 -459 500 459
rect -500 -500 500 -459
<< via4 >>
rect -459 -459 459 459
<< metal5 >>
rect -500 459 500 500
rect -500 -459 -459 459
rect 459 -459 500 459
rect -500 -500 500 -459
<< end >>
