magic
tech sky130A
timestamp 1656729169
<< metal4 >>
rect -90 379 90 406
rect -90 261 -59 379
rect 59 261 90 379
rect -90 219 90 261
rect -90 101 -59 219
rect 59 101 90 219
rect -90 59 90 101
rect -90 -59 -59 59
rect 59 -59 90 59
rect -90 -101 90 -59
rect -90 -219 -59 -101
rect 59 -219 90 -101
rect -90 -261 90 -219
rect -90 -379 -59 -261
rect 59 -379 90 -261
rect -90 -406 90 -379
<< via4 >>
rect -59 261 59 379
rect -59 101 59 219
rect -59 -59 59 59
rect -59 -219 59 -101
rect -59 -379 59 -261
<< metal5 >>
rect -90 379 90 406
rect -90 261 -59 379
rect 59 261 90 379
rect -90 219 90 261
rect -90 101 -59 219
rect 59 101 90 219
rect -90 59 90 101
rect -90 -59 -59 59
rect 59 -59 90 59
rect -90 -101 90 -59
rect -90 -219 -59 -101
rect 59 -219 90 -101
rect -90 -261 90 -219
rect -90 -379 -59 -261
rect 59 -379 90 -261
rect -90 -406 90 -379
<< properties >>
string GDS_END 9314460
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/merge/design_merged.gds
string GDS_START 9314008
<< end >>
