magic
tech sky130A
timestamp 1655323538
<< metal4 >>
rect -196 459 196 500
rect -196 -459 -139 459
rect 139 -459 196 459
rect -196 -500 196 -459
<< via4 >>
rect -139 -459 139 459
<< metal5 >>
rect -196 459 196 500
rect -196 -459 -139 459
rect 139 -459 196 459
rect -196 -500 196 -459
<< end >>
