magic
tech sky130A
magscale 1 2
timestamp 1656729169
<< error_p >>
rect -403 142 403 178
<< metal4 >>
rect -403 118 403 142
rect -403 -118 -278 118
rect -42 -118 403 118
rect -403 -142 403 -118
<< via4 >>
rect -278 -118 -42 118
<< metal5 >>
rect -403 118 403 142
rect -403 -118 -278 118
rect -42 -118 403 118
rect -403 -142 403 -118
<< properties >>
string GDS_END 9322338
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/merge/design_merged.gds
string GDS_START 9322142
<< end >>
