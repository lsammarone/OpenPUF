magic
tech sky130A
timestamp 1655322987
<< metal2 >>
rect -90 74 90 90
rect -90 -74 -74 74
rect 74 -74 90 74
rect -90 -90 90 -74
<< via2 >>
rect -74 -74 74 74
<< metal3 >>
rect -90 74 90 90
rect -90 -74 -74 74
rect 74 -74 90 74
rect -90 -90 90 -74
<< end >>
