magic
tech sky130A
timestamp 1656729169
<< metal4 >>
rect -90 139 90 226
rect -90 21 -59 139
rect 59 21 90 139
rect -90 -21 90 21
rect -90 -139 -59 -21
rect 59 -139 90 -21
rect -90 -226 90 -139
<< via4 >>
rect -59 21 59 139
rect -59 -139 59 -21
<< metal5 >>
rect -90 139 90 226
rect -90 21 -59 139
rect 59 21 90 139
rect -90 -21 90 21
rect -90 -139 -59 -21
rect 59 -139 90 -21
rect -90 -226 90 -139
<< properties >>
string GDS_END 9361570
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/merge/design_merged.gds
string GDS_START 9361310
<< end >>
