magic
tech sky130A
magscale 1 2
timestamp 1483428465
<< checkpaint >>
rect -1440 -1637 1440 1637
<< metal4 >>
rect -180 278 180 377
rect -180 42 -118 278
rect 118 42 180 278
rect -180 -42 180 42
rect -180 -278 -118 -42
rect 118 -278 180 -42
rect -180 -377 180 -278
<< via4 >>
rect -118 42 118 278
rect -118 -278 118 -42
<< metal5 >>
rect -180 278 180 377
rect -180 42 -118 278
rect 118 42 180 278
rect -180 -42 180 42
rect -180 -278 -118 -42
rect 118 -278 180 -42
rect -180 -377 180 -278
<< end >>
