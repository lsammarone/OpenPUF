magic
tech sky130A
timestamp 1483428465
<< checkpaint >>
rect -826 -701 826 701
<< metal4 >>
rect -196 59 196 71
rect -196 -59 -139 59
rect -21 -59 21 59
rect 139 -59 196 59
rect -196 -71 196 -59
<< via4 >>
rect -139 -59 -21 59
rect 21 -59 139 59
<< metal5 >>
rect -196 59 196 71
rect -196 -59 -139 59
rect -21 -59 21 59
rect 139 -59 196 59
rect -196 -71 196 -59
<< end >>
