* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_1 Y A VGND VPWR VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_1 Y B A VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VNB VPB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 X A VGND VPWR VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_8 Y A VGND VPWR VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 Q RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_1 B Y A VGND VPWR VNB VPB a_109_297#
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 X A VGND VPWR VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_16 Y A VGND VPWR VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_4 Y A VPWR VGND VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_1#0 a_150_47# w_n38_261# a_68_47# a_68_297# a_64_199#
+ VSUBS
X0 a_150_47# a_64_199# a_68_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_150_47# a_64_199# a_68_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_hvt_UUWA33 a_n73_n100# a_15_n100# w_n109_n200# a_n33_n197#
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n109_n200# sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_hvt_SH6FHF w_n161_n200# a_n125_n100# a_63_n100# a_15_131#
+ a_n33_n100# a_n81_n197#
X0 a_63_n100# a_15_131# a_n33_n100# w_n161_n200# sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n33_n100# a_n81_n197# a_n125_n100# w_n161_n200# sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_PX9ZJG a_63_n65# a_n125_n65# a_15_87# a_n81_n153#
+ a_n33_n65# VSUBS
X0 a_n33_n65# a_n81_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_63_n65# a_15_87# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt mux 2/VSUBS w_n54_614# m1_188_418# m1_76_558# a_28_318# m1_n50_88# m1_46_n2#
Xsky130_fd_pr__pfet_01v8_hvt_SH6FHF_4 w_n54_614# m1_n50_88# m1_188_418# m1_46_n2#
+ m1_76_558# a_28_318# sky130_fd_pr__pfet_01v8_hvt_SH6FHF
X1 m1_188_418# m1_n50_88# a_28_318# m1_46_n2# m1_76_558# 2/VSUBS sky130_fd_pr__nfet_01v8_PX9ZJG
X2 w_n54_614# m1_n50_88# m1_188_418# m1_46_n2# m1_76_558# a_28_318# sky130_fd_pr__pfet_01v8_hvt_SH6FHF
Xsky130_fd_pr__nfet_01v8_PX9ZJG_0 m1_188_418# m1_n50_88# a_28_318# m1_46_n2# m1_76_558#
+ 2/VSUBS sky130_fd_pr__nfet_01v8_PX9ZJG
Xsky130_fd_pr__nfet_01v8_PX9ZJG_1 m1_188_418# m1_n50_88# a_28_318# m1_46_n2# m1_76_558#
+ 2/VSUBS sky130_fd_pr__nfet_01v8_PX9ZJG
Xsky130_fd_pr__nfet_01v8_PX9ZJG_2 m1_188_418# m1_n50_88# a_28_318# m1_46_n2# m1_76_558#
+ 2/VSUBS sky130_fd_pr__nfet_01v8_PX9ZJG
Xsky130_fd_pr__nfet_01v8_PX9ZJG_4 m1_188_418# m1_n50_88# a_28_318# m1_46_n2# m1_76_558#
+ 2/VSUBS sky130_fd_pr__nfet_01v8_PX9ZJG
Xsky130_fd_pr__nfet_01v8_PX9ZJG_3 m1_188_418# m1_n50_88# a_28_318# m1_46_n2# m1_76_558#
+ 2/VSUBS sky130_fd_pr__nfet_01v8_PX9ZJG
Xsky130_fd_pr__pfet_01v8_hvt_SH6FHF_0 w_n54_614# m1_n50_88# m1_188_418# m1_46_n2#
+ m1_76_558# a_28_318# sky130_fd_pr__pfet_01v8_hvt_SH6FHF
Xsky130_fd_pr__pfet_01v8_hvt_SH6FHF_1 w_n54_614# m1_n50_88# m1_188_418# m1_46_n2#
+ m1_76_558# a_28_318# sky130_fd_pr__pfet_01v8_hvt_SH6FHF
Xsky130_fd_pr__pfet_01v8_hvt_SH6FHF_2 w_n54_614# m1_n50_88# m1_188_418# m1_46_n2#
+ m1_76_558# a_28_318# sky130_fd_pr__pfet_01v8_hvt_SH6FHF
Xsky130_fd_pr__pfet_01v8_hvt_SH6FHF_3 w_n54_614# m1_n50_88# m1_188_418# m1_46_n2#
+ m1_76_558# a_28_318# sky130_fd_pr__pfet_01v8_hvt_SH6FHF
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VNB VPB a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt demux m1_188_418# 2/VSUBS w_n54_614# m1_46_n2# m1_76_558# a_28_318# m1_n50_88#
X1 m1_188_418# m1_n50_88# a_28_318# m1_46_n2# m1_76_558# 2/VSUBS sky130_fd_pr__nfet_01v8_PX9ZJG
X2 w_n54_614# m1_n50_88# m1_188_418# m1_46_n2# m1_76_558# a_28_318# sky130_fd_pr__pfet_01v8_hvt_SH6FHF
Xsky130_fd_pr__nfet_01v8_PX9ZJG_0 m1_188_418# m1_n50_88# a_28_318# m1_46_n2# m1_76_558#
+ 2/VSUBS sky130_fd_pr__nfet_01v8_PX9ZJG
Xsky130_fd_pr__nfet_01v8_PX9ZJG_1 m1_188_418# m1_n50_88# a_28_318# m1_46_n2# m1_76_558#
+ 2/VSUBS sky130_fd_pr__nfet_01v8_PX9ZJG
Xsky130_fd_pr__pfet_01v8_hvt_SH6FHF_0 w_n54_614# m1_n50_88# m1_188_418# m1_46_n2#
+ m1_76_558# a_28_318# sky130_fd_pr__pfet_01v8_hvt_SH6FHF
Xsky130_fd_pr__pfet_01v8_hvt_SH6FHF_1 w_n54_614# m1_n50_88# m1_188_418# m1_46_n2#
+ m1_76_558# a_28_318# sky130_fd_pr__pfet_01v8_hvt_SH6FHF
.ends

.subckt unitcell2buf sky130_fd_sc_hd__nor2_1_3/a_109_297# sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ sky130_fd_sc_hd__buf_1_1/X li_n460_n386# sky130_fd_sc_hd__buf_1_1/a_27_47# sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nor2_1_2/Y li_80_172# m2_136_462# sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__nor2_1_3/A a_24_n198# sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__buf_1_1/A VSUBS
Xsky130_fd_sc_hd__inv_1#0_0 li_80_172# sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ a_24_n198# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1#0_1 a_24_n198# sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ li_n460_n386# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__nor2_1_3/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__nor2_1_3/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__nor2_1_2/Y
+ sky130_fd_sc_hd__nor2_1_3/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__nor2_1_2/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_2 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__nor2_1_2/Y
+ sky130_fd_sc_hd__nor2_1_3/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__nor2_1_2/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_3 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__nor2_1_3/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__nor2_1_3/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_pr__pfet_01v8_hvt_UUWA33_0 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__buf_1_1/VPB li_80_172# sky130_fd_pr__pfet_01v8_hvt_UUWA33
X1 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/VPB
+ li_80_172# sky130_fd_pr__pfet_01v8_hvt_UUWA33
Xsky130_fd_pr__pfet_01v8_hvt_UUWA33_1 sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__buf_1_1/VPB a_24_n198# sky130_fd_pr__pfet_01v8_hvt_UUWA33
X2 sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__buf_1_1/VPB
+ a_24_n198# sky130_fd_pr__pfet_01v8_hvt_UUWA33
Xmux_0 VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__buf_1_1/A
+ a_24_n198# sky130_fd_sc_hd__nor2_1_2/Y li_80_172# mux
Xmux_1 VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__buf_1_1/A
+ a_24_n198# sky130_fd_sc_hd__nor2_1_2/Y li_80_172# mux
Xsky130_fd_sc_hd__buf_1_0 VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/X
+ sky130_fd_sc_hd__buf_1_1/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__buf_1_1 VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/X
+ sky130_fd_sc_hd__buf_1_1/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__inv_1_0 li_80_172# sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ a_24_n198# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1_1 a_24_n198# sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ li_n460_n386# VSUBS sky130_fd_sc_hd__inv_1#0
Xdemux_0 sky130_fd_sc_hd__nor2_1_3/B VSUBS sky130_fd_sc_hd__buf_1_1/VPB li_80_172#
+ m2_136_462# a_24_n198# sky130_fd_sc_hd__nor2_1_2/B demux
Xdemux_1 sky130_fd_sc_hd__nor2_1_3/B VSUBS sky130_fd_sc_hd__buf_1_1/VPB li_80_172#
+ m2_136_462# a_24_n198# sky130_fd_sc_hd__nor2_1_2/B demux
.ends

.subckt unitcell2bufcut sky130_fd_sc_hd__nor2_1_3/a_109_297# sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ sky130_fd_sc_hd__nor2_1_2/B a_24_n198# li_n460_n386# sky130_fd_sc_hd__buf_1_1/a_27_47#
+ sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__nor2_1_2/Y m2_136_462# li_80_172# sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__buf_1_1/X sky130_fd_sc_hd__nor2_1_3/A sky130_fd_sc_hd__nor2_1_3/B
+ VSUBS sky130_fd_sc_hd__buf_1_1/A
Xsky130_fd_sc_hd__inv_1#0_0 li_80_172# sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ a_24_n198# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1#0_1 a_24_n198# sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ li_n460_n386# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__nor2_1_3/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__nor2_1_3/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__nor2_1_2/Y
+ sky130_fd_sc_hd__nor2_1_3/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__nor2_1_2/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_2 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__nor2_1_2/Y
+ sky130_fd_sc_hd__nor2_1_3/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__nor2_1_2/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_3 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__nor2_1_3/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__nor2_1_3/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_pr__pfet_01v8_hvt_UUWA33_0 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__buf_1_1/VPB li_80_172# sky130_fd_pr__pfet_01v8_hvt_UUWA33
X1 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/VPB
+ li_80_172# sky130_fd_pr__pfet_01v8_hvt_UUWA33
Xsky130_fd_pr__pfet_01v8_hvt_UUWA33_1 sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__buf_1_1/VPB a_24_n198# sky130_fd_pr__pfet_01v8_hvt_UUWA33
X2 sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__buf_1_1/VPB
+ a_24_n198# sky130_fd_pr__pfet_01v8_hvt_UUWA33
Xmux_0 VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__buf_1_1/A
+ a_24_n198# sky130_fd_sc_hd__nor2_1_2/Y li_80_172# mux
Xmux_1 VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__buf_1_1/A
+ a_24_n198# sky130_fd_sc_hd__nor2_1_2/Y li_80_172# mux
Xsky130_fd_sc_hd__buf_1_0 VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/X
+ sky130_fd_sc_hd__buf_1_1/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__buf_1_1 VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/X
+ sky130_fd_sc_hd__buf_1_1/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__inv_1_0 li_80_172# sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ a_24_n198# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1_1 a_24_n198# sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ li_n460_n386# VSUBS sky130_fd_sc_hd__inv_1#0
Xdemux_0 sky130_fd_sc_hd__nor2_1_3/B VSUBS sky130_fd_sc_hd__buf_1_1/VPB li_80_172#
+ m2_136_462# a_24_n198# sky130_fd_sc_hd__nor2_1_2/B demux
Xdemux_1 sky130_fd_sc_hd__nor2_1_3/B VSUBS sky130_fd_sc_hd__buf_1_1/VPB li_80_172#
+ m2_136_462# a_24_n198# sky130_fd_sc_hd__nor2_1_2/B demux
.ends

.subckt brbufhalf unitcell2buf_7/li_n460_n386# unitcell2bufcut_3/li_n460_n386# sky130_fd_sc_hd__inv_16_7/A
+ unitcell2buf_2/li_n460_n386# unitcell2buf_24/li_n460_n386# sky130_fd_sc_hd__inv_16_6/VGND
+ unitcell2buf_5/li_n460_n386# unitcell2buf_27/li_n460_n386# unitcell2buf_8/li_n460_n386#
+ unitcell2buf_0/li_n460_n386# unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_7/VGND unitcell2buf_25/li_n460_n386# unitcell2bufcut_2/li_n460_n386#
+ unitcell2buf_6/li_n460_n386# sky130_fd_sc_hd__inv_16_4/VGND unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_9/li_n460_n386# unitcell2buf_1/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_5/A
+ unitcell2buf_26/m2_136_462# sky130_fd_sc_hd__inv_16_5/VGND VSUBS unitcell2buf_26/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_7/VPB
Xunitcell2buf_1 unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_1/li_n460_n386# unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_1/li_80_172# unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_1/a_24_n198#
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/A
+ sky130_fd_sc_hd__inv_16_7/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_2 unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_2/li_n460_n386# unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_2/li_80_172# unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_2/a_24_n198#
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_4 sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_5/A
+ sky130_fd_sc_hd__inv_16_4/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_5 sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_5/A
+ sky130_fd_sc_hd__inv_16_5/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_3 unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_3/li_n460_n386# unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_3/li_80_172# unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_3/a_24_n198#
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_6 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/A
+ sky130_fd_sc_hd__inv_16_6/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_4 unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_4/li_n460_n386# unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_4/li_80_172# unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_4/a_24_n198#
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_7 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/A
+ sky130_fd_sc_hd__inv_16_7/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_5 unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_5/li_n460_n386# unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_5/li_80_172# unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_5/a_24_n198#
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_6 unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_6/li_n460_n386# unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_6/li_80_172# unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_6/a_24_n198#
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_7 unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_7/li_n460_n386# unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_7/li_80_172# unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_7/a_24_n198#
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_8 unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_8/li_n460_n386# unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_8/li_80_172# unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_8/a_24_n198#
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_9 unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_9/li_n460_n386# unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_9/li_80_172# unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_9/a_24_n198#
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_20 unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_6/li_n460_n386# unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_6/li_80_172# unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_6/a_24_n198#
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_21 unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_7/li_n460_n386# unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_7/li_80_172# unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_7/a_24_n198#
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_22 unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_8/li_n460_n386# unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_8/li_80_172# unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_8/a_24_n198#
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_10 unitcell2buf_24/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_24/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_24/li_n460_n386# unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_24/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_24/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_24/li_80_172# unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_24/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_24/a_24_n198#
+ unitcell2buf_24/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_11 unitcell2buf_25/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_25/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_25/li_n460_n386# unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_25/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_25/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_25/li_80_172# unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_25/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_25/a_24_n198#
+ unitcell2buf_25/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_23 unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_9/li_n460_n386# unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_9/li_80_172# unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_9/a_24_n198#
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_12 unitcell2buf_26/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_26/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_26/li_n460_n386# unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_26/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_26/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_26/li_80_172# unitcell2buf_26/m2_136_462# sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_26/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_26/a_24_n198#
+ unitcell2buf_26/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_24 unitcell2buf_24/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_24/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_24/li_n460_n386# unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_24/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_24/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_24/li_80_172# unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_24/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_24/a_24_n198#
+ unitcell2buf_24/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_13 unitcell2buf_27/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_27/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_27/li_n460_n386# unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_27/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_27/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_27/li_80_172# unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_27/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_27/a_24_n198#
+ unitcell2buf_27/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_14 unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_0/li_n460_n386# unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_0/li_80_172# unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_0/a_24_n198#
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_25 unitcell2buf_25/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_25/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_25/li_n460_n386# unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_25/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_25/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_25/li_80_172# unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_25/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_25/a_24_n198#
+ unitcell2buf_25/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_15 unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_1/li_n460_n386# unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_1/li_80_172# unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_1/a_24_n198#
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_26 unitcell2buf_26/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_26/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_26/li_n460_n386# unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_26/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_26/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_26/li_80_172# unitcell2buf_26/m2_136_462# sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_26/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_26/a_24_n198#
+ unitcell2buf_26/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_16 unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_2/li_n460_n386# unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_2/li_80_172# unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_2/a_24_n198#
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_27 unitcell2buf_27/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_27/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_27/li_n460_n386# unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_27/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_27/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_27/li_80_172# unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_27/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_27/a_24_n198#
+ unitcell2buf_27/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_17 unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_3/li_n460_n386# unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_3/li_80_172# unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_3/a_24_n198#
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_18 unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_4/li_n460_n386# unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_4/li_80_172# unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_4/a_24_n198#
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_19 unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_5/li_n460_n386# unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_5/li_80_172# unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_5/a_24_n198#
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2bufcut_0 unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_2/B unitcell2bufcut_2/a_24_n198# unitcell2bufcut_2/li_n460_n386#
+ unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2bufcut_2/li_80_172# sky130_fd_sc_hd__inv_16_7/VPB unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_3/B VSUBS
+ unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_5/A
+ sky130_fd_sc_hd__inv_16_4/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2bufcut_1 unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_2/B unitcell2bufcut_3/a_24_n198# unitcell2bufcut_3/li_n460_n386#
+ unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2bufcut_3/li_80_172# sky130_fd_sc_hd__inv_16_7/VPB unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/X
+ sky130_fd_sc_hd__inv_16_7/Y unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_3/B VSUBS
+ unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut
Xunitcell2bufcut_2 unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_2/B unitcell2bufcut_2/a_24_n198# unitcell2bufcut_2/li_n460_n386#
+ unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2bufcut_2/li_80_172# sky130_fd_sc_hd__inv_16_7/VPB unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_3/B VSUBS
+ unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_5/A
+ sky130_fd_sc_hd__inv_16_5/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_0 unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_0/li_n460_n386# unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_0/li_80_172# unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_0/a_24_n198#
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2bufcut_3 unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_2/B unitcell2bufcut_3/a_24_n198# unitcell2bufcut_3/li_n460_n386#
+ unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2bufcut_3/li_80_172# sky130_fd_sc_hd__inv_16_7/VPB unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/X
+ sky130_fd_sc_hd__inv_16_7/Y unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_3/B VSUBS
+ unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/A
+ sky130_fd_sc_hd__inv_16_6/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
.ends

.subckt brbufhalf_64 unitcell2buf_7/li_n460_n386# unitcell2buf_2/li_n460_n386# unitcell2buf_10/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_2/VGND unitcell2buf_5/li_n460_n386# unitcell2buf_13/li_n460_n386#
+ unitcell2buf_8/li_n460_n386# sky130_fd_sc_hd__inv_16_1/A unitcell2buf_0/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/A unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/VGND unitcell2buf_11/li_n460_n386# sky130_fd_sc_hd__inv_16_0/VGND
+ unitcell2bufcut_0/li_n460_n386# unitcell2buf_6/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_9/li_n460_n386# unitcell2buf_1/li_n460_n386# unitcell2buf_4/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_1/VGND unitcell2buf_12/m2_136_462# VSUBS unitcell2buf_12/li_n460_n386#
Xunitcell2buf_1 unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_1/li_n460_n386# unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_1/li_80_172# unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_1/a_24_n198#
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16_3/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_2 unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_2/li_n460_n386# unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_2/li_80_172# unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_2/a_24_n198#
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_3 unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_3/li_n460_n386# unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_3/li_80_172# unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_3/a_24_n198#
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_4 unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_4/li_n460_n386# unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_4/li_80_172# unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_4/a_24_n198#
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_5 unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_5/li_n460_n386# unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_5/li_80_172# unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_5/a_24_n198#
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_6 unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_6/li_n460_n386# unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_6/li_80_172# unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_6/a_24_n198#
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_7 unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_7/li_n460_n386# unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_7/li_80_172# unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_7/a_24_n198#
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_8 unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_8/li_n460_n386# unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_8/li_80_172# unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_8/a_24_n198#
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_9 unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_9/li_n460_n386# unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_9/li_80_172# unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_9/a_24_n198#
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_10 unitcell2buf_10/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_10/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_10/li_n460_n386# unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_10/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_10/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_10/li_80_172# unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_10/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_10/a_24_n198#
+ unitcell2buf_10/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_11 unitcell2buf_11/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_11/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_11/li_n460_n386# unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_11/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_11/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_11/li_80_172# unitcell2buf_13/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_11/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_11/a_24_n198#
+ unitcell2buf_11/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_12 unitcell2buf_12/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_12/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_12/li_n460_n386# unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_12/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_12/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_12/li_80_172# unitcell2buf_12/m2_136_462# sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_12/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_12/a_24_n198#
+ unitcell2buf_12/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_13 unitcell2buf_13/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_13/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_13/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_13/li_n460_n386# unitcell2buf_13/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_13/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_13/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_13/li_80_172# unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_13/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_13/a_24_n198#
+ unitcell2buf_13/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_13/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2bufcut_0 unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_2/B unitcell2bufcut_0/a_24_n198# unitcell2bufcut_0/li_n460_n386#
+ unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2bufcut_0/li_80_172# sky130_fd_sc_hd__inv_16_3/VPB unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/X
+ sky130_fd_sc_hd__inv_16_3/Y unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_3/B VSUBS
+ unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_0/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_1/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_0 unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_0/li_n460_n386# unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_0/li_80_172# unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_0/a_24_n198#
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16_2/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
.ends

.subckt BR64 OUT VDD RESET C[0] C[1] C[2] C[3] C[4] C[5] C[6] C[7] C[8] C[9] C[10]
+ C[11] C[12] C[13] C[14] C[15] C[16] C[17] C[18] C[19] C[20] C[21] C[22] C[23] C[24]
+ C[25] C[26] C[27] C[28] C[29] C[30] C[31] C[32] C[33] C[34] C[35] C[36] C[37] C[38]
+ C[39] C[40] C[41] C[42] C[43] C[44] C[45] C[46] C[47] C[48] C[49] C[50] C[51] C[52]
+ C[53] C[54] C[55] C[56] C[57] C[58] C[59] C[60] C[61] C[62] C[63] VSS
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__inv_16_4/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_4 sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__inv_16_4/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_4_0 sky130_fd_sc_hd__inv_4_0/Y RESET VDD VSS VSS VDD sky130_fd_sc_hd__inv_4
Xbrbufhalf_0 C[6] C[7] sky130_fd_sc_hd__inv_16_1/Y C[12] C[3] VSS C[9] C[1] C[5] C[14]
+ brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X C[11] VSS C[2] C[15] C[8]
+ VSS brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A brbufhalf_0/sky130_fd_sc_hd__inv_16_7/Y
+ C[4] C[13] brbufhalf_0/sky130_fd_sc_hd__inv_16_5/Y C[10] sky130_fd_sc_hd__inv_16_1/Y
+ brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A VSS VSS C[0] VDD brbufhalf
Xbrbufhalf_1 C[54] C[55] sky130_fd_sc_hd__inv_16_1/Y C[60] C[51] VSS C[57] C[49] C[53]
+ C[62] OUT C[59] VSS C[50] C[63] C[56] VSS brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_1/sky130_fd_sc_hd__inv_16_7/Y C[52] C[61] brbufhalf_1/sky130_fd_sc_hd__inv_16_5/Y
+ C[58] sky130_fd_sc_hd__inv_16_1/Y brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ VSS VSS C[48] VDD brbufhalf
Xbrbufhalf_2 C[38] C[39] sky130_fd_sc_hd__inv_16_4/Y C[44] C[35] VSS C[41] C[33] C[37]
+ C[46] brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X C[43] VSS C[34] C[47]
+ C[40] VSS brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A brbufhalf_2/sky130_fd_sc_hd__inv_16_7/Y
+ C[36] C[45] brbufhalf_2/sky130_fd_sc_hd__inv_16_5/Y C[42] sky130_fd_sc_hd__inv_16_4/Y
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A VSS VSS C[32] VDD brbufhalf
Xbrbufhalf_64_0 C[22] C[28] C[19] VSS C[25] C[17] C[21] sky130_fd_sc_hd__inv_16_4/Y
+ C[30] sky130_fd_sc_hd__inv_16_4/Y brbufhalf_64_0/unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ C[27] VSS C[18] VSS C[23] C[24] VDD C[20] C[29] C[26] VSS brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ VSS C[16] brbufhalf_64
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_4/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_4/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_4_0/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xunitcell2buf_0 unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/X C[31] unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_0/li_80_172# brbufhalf_64_0/unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ VDD unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/Y brbufhalf_2/sky130_fd_sc_hd__inv_16_7/Y
+ unitcell2buf_0/a_24_n198# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ VSS unitcell2buf
.ends

.subckt sky130_fd_sc_hd__nand2_2 Y A B VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt unitcell2bufcut_32 IN C VDD OUT buf_out sky130_fd_sc_hd__nor2_1_1/A VSS
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_1_0/B sky130_fd_sc_hd__nor2_1_0/Y
+ sky130_fd_sc_hd__nor2_1_1/A VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1_0/a_109_297#
+ sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_1/B sky130_fd_sc_hd__nor2_1_1/Y
+ sky130_fd_sc_hd__nor2_1_1/A VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1_1/a_109_297#
+ sky130_fd_sc_hd__nor2_1
X1 sky130_fd_sc_hd__nor2_1_0/B VDD VDD li_80_172# sky130_fd_pr__pfet_01v8_hvt_UUWA33
X2 VDD sky130_fd_sc_hd__nor2_1_1/B VDD a_24_n198# sky130_fd_pr__pfet_01v8_hvt_UUWA33
Xmux_0 VSS VDD sky130_fd_sc_hd__nor2_1_1/Y OUT a_24_n198# sky130_fd_sc_hd__nor2_1_0/Y
+ li_80_172# mux
Xsky130_fd_sc_hd__buf_1_0 VSS VDD buf_out OUT VSS VDD sky130_fd_sc_hd__buf_1_0/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__inv_1_0 li_80_172# VDD VSS VDD a_24_n198# VSS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1_1 a_24_n198# VDD VSS VDD C VSS sky130_fd_sc_hd__inv_1#0
Xdemux_0 sky130_fd_sc_hd__nor2_1_1/B VSS VDD li_80_172# IN a_24_n198# sky130_fd_sc_hd__nor2_1_0/B
+ demux
.ends

.subckt unitcell2buf_32 IN C OUT buf_out VDD RESET VSS
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_1_0/B sky130_fd_sc_hd__nor2_1_0/Y
+ RESET VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_1/B sky130_fd_sc_hd__nor2_1_1/Y
+ RESET VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1_1/a_109_297# sky130_fd_sc_hd__nor2_1
X1 sky130_fd_sc_hd__nor2_1_0/B VDD VDD li_80_172# sky130_fd_pr__pfet_01v8_hvt_UUWA33
X2 VDD sky130_fd_sc_hd__nor2_1_1/B VDD a_24_n198# sky130_fd_pr__pfet_01v8_hvt_UUWA33
Xmux_0 VSS VDD sky130_fd_sc_hd__nor2_1_1/Y OUT a_24_n198# sky130_fd_sc_hd__nor2_1_0/Y
+ li_80_172# mux
Xsky130_fd_sc_hd__buf_1_0 VSS VDD buf_out OUT VSS VDD sky130_fd_sc_hd__buf_1_0/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__inv_1_0 li_80_172# VDD VSS VDD a_24_n198# VSS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1_1 a_24_n198# VDD VSS VDD C VSS sky130_fd_sc_hd__inv_1#0
Xdemux_0 sky130_fd_sc_hd__nor2_1_1/B VSS VDD li_80_172# IN a_24_n198# sky130_fd_sc_hd__nor2_1_0/B
+ demux
.ends

.subckt brbufhalf_32 unitcell2buf_32_9/C unitcell2buf_32_0/C unitcell2bufcut_32_0/buf_out
+ unitcell2buf_32_10/C unitcell2buf_32_2/C unitcell2buf_32_12/C unitcell2buf_32_4/C
+ unitcell2bufcut_32_1/C unitcell2buf_32_6/C unitcell2buf_32_8/C sky130_fd_sc_hd__inv_16_3/A
+ unitcell2buf_32_1/C unitcell2buf_32_11/C sky130_fd_sc_hd__inv_16_3/VGND unitcell2buf_32_3/C
+ unitcell2bufcut_32_0/C unitcell2buf_32_5/C unitcell2buf_32_11/IN unitcell2bufcut_32_0/OUT
+ unitcell2buf_32_7/C sky130_fd_sc_hd__inv_16_1/A unitcell2buf_32_9/RESET sky130_fd_sc_hd__inv_16_1/VGND
+ unitcell2buf_32_9/VDD VSUBS
Xsky130_fd_sc_hd__inv_16_3 unitcell2buf_32_9/RESET sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__inv_16_3/VGND
+ unitcell2buf_32_9/VDD VSUBS unitcell2buf_32_9/VDD sky130_fd_sc_hd__inv_16
Xunitcell2bufcut_32_0 unitcell2buf_32_0/OUT unitcell2bufcut_32_0/C unitcell2buf_32_9/VDD
+ unitcell2bufcut_32_0/OUT unitcell2bufcut_32_0/buf_out unitcell2buf_32_6/RESET VSUBS
+ unitcell2bufcut_32
Xunitcell2buf_32_0 unitcell2buf_32_0/IN unitcell2buf_32_0/C unitcell2buf_32_0/OUT
+ unitcell2buf_32_0/buf_out unitcell2buf_32_9/VDD unitcell2buf_32_6/RESET VSUBS unitcell2buf_32
Xunitcell2buf_32_1 unitcell2buf_32_1/IN unitcell2buf_32_1/C unitcell2buf_32_0/IN unitcell2buf_32_1/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_6/RESET VSUBS unitcell2buf_32
Xunitcell2bufcut_32_1 unitcell2buf_32_7/OUT unitcell2bufcut_32_1/C unitcell2buf_32_9/VDD
+ unitcell2buf_32_6/IN unitcell2bufcut_32_1/buf_out unitcell2buf_32_9/RESET VSUBS
+ unitcell2bufcut_32
Xunitcell2buf_32_10 unitcell2buf_32_10/IN unitcell2buf_32_10/C unitcell2buf_32_9/IN
+ unitcell2buf_32_10/buf_out unitcell2buf_32_9/VDD unitcell2buf_32_9/RESET VSUBS unitcell2buf_32
Xunitcell2buf_32_2 unitcell2buf_32_2/IN unitcell2buf_32_2/C unitcell2buf_32_1/IN unitcell2buf_32_2/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_6/RESET VSUBS unitcell2buf_32
Xunitcell2buf_32_12 unitcell2buf_32_12/IN unitcell2buf_32_12/C unitcell2buf_32_10/IN
+ unitcell2buf_32_12/buf_out unitcell2buf_32_9/VDD unitcell2buf_32_9/RESET VSUBS unitcell2buf_32
Xunitcell2buf_32_11 unitcell2buf_32_11/IN unitcell2buf_32_11/C unitcell2buf_32_12/IN
+ unitcell2buf_32_11/buf_out unitcell2buf_32_9/VDD unitcell2buf_32_9/RESET VSUBS unitcell2buf_32
Xunitcell2buf_32_3 unitcell2buf_32_3/IN unitcell2buf_32_3/C unitcell2buf_32_2/IN unitcell2buf_32_3/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_6/RESET VSUBS unitcell2buf_32
Xunitcell2buf_32_4 unitcell2buf_32_4/IN unitcell2buf_32_4/C unitcell2buf_32_3/IN unitcell2buf_32_4/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_6/RESET VSUBS unitcell2buf_32
Xunitcell2buf_32_5 unitcell2buf_32_5/IN unitcell2buf_32_5/C unitcell2buf_32_4/IN unitcell2buf_32_5/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_6/RESET VSUBS unitcell2buf_32
Xunitcell2buf_32_6 unitcell2buf_32_6/IN unitcell2buf_32_6/C unitcell2buf_32_5/IN unitcell2buf_32_6/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_6/RESET VSUBS unitcell2buf_32
Xunitcell2buf_32_7 unitcell2buf_32_7/IN unitcell2buf_32_7/C unitcell2buf_32_7/OUT
+ unitcell2buf_32_7/buf_out unitcell2buf_32_9/VDD unitcell2buf_32_9/RESET VSUBS unitcell2buf_32
Xunitcell2buf_32_8 unitcell2buf_32_8/IN unitcell2buf_32_8/C unitcell2buf_32_7/IN unitcell2buf_32_8/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_9/RESET VSUBS unitcell2buf_32
Xunitcell2buf_32_9 unitcell2buf_32_9/IN unitcell2buf_32_9/C unitcell2buf_32_8/IN unitcell2buf_32_9/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_9/RESET VSUBS unitcell2buf_32
Xsky130_fd_sc_hd__inv_16_0 unitcell2buf_32_6/RESET sky130_fd_sc_hd__inv_16_1/A sky130_fd_sc_hd__inv_16_1/VGND
+ unitcell2buf_32_9/VDD VSUBS unitcell2buf_32_9/VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 unitcell2buf_32_6/RESET sky130_fd_sc_hd__inv_16_1/A sky130_fd_sc_hd__inv_16_1/VGND
+ unitcell2buf_32_9/VDD VSUBS unitcell2buf_32_9/VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 unitcell2buf_32_9/RESET sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__inv_16_3/VGND
+ unitcell2buf_32_9/VDD VSUBS unitcell2buf_32_9/VDD sky130_fd_sc_hd__inv_16
.ends

.subckt sky130_fd_sc_hd__inv_8 A Y VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_2 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt invcell sky130_fd_sc_hd__inv_8_1/VGND sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_8_1/VPB
+ sky130_fd_sc_hd__inv_8_1/VPWR sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__inv_16_2/Y
+ VSUBS
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__inv_8_1/VGND sky130_fd_sc_hd__inv_8_1/VPWR VSUBS sky130_fd_sc_hd__inv_8_1/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_8_0 sky130_fd_sc_hd__inv_8_1/A sky130_fd_sc_hd__inv_8_1/Y sky130_fd_sc_hd__inv_8_1/VGND
+ sky130_fd_sc_hd__inv_8_1/VPWR VSUBS sky130_fd_sc_hd__inv_8_1/VPB sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__inv_8_1 sky130_fd_sc_hd__inv_8_1/A sky130_fd_sc_hd__inv_8_1/Y sky130_fd_sc_hd__inv_8_1/VGND
+ sky130_fd_sc_hd__inv_8_1/VPWR VSUBS sky130_fd_sc_hd__inv_8_1/VPB sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__inv_2_0 sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__inv_8_1/A sky130_fd_sc_hd__inv_8_1/VPWR
+ sky130_fd_sc_hd__inv_8_1/VGND VSUBS sky130_fd_sc_hd__inv_8_1/VPB sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_1 sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__inv_8_1/A sky130_fd_sc_hd__inv_8_1/VPWR
+ sky130_fd_sc_hd__inv_8_1/VGND VSUBS sky130_fd_sc_hd__inv_8_1/VPB sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__inv_8_1/VGND sky130_fd_sc_hd__inv_8_1/VPWR VSUBS sky130_fd_sc_hd__inv_8_1/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__inv_8_1/VGND sky130_fd_sc_hd__inv_8_1/VPWR VSUBS sky130_fd_sc_hd__inv_8_1/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__inv_8_1/Y
+ sky130_fd_sc_hd__inv_8_1/VGND sky130_fd_sc_hd__inv_8_1/VPWR VSUBS sky130_fd_sc_hd__inv_8_1/VPB
+ sky130_fd_sc_hd__inv_16
.ends

.subckt BR32 C[31] C[30] C[29] C[28] C[27] C[26] C[25] C[24] C[23] C[22] C[21] C[20]
+ C[19] C[18] C[17] C[16] C[15] C[14] C[13] C[12] C[11] C[10] C[9] C[8] C[7] C[6]
+ C[5] C[4] C[3] C[2] C[1] C[0] VSS VDD RESET OUT
Xbrbufhalf_32_0 C[20] C[30] OUT C[19] C[28] C[18] C[26] C[23] C[24] C[21] invcell_0/sky130_fd_sc_hd__inv_16_3/Y
+ C[29] C[17] VSS C[27] C[31] C[25] unitcell2buf_32_1/OUT brbufhalf_32_1/unitcell2buf_32_11/IN
+ C[22] invcell_0/sky130_fd_sc_hd__inv_16_2/Y unitcell2buf_32_1/RESET VSS VDD VSS
+ brbufhalf_32
Xbrbufhalf_32_1 C[3] C[13] brbufhalf_32_1/unitcell2bufcut_32_0/buf_out C[2] C[11]
+ C[1] C[9] C[6] C[7] C[4] invcell_0/sky130_fd_sc_hd__inv_16_2/Y C[12] C[0] VSS C[10]
+ C[14] C[8] brbufhalf_32_1/unitcell2buf_32_11/IN unitcell2buf_32_0/IN C[5] invcell_0/sky130_fd_sc_hd__inv_16_3/Y
+ brbufhalf_32_1/unitcell2buf_32_9/RESET VSS VDD VSS brbufhalf_32
Xinvcell_0 VSS invcell_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD RESET invcell_0/sky130_fd_sc_hd__inv_16_2/Y
+ VSS invcell
Xunitcell2buf_32_0 unitcell2buf_32_0/IN C[15] unitcell2buf_32_1/IN unitcell2buf_32_0/buf_out
+ VDD unitcell2buf_32_1/RESET VSS unitcell2buf_32
Xunitcell2buf_32_1 unitcell2buf_32_1/IN C[16] unitcell2buf_32_1/OUT unitcell2buf_32_1/buf_out
+ VDD unitcell2buf_32_1/RESET VSS unitcell2buf_32
.ends

.subckt sky130_fd_sc_hd__o22ai_1 A2 B1 Y A1 B2 VGND VPWR VNB VPB
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A1 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_307_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 A1 B1 Y VNB VPB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt unitcell_nbr sky130_fd_sc_hd__nor2_1_4/a_109_297# sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ sky130_fd_sc_hd__buf_1_4/X sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__buf_1_4/a_27_47#
+ sky130_fd_sc_hd__buf_1_4/A m1_746_156# sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__nor2_1_5/Y
+ sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__nor2_1_5/A sky130_fd_sc_hd__buf_1_5/VPB
+ li_n384_n810# li_n176_n810# sky130_fd_sc_hd__buf_1_5/X VSUBS sky130_fd_sc_hd__buf_1_5/A
+ sky130_fd_sc_hd__buf_1_5/a_27_47#
Xsky130_fd_sc_hd__buf_1_4 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_4/X
+ sky130_fd_sc_hd__buf_1_4/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_4/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__buf_1_5 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_5/X
+ sky130_fd_sc_hd__buf_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_5/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__inv_1#0_0 m1_746_156# sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ li_n176_n810# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1#0_1 li_n176_n810# sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ li_n384_n810# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__nor2_1_4/Y
+ sky130_fd_sc_hd__nor2_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ sky130_fd_sc_hd__nor2_1_4/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__nor2_1_5/Y
+ sky130_fd_sc_hd__nor2_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ sky130_fd_sc_hd__nor2_1_5/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__inv_1#0_3 li_n176_n810# sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ li_n384_n810# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1#0_2 m1_746_156# sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ li_n176_n810# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__nor2_1_2 sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__nor2_1_4/Y
+ sky130_fd_sc_hd__nor2_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ sky130_fd_sc_hd__nor2_1_4/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_3 sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__nor2_1_5/Y
+ sky130_fd_sc_hd__nor2_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ sky130_fd_sc_hd__nor2_1_5/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_4 sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__nor2_1_4/Y
+ sky130_fd_sc_hd__nor2_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ sky130_fd_sc_hd__nor2_1_4/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_5 sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__nor2_1_5/Y
+ sky130_fd_sc_hd__nor2_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ sky130_fd_sc_hd__nor2_1_5/a_109_297# sky130_fd_sc_hd__nor2_1
Xmux_0 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__buf_1_5/A
+ li_n176_n810# sky130_fd_sc_hd__nor2_1_5/Y m1_746_156# mux
Xmux_1 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__nor2_1_5/Y sky130_fd_sc_hd__buf_1_4/A
+ li_n176_n810# sky130_fd_sc_hd__nor2_1_4/Y m1_746_156# mux
Xmux_2 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__buf_1_5/A
+ li_n176_n810# sky130_fd_sc_hd__nor2_1_5/Y m1_746_156# mux
Xmux_3 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__nor2_1_5/Y sky130_fd_sc_hd__buf_1_4/A
+ li_n176_n810# sky130_fd_sc_hd__nor2_1_4/Y m1_746_156# mux
Xmux_4 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__buf_1_5/A
+ li_n176_n810# sky130_fd_sc_hd__nor2_1_5/Y m1_746_156# mux
Xmux_5 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__nor2_1_5/Y sky130_fd_sc_hd__buf_1_4/A
+ li_n176_n810# sky130_fd_sc_hd__nor2_1_4/Y m1_746_156# mux
Xsky130_fd_sc_hd__buf_1_0 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_4/X
+ sky130_fd_sc_hd__buf_1_4/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_4/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__buf_1_1 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_5/X
+ sky130_fd_sc_hd__buf_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_5/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__inv_1_1 li_n176_n810# sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ li_n384_n810# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1_0 m1_746_156# sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ li_n176_n810# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__buf_1_2 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_4/X
+ sky130_fd_sc_hd__buf_1_4/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_4/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__buf_1_3 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_5/X
+ sky130_fd_sc_hd__buf_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_5/a_27_47#
+ sky130_fd_sc_hd__buf_1
.ends

.subckt unitcell_nbr_cut sky130_fd_sc_hd__nor2_1_4/a_109_297# sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ sky130_fd_sc_hd__buf_1_4/X sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__buf_1_4/a_27_47#
+ li_n176_n810# sky130_fd_sc_hd__buf_1_4/A sky130_fd_sc_hd__nor2_1_5/Y m1_746_156#
+ sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__nor2_1_4/Y
+ sky130_fd_sc_hd__nor2_1_5/A li_n384_n810# sky130_fd_sc_hd__buf_1_5/X VSUBS sky130_fd_sc_hd__buf_1_5/A
+ sky130_fd_sc_hd__buf_1_5/a_27_47#
Xsky130_fd_sc_hd__buf_1_4 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_4/X
+ sky130_fd_sc_hd__buf_1_4/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_4/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__buf_1_5 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_5/X
+ sky130_fd_sc_hd__buf_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_5/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__inv_1#0_0 m1_746_156# sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ li_n176_n810# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1#0_1 li_n176_n810# sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ li_n384_n810# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__nor2_1_4/Y
+ sky130_fd_sc_hd__nor2_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ sky130_fd_sc_hd__nor2_1_4/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__nor2_1_5/Y
+ sky130_fd_sc_hd__nor2_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ sky130_fd_sc_hd__nor2_1_5/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__inv_1#0_3 li_n176_n810# sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ li_n384_n810# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1#0_2 m1_746_156# sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ li_n176_n810# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__nor2_1_2 sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__nor2_1_4/Y
+ sky130_fd_sc_hd__nor2_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ sky130_fd_sc_hd__nor2_1_4/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_3 sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__nor2_1_5/Y
+ sky130_fd_sc_hd__nor2_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ sky130_fd_sc_hd__nor2_1_5/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_4 sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__nor2_1_4/Y
+ sky130_fd_sc_hd__nor2_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ sky130_fd_sc_hd__nor2_1_4/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_5 sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__nor2_1_5/Y
+ sky130_fd_sc_hd__nor2_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ sky130_fd_sc_hd__nor2_1_5/a_109_297# sky130_fd_sc_hd__nor2_1
Xmux_0 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__buf_1_5/A
+ li_n176_n810# sky130_fd_sc_hd__nor2_1_5/Y m1_746_156# mux
Xmux_1 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__nor2_1_5/Y sky130_fd_sc_hd__buf_1_4/A
+ li_n176_n810# sky130_fd_sc_hd__nor2_1_4/Y m1_746_156# mux
Xmux_2 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__buf_1_5/A
+ li_n176_n810# sky130_fd_sc_hd__nor2_1_5/Y m1_746_156# mux
Xmux_3 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__nor2_1_5/Y sky130_fd_sc_hd__buf_1_4/A
+ li_n176_n810# sky130_fd_sc_hd__nor2_1_4/Y m1_746_156# mux
Xmux_4 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__buf_1_5/A
+ li_n176_n810# sky130_fd_sc_hd__nor2_1_5/Y m1_746_156# mux
Xmux_5 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__nor2_1_5/Y sky130_fd_sc_hd__buf_1_4/A
+ li_n176_n810# sky130_fd_sc_hd__nor2_1_4/Y m1_746_156# mux
Xsky130_fd_sc_hd__buf_1_0 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_4/X
+ sky130_fd_sc_hd__buf_1_4/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_4/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__buf_1_1 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_5/X
+ sky130_fd_sc_hd__buf_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_5/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__inv_1_1 li_n176_n810# sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ li_n384_n810# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1_0 m1_746_156# sky130_fd_sc_hd__buf_1_5/VPB VSUBS sky130_fd_sc_hd__buf_1_5/VPB
+ li_n176_n810# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__buf_1_2 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_4/X
+ sky130_fd_sc_hd__buf_1_4/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_4/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__buf_1_3 VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_5/X
+ sky130_fd_sc_hd__buf_1_5/A VSUBS sky130_fd_sc_hd__buf_1_5/VPB sky130_fd_sc_hd__buf_1_5/a_27_47#
+ sky130_fd_sc_hd__buf_1
.ends

.subckt nbrhalf unitcell_nbr_7/li_n384_n810# sky130_fd_sc_hd__inv_16_7/A unitcell_nbr_24/li_n384_n810#
+ unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/A unitcell_nbr_2/li_n384_n810# unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B
+ sky130_fd_sc_hd__inv_16_6/VGND unitcell_nbr_27/li_n384_n810# unitcell_nbr_5/li_n384_n810#
+ unitcell_nbr_cut_2/li_n384_n810# unitcell_nbr_8/li_n384_n810# unitcell_nbr_0/li_n384_n810#
+ unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/X sky130_fd_sc_hd__inv_16_7/VGND unitcell_nbr_25/li_n384_n810#
+ unitcell_nbr_3/li_n384_n810# sky130_fd_sc_hd__inv_16_4/VGND unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/A
+ unitcell_nbr_6/li_n384_n810# sky130_fd_sc_hd__inv_16_7/Y unitcell_nbr_cut_3/li_n384_n810#
+ unitcell_nbr_9/li_n384_n810# sky130_fd_sc_hd__inv_16_5/Y unitcell_nbr_1/li_n384_n810#
+ unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B unitcell_nbr_26/li_n384_n810# sky130_fd_sc_hd__inv_16_5/A
+ sky130_fd_sc_hd__inv_16_5/VGND unitcell_nbr_4/li_n384_n810# sky130_fd_sc_hd__inv_16_7/VPB
+ VSUBS
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/A
+ sky130_fd_sc_hd__inv_16_7/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_4 sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_5/A
+ sky130_fd_sc_hd__inv_16_4/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_5 sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_5/A
+ sky130_fd_sc_hd__inv_16_5/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_6 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/A
+ sky130_fd_sc_hd__inv_16_6/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_7 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/A
+ sky130_fd_sc_hd__inv_16_7/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell_nbr_20 unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_6/m1_746_156# unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_6/li_n384_n810# unitcell_nbr_6/li_n176_n810# unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_21 unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_7/m1_746_156# unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_7/li_n384_n810# unitcell_nbr_7/li_n176_n810# unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_10 unitcell_nbr_24/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_24/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_24/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_25/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_24/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_24/m1_746_156# unitcell_nbr_25/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_24/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_24/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_24/li_n384_n810# unitcell_nbr_24/li_n176_n810# unitcell_nbr_24/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_24/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_22 unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_8/m1_746_156# unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_8/li_n384_n810# unitcell_nbr_8/li_n176_n810# unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_11 unitcell_nbr_25/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_25/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_25/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_26/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_25/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_25/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_25/m1_746_156# unitcell_nbr_26/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_25/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_25/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_25/li_n384_n810# unitcell_nbr_25/li_n176_n810# unitcell_nbr_25/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_25/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_25/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_23 unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_9/m1_746_156# unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_9/li_n384_n810# unitcell_nbr_9/li_n176_n810# unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_24 unitcell_nbr_24/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_24/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_24/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_25/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_24/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_24/m1_746_156# unitcell_nbr_25/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_24/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_24/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_24/li_n384_n810# unitcell_nbr_24/li_n176_n810# unitcell_nbr_24/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_24/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_13 unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_27/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_27/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_27/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_27/m1_746_156# unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_27/li_n384_n810# unitcell_nbr_27/li_n176_n810# unitcell_nbr_27/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_27/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_27/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_12 unitcell_nbr_26/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_26/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_26/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_27/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_26/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_26/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_26/m1_746_156# unitcell_nbr_27/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_26/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_26/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_26/li_n384_n810# unitcell_nbr_26/li_n176_n810# unitcell_nbr_26/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_26/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_26/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_14 unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_0/m1_746_156# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_0/li_n384_n810# unitcell_nbr_0/li_n176_n810# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_25 unitcell_nbr_25/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_25/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_25/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_26/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_25/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_25/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_25/m1_746_156# unitcell_nbr_26/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_25/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_25/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_25/li_n384_n810# unitcell_nbr_25/li_n176_n810# unitcell_nbr_25/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_25/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_25/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_15 unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_1/m1_746_156# unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_1/li_n384_n810# unitcell_nbr_1/li_n176_n810# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_26 unitcell_nbr_26/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_26/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_26/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_27/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_26/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_26/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_26/m1_746_156# unitcell_nbr_27/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_26/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_26/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_26/li_n384_n810# unitcell_nbr_26/li_n176_n810# unitcell_nbr_26/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_26/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_26/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_16 unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_2/m1_746_156# unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_2/li_n384_n810# unitcell_nbr_2/li_n176_n810# unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_27 unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_27/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_27/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_27/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_27/m1_746_156# unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_27/li_n384_n810# unitcell_nbr_27/li_n176_n810# unitcell_nbr_27/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_27/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_27/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_17 unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_3/m1_746_156# unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_3/li_n384_n810# unitcell_nbr_3/li_n176_n810# unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_18 unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_4/m1_746_156# unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_4/li_n384_n810# unitcell_nbr_4/li_n176_n810# unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_0 unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_0/m1_746_156# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_0/li_n384_n810# unitcell_nbr_0/li_n176_n810# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_1 unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_1/m1_746_156# unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_1/li_n384_n810# unitcell_nbr_1/li_n176_n810# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_19 unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_5/m1_746_156# unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_5/li_n384_n810# unitcell_nbr_5/li_n176_n810# unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_2 unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_2/m1_746_156# unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_2/li_n384_n810# unitcell_nbr_2/li_n176_n810# unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_3 unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_3/m1_746_156# unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_3/li_n384_n810# unitcell_nbr_3/li_n176_n810# unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_4 unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_4/m1_746_156# unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_4/li_n384_n810# unitcell_nbr_4/li_n176_n810# unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_5 unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_5/m1_746_156# unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_5/li_n384_n810# unitcell_nbr_5/li_n176_n810# unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_cut_0 unitcell_nbr_cut_2/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_cut_2/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_cut_2/li_n176_n810#
+ unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/A unitcell_nbr_cut_2/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_cut_2/m1_746_156# sky130_fd_sc_hd__inv_16_7/VPB unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A
+ unitcell_nbr_cut_2/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y unitcell_nbr_cut_2/li_n384_n810#
+ unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/X VSUBS unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/A
+ unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/a_27_47# unitcell_nbr_cut
Xunitcell_nbr_6 unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_6/m1_746_156# unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_6/li_n384_n810# unitcell_nbr_6/li_n176_n810# unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_cut_2 unitcell_nbr_cut_2/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_cut_2/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_cut_2/li_n176_n810#
+ unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/A unitcell_nbr_cut_2/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_cut_2/m1_746_156# sky130_fd_sc_hd__inv_16_7/VPB unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A
+ unitcell_nbr_cut_2/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_5/Y unitcell_nbr_cut_2/li_n384_n810#
+ unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/X VSUBS unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/A
+ unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/a_27_47# unitcell_nbr_cut
Xunitcell_nbr_cut_1 unitcell_nbr_cut_3/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_cut_3/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_cut_3/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_cut_3/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_cut_3/li_n176_n810#
+ unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/B unitcell_nbr_cut_3/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_cut_3/m1_746_156# sky130_fd_sc_hd__inv_16_7/VPB unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/A
+ unitcell_nbr_cut_3/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y unitcell_nbr_cut_3/li_n384_n810#
+ unitcell_nbr_cut_3/sky130_fd_sc_hd__buf_1_5/X VSUBS unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/B
+ unitcell_nbr_cut_3/sky130_fd_sc_hd__buf_1_5/a_27_47# unitcell_nbr_cut
Xunitcell_nbr_7 unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_7/m1_746_156# unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_7/li_n384_n810# unitcell_nbr_7/li_n176_n810# unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_cut_3 unitcell_nbr_cut_3/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_cut_3/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_cut_3/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_cut_3/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_cut_3/li_n176_n810#
+ unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/B unitcell_nbr_cut_3/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_cut_3/m1_746_156# sky130_fd_sc_hd__inv_16_7/VPB unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/A
+ unitcell_nbr_cut_3/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y unitcell_nbr_cut_3/li_n384_n810#
+ unitcell_nbr_cut_3/sky130_fd_sc_hd__buf_1_5/X VSUBS unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/B
+ unitcell_nbr_cut_3/sky130_fd_sc_hd__buf_1_5/a_27_47# unitcell_nbr_cut
Xunitcell_nbr_8 unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_8/m1_746_156# unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_8/li_n384_n810# unitcell_nbr_8/li_n176_n810# unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_9 unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_9/m1_746_156# unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/VPB
+ unitcell_nbr_9/li_n384_n810# unitcell_nbr_9/li_n176_n810# unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_5/A
+ sky130_fd_sc_hd__inv_16_4/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_5/A
+ sky130_fd_sc_hd__inv_16_5/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/A
+ sky130_fd_sc_hd__inv_16_6/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
.ends

.subckt NBR128half nbrhalf_3/unitcell_nbr_9/li_n384_n810# nbrhalf_2/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/A
+ nbrhalf_3/unitcell_nbr_cut_2/li_n384_n810# nbrhalf_2/unitcell_nbr_3/li_n384_n810#
+ nbrhalf_3/unitcell_nbr_24/li_n384_n810# nbrhalf_0/unitcell_nbr_cut_3/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_2/li_n384_n810# nbrhalf_3/unitcell_nbr_1/li_n384_n810# nbrhalf_1/unitcell_nbr_8/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_6/li_n384_n810# nbrhalf_1/unitcell_nbr_0/li_n384_n810# nbrhalf_3/unitcell_nbr_27/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_25/li_n384_n810# nbrhalf_0/unitcell_nbr_5/li_n384_n810# nbrhalf_3/unitcell_nbr_4/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_3/li_n384_n810# nbrhalf_2/unitcell_nbr_9/li_n384_n810# nbrhalf_2/unitcell_nbr_cut_2/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_25/li_n384_n810# nbrhalf_2/unitcell_nbr_1/li_n384_n810# sky130_fd_sc_hd__inv_16_3/A
+ nbrhalf_3/unitcell_nbr_7/li_n384_n810# nbrhalf_0/unitcell_nbr_8/li_n384_n810# nbrhalf_0/unitcell_nbr_0/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_6/li_n384_n810# nbrhalf_0/unitcell_nbr_26/li_n384_n810# nbrhalf_3/unitcell_nbr_cut_3/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_4/li_n384_n810# nbrhalf_3/unitcell_nbr_25/li_n384_n810# nbrhalf_0/unitcell_nbr_3/li_n384_n810#
+ nbrhalf_3/unitcell_nbr_2/li_n384_n810# nbrhalf_1/unitcell_nbr_9/li_n384_n810# nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/A
+ nbrhalf_1/unitcell_nbr_cut_2/li_n384_n810# nbrhalf_1/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B
+ nbrhalf_2/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/A nbrhalf_1/unitcell_nbr_1/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_7/li_n384_n810# nbrhalf_3/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B
+ nbrhalf_1/unitcell_nbr_26/li_n384_n810# nbrhalf_3/unitcell_nbr_5/li_n384_n810# nbrhalf_0/unitcell_nbr_6/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_4/li_n384_n810# nbrhalf_2/unitcell_nbr_cut_3/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_2/li_n384_n810# nbrhalf_2/unitcell_nbr_26/li_n384_n810# nbrhalf_0/unitcell_nbr_24/li_n384_n810#
+ nbrhalf_3/unitcell_nbr_8/li_n384_n810# nbrhalf_0/unitcell_nbr_9/li_n384_n810# nbrhalf_0/unitcell_nbr_1/li_n384_n810#
+ nbrhalf_3/unitcell_nbr_0/li_n384_n810# nbrhalf_0/unitcell_nbr_cut_2/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_7/li_n384_n810# nbrhalf_3/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B
+ nbrhalf_2/unitcell_nbr_5/li_n384_n810# nbrhalf_0/unitcell_nbr_27/li_n384_n810# nbrhalf_1/unitcell_nbr_24/li_n384_n810#
+ nbrhalf_3/unitcell_nbr_26/li_n384_n810# nbrhalf_2/sky130_fd_sc_hd__inv_16_5/Y nbrhalf_0/unitcell_nbr_4/li_n384_n810#
+ nbrhalf_3/unitcell_nbr_3/li_n384_n810# nbrhalf_1/unitcell_nbr_cut_3/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_2/li_n384_n810# nbrhalf_2/unitcell_nbr_8/li_n384_n810# nbrhalf_1/unitcell_nbr_27/li_n384_n810#
+ sky130_fd_sc_hd__inv_16_3/VPB nbrhalf_2/unitcell_nbr_24/li_n384_n810# nbrhalf_2/unitcell_nbr_0/li_n384_n810#
+ nbrhalf_3/unitcell_nbr_6/li_n384_n810# nbrhalf_0/unitcell_nbr_7/li_n384_n810# nbrhalf_1/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B
+ nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/A nbrhalf_1/unitcell_nbr_5/li_n384_n810#
+ VSUBS nbrhalf_0/unitcell_nbr_25/li_n384_n810# nbrhalf_2/unitcell_nbr_27/li_n384_n810#
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xnbrhalf_0 nbrhalf_0/unitcell_nbr_7/li_n384_n810# sky130_fd_sc_hd__inv_16_3/Y nbrhalf_0/unitcell_nbr_24/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/A nbrhalf_0/unitcell_nbr_2/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B VSUBS nbrhalf_0/unitcell_nbr_27/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_5/li_n384_n810# nbrhalf_0/unitcell_nbr_cut_2/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_8/li_n384_n810# nbrhalf_0/unitcell_nbr_0/li_n384_n810# nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS nbrhalf_0/unitcell_nbr_25/li_n384_n810# nbrhalf_0/unitcell_nbr_3/li_n384_n810#
+ VSUBS nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/A nbrhalf_0/unitcell_nbr_6/li_n384_n810#
+ nbrhalf_0/sky130_fd_sc_hd__inv_16_7/Y nbrhalf_0/unitcell_nbr_cut_3/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_9/li_n384_n810# nbrhalf_0/sky130_fd_sc_hd__inv_16_5/Y nbrhalf_0/unitcell_nbr_1/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B nbrhalf_0/unitcell_nbr_26/li_n384_n810#
+ sky130_fd_sc_hd__inv_16_3/Y VSUBS nbrhalf_0/unitcell_nbr_4/li_n384_n810# sky130_fd_sc_hd__inv_16_3/VPB
+ VSUBS nbrhalf
Xnbrhalf_1 nbrhalf_1/unitcell_nbr_7/li_n384_n810# sky130_fd_sc_hd__inv_16_1/Y nbrhalf_1/unitcell_nbr_24/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B nbrhalf_1/unitcell_nbr_2/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B VSUBS nbrhalf_1/unitcell_nbr_27/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_5/li_n384_n810# nbrhalf_1/unitcell_nbr_cut_2/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_8/li_n384_n810# nbrhalf_1/unitcell_nbr_0/li_n384_n810# nbrhalf_1/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS nbrhalf_1/unitcell_nbr_25/li_n384_n810# nbrhalf_1/unitcell_nbr_3/li_n384_n810#
+ VSUBS nbrhalf_0/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B nbrhalf_1/unitcell_nbr_6/li_n384_n810#
+ nbrhalf_1/sky130_fd_sc_hd__inv_16_7/Y nbrhalf_1/unitcell_nbr_cut_3/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_9/li_n384_n810# nbrhalf_1/sky130_fd_sc_hd__inv_16_5/Y nbrhalf_1/unitcell_nbr_1/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B nbrhalf_1/unitcell_nbr_26/li_n384_n810#
+ sky130_fd_sc_hd__inv_16_1/Y VSUBS nbrhalf_1/unitcell_nbr_4/li_n384_n810# sky130_fd_sc_hd__inv_16_3/VPB
+ VSUBS nbrhalf
Xnbrhalf_2 nbrhalf_2/unitcell_nbr_7/li_n384_n810# sky130_fd_sc_hd__inv_16_1/Y nbrhalf_2/unitcell_nbr_24/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/A nbrhalf_2/unitcell_nbr_2/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B VSUBS nbrhalf_2/unitcell_nbr_27/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_5/li_n384_n810# nbrhalf_2/unitcell_nbr_cut_2/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_8/li_n384_n810# nbrhalf_2/unitcell_nbr_0/li_n384_n810# nbrhalf_2/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS nbrhalf_2/unitcell_nbr_25/li_n384_n810# nbrhalf_2/unitcell_nbr_3/li_n384_n810#
+ VSUBS nbrhalf_2/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/A nbrhalf_2/unitcell_nbr_6/li_n384_n810#
+ nbrhalf_2/sky130_fd_sc_hd__inv_16_7/Y nbrhalf_2/unitcell_nbr_cut_3/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_9/li_n384_n810# nbrhalf_2/sky130_fd_sc_hd__inv_16_5/Y nbrhalf_2/unitcell_nbr_1/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B nbrhalf_2/unitcell_nbr_26/li_n384_n810#
+ sky130_fd_sc_hd__inv_16_1/Y VSUBS nbrhalf_2/unitcell_nbr_4/li_n384_n810# sky130_fd_sc_hd__inv_16_3/VPB
+ VSUBS nbrhalf
Xnbrhalf_3 nbrhalf_3/unitcell_nbr_7/li_n384_n810# sky130_fd_sc_hd__inv_16_3/Y nbrhalf_3/unitcell_nbr_24/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B nbrhalf_3/unitcell_nbr_2/li_n384_n810#
+ nbrhalf_3/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B VSUBS nbrhalf_3/unitcell_nbr_27/li_n384_n810#
+ nbrhalf_3/unitcell_nbr_5/li_n384_n810# nbrhalf_3/unitcell_nbr_cut_2/li_n384_n810#
+ nbrhalf_3/unitcell_nbr_8/li_n384_n810# nbrhalf_3/unitcell_nbr_0/li_n384_n810# nbrhalf_3/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS nbrhalf_3/unitcell_nbr_25/li_n384_n810# nbrhalf_3/unitcell_nbr_3/li_n384_n810#
+ VSUBS nbrhalf_2/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B nbrhalf_3/unitcell_nbr_6/li_n384_n810#
+ nbrhalf_3/sky130_fd_sc_hd__inv_16_7/Y nbrhalf_3/unitcell_nbr_cut_3/li_n384_n810#
+ nbrhalf_3/unitcell_nbr_9/li_n384_n810# nbrhalf_3/sky130_fd_sc_hd__inv_16_5/Y nbrhalf_3/unitcell_nbr_1/li_n384_n810#
+ nbrhalf_3/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B nbrhalf_3/unitcell_nbr_26/li_n384_n810#
+ sky130_fd_sc_hd__inv_16_3/Y VSUBS nbrhalf_3/unitcell_nbr_4/li_n384_n810# sky130_fd_sc_hd__inv_16_3/VPB
+ VSUBS nbrhalf
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
.ends

.subckt nbrhalf_128 unitcell_nbr_7/li_n384_n810# sky130_fd_sc_hd__inv_16_3/A unitcell_nbr_10/li_n384_n810#
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_4/A unitcell_nbr_2/li_n384_n810# unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_5/B
+ sky130_fd_sc_hd__inv_16_2/VGND unitcell_nbr_5/li_n384_n810# unitcell_nbr_8/li_n384_n810#
+ unitcell_nbr_cut_0/li_n384_n810# unitcell_nbr_0/li_n384_n810# sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_3/VGND unitcell_nbr_11/li_n384_n810# unitcell_nbr_3/li_n384_n810#
+ sky130_fd_sc_hd__inv_16_0/VGND unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_4/B
+ unitcell_nbr_6/li_n384_n810# sky130_fd_sc_hd__inv_16_3/VPB unitcell_nbr_9/li_n384_n810#
+ unitcell_nbr_cut_1/li_n384_n810# unitcell_nbr_1/li_n384_n810# unitcell_nbr_12/li_n384_n810#
+ sky130_fd_sc_hd__inv_16_1/VGND unitcell_nbr_4/li_n384_n810# VSUBS
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16_3/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell_nbr_10 unitcell_nbr_10/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_10/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_10/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_11/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_10/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_10/m1_746_156# unitcell_nbr_11/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_10/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_10/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_10/li_n384_n810# unitcell_nbr_10/li_n176_n810# unitcell_nbr_10/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_10/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_11 unitcell_nbr_11/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_11/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_11/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_12/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_11/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_11/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_11/m1_746_156# unitcell_nbr_12/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_11/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_11/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_11/li_n384_n810# unitcell_nbr_11/li_n176_n810# unitcell_nbr_11/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_11/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_11/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_12 unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_12/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_12/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_12/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_12/m1_746_156# unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_12/li_n384_n810# unitcell_nbr_12/li_n176_n810# unitcell_nbr_12/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_12/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_12/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_0 unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_0/m1_746_156# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_0/li_n384_n810# unitcell_nbr_0/li_n176_n810# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_1 unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_1/m1_746_156# unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_1/li_n384_n810# unitcell_nbr_1/li_n176_n810# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_2 unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_2/m1_746_156# unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_2/li_n384_n810# unitcell_nbr_2/li_n176_n810# unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_3 unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_3/m1_746_156# unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_3/li_n384_n810# unitcell_nbr_3/li_n176_n810# unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_4 unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_4/m1_746_156# unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_4/li_n384_n810# unitcell_nbr_4/li_n176_n810# unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_5 unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_5/m1_746_156# unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_5/li_n384_n810# unitcell_nbr_5/li_n176_n810# unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_cut_0 unitcell_nbr_cut_0/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_cut_0/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_cut_0/li_n176_n810#
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_4/A unitcell_nbr_cut_0/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_cut_0/m1_746_156# sky130_fd_sc_hd__inv_16_3/VPB unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y unitcell_nbr_cut_0/li_n384_n810#
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_5/X VSUBS unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_5/A
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_5/a_27_47# unitcell_nbr_cut
Xunitcell_nbr_6 unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_6/m1_746_156# unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_6/li_n384_n810# unitcell_nbr_6/li_n176_n810# unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_cut_1 unitcell_nbr_cut_1/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_cut_1/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_cut_1/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_cut_1/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_cut_1/li_n176_n810#
+ unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/B unitcell_nbr_cut_1/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_cut_1/m1_746_156# sky130_fd_sc_hd__inv_16_3/VPB unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/A
+ unitcell_nbr_cut_1/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y unitcell_nbr_cut_1/li_n384_n810#
+ unitcell_nbr_cut_1/sky130_fd_sc_hd__buf_1_5/X VSUBS unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/B
+ unitcell_nbr_cut_1/sky130_fd_sc_hd__buf_1_5/a_27_47# unitcell_nbr_cut
Xunitcell_nbr_7 unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_7/m1_746_156# unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_7/li_n384_n810# unitcell_nbr_7/li_n176_n810# unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_8 unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_8/m1_746_156# unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_8/li_n384_n810# unitcell_nbr_8/li_n176_n810# unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_9 unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_9/m1_746_156# unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_9/li_n384_n810# unitcell_nbr_9/li_n176_n810# unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_0/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_1/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16_2/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
.ends

.subckt NBR128half_bottom nbrhalf_2/unitcell_nbr_3/li_n384_n810# nbrhalf_128_0/unitcell_nbr_0/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_cut_3/li_n384_n810# nbrhalf_0/unitcell_nbr_2/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_8/li_n384_n810# nbrhalf_1/unitcell_nbr_0/li_n384_n810# nbrhalf_2/unitcell_nbr_6/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_25/li_n384_n810# nbrhalf_128_0/unitcell_nbr_3/li_n384_n810#
+ nbrhalf_128_0/unitcell_nbr_10/li_n384_n810# nbrhalf_0/unitcell_nbr_5/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_3/li_n384_n810# nbrhalf_2/unitcell_nbr_9/li_n384_n810# nbrhalf_2/unitcell_nbr_cut_2/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/A nbrhalf_128_0/unitcell_nbr_6/li_n384_n810#
+ nbrhalf_128_0/unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_4/B nbrhalf_2/unitcell_nbr_25/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_1/li_n384_n810# sky130_fd_sc_hd__inv_16_3/A nbrhalf_0/unitcell_nbr_8/li_n384_n810#
+ nbrhalf_128_0/unitcell_nbr_cut_0/li_n384_n810# nbrhalf_0/unitcell_nbr_0/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_6/li_n384_n810# nbrhalf_128_0/unitcell_nbr_9/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_26/li_n384_n810# nbrhalf_2/unitcell_nbr_4/li_n384_n810# nbrhalf_128_0/unitcell_nbr_1/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_3/li_n384_n810# nbrhalf_1/unitcell_nbr_9/li_n384_n810# nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/A
+ nbrhalf_1/unitcell_nbr_cut_2/li_n384_n810# nbrhalf_1/unitcell_nbr_1/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_7/li_n384_n810# nbrhalf_1/unitcell_nbr_26/li_n384_n810# nbrhalf_128_0/unitcell_nbr_4/li_n384_n810#
+ nbrhalf_128_0/unitcell_nbr_11/li_n384_n810# nbrhalf_0/unitcell_nbr_6/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_4/li_n384_n810# nbrhalf_2/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B
+ nbrhalf_2/unitcell_nbr_cut_3/li_n384_n810# nbrhalf_128_0/unitcell_nbr_7/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_26/li_n384_n810# nbrhalf_0/unitcell_nbr_24/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_2/li_n384_n810# nbrhalf_0/unitcell_nbr_9/li_n384_n810# nbrhalf_0/unitcell_nbr_cut_2/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_1/li_n384_n810# nbrhalf_128_0/unitcell_nbr_cut_1/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_7/li_n384_n810# nbrhalf_1/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/A
+ nbrhalf_2/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B nbrhalf_0/unitcell_nbr_27/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_5/li_n384_n810# nbrhalf_1/unitcell_nbr_24/li_n384_n810# nbrhalf_128_0/unitcell_nbr_2/li_n384_n810#
+ nbrhalf_128_0/unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_5/B nbrhalf_0/unitcell_nbr_4/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_cut_3/li_n384_n810# nbrhalf_1/unitcell_nbr_2/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_8/li_n384_n810# nbrhalf_1/unitcell_nbr_27/li_n384_n810# nbrhalf_128_0/unitcell_nbr_5/li_n384_n810#
+ nbrhalf_128_0/unitcell_nbr_12/li_n384_n810# nbrhalf_2/unitcell_nbr_24/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_0/li_n384_n810# nbrhalf_0/unitcell_nbr_7/li_n384_n810# nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/A
+ nbrhalf_1/unitcell_nbr_5/li_n384_n810# sky130_fd_sc_hd__inv_16_3/VPB nbrhalf_128_0/unitcell_nbr_8/li_n384_n810#
+ VSUBS nbrhalf_2/unitcell_nbr_27/li_n384_n810# nbrhalf_0/unitcell_nbr_25/li_n384_n810#
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xnbrhalf_0 nbrhalf_0/unitcell_nbr_7/li_n384_n810# sky130_fd_sc_hd__inv_16_3/Y nbrhalf_0/unitcell_nbr_24/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/A nbrhalf_0/unitcell_nbr_2/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B VSUBS nbrhalf_0/unitcell_nbr_27/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_5/li_n384_n810# nbrhalf_0/unitcell_nbr_cut_2/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_8/li_n384_n810# nbrhalf_0/unitcell_nbr_0/li_n384_n810# nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS nbrhalf_0/unitcell_nbr_25/li_n384_n810# nbrhalf_0/unitcell_nbr_3/li_n384_n810#
+ VSUBS nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/A nbrhalf_0/unitcell_nbr_6/li_n384_n810#
+ nbrhalf_0/sky130_fd_sc_hd__inv_16_7/Y nbrhalf_0/unitcell_nbr_cut_3/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_9/li_n384_n810# nbrhalf_0/sky130_fd_sc_hd__inv_16_5/Y nbrhalf_0/unitcell_nbr_1/li_n384_n810#
+ nbrhalf_0/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B nbrhalf_0/unitcell_nbr_26/li_n384_n810#
+ sky130_fd_sc_hd__inv_16_3/Y VSUBS nbrhalf_0/unitcell_nbr_4/li_n384_n810# sky130_fd_sc_hd__inv_16_3/VPB
+ VSUBS nbrhalf
Xnbrhalf_1 nbrhalf_1/unitcell_nbr_7/li_n384_n810# sky130_fd_sc_hd__inv_16_1/Y nbrhalf_1/unitcell_nbr_24/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/A nbrhalf_1/unitcell_nbr_2/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B VSUBS nbrhalf_1/unitcell_nbr_27/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_5/li_n384_n810# nbrhalf_1/unitcell_nbr_cut_2/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_8/li_n384_n810# nbrhalf_1/unitcell_nbr_0/li_n384_n810# nbrhalf_1/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS nbrhalf_1/unitcell_nbr_25/li_n384_n810# nbrhalf_1/unitcell_nbr_3/li_n384_n810#
+ VSUBS nbrhalf_1/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/A nbrhalf_1/unitcell_nbr_6/li_n384_n810#
+ nbrhalf_1/sky130_fd_sc_hd__inv_16_7/Y nbrhalf_1/unitcell_nbr_cut_3/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_9/li_n384_n810# nbrhalf_1/sky130_fd_sc_hd__inv_16_5/Y nbrhalf_1/unitcell_nbr_1/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B nbrhalf_1/unitcell_nbr_26/li_n384_n810#
+ sky130_fd_sc_hd__inv_16_1/Y VSUBS nbrhalf_1/unitcell_nbr_4/li_n384_n810# sky130_fd_sc_hd__inv_16_3/VPB
+ VSUBS nbrhalf
Xnbrhalf_2 nbrhalf_2/unitcell_nbr_7/li_n384_n810# sky130_fd_sc_hd__inv_16_3/Y nbrhalf_2/unitcell_nbr_24/li_n384_n810#
+ nbrhalf_1/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B nbrhalf_2/unitcell_nbr_2/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B VSUBS nbrhalf_2/unitcell_nbr_27/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_5/li_n384_n810# nbrhalf_2/unitcell_nbr_cut_2/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_8/li_n384_n810# nbrhalf_2/unitcell_nbr_0/li_n384_n810# nbrhalf_2/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS nbrhalf_2/unitcell_nbr_25/li_n384_n810# nbrhalf_2/unitcell_nbr_3/li_n384_n810#
+ VSUBS nbrhalf_1/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B nbrhalf_2/unitcell_nbr_6/li_n384_n810#
+ nbrhalf_2/sky130_fd_sc_hd__inv_16_7/Y nbrhalf_2/unitcell_nbr_cut_3/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_9/li_n384_n810# nbrhalf_2/sky130_fd_sc_hd__inv_16_5/Y nbrhalf_2/unitcell_nbr_1/li_n384_n810#
+ nbrhalf_2/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B nbrhalf_2/unitcell_nbr_26/li_n384_n810#
+ sky130_fd_sc_hd__inv_16_3/Y VSUBS nbrhalf_2/unitcell_nbr_4/li_n384_n810# sky130_fd_sc_hd__inv_16_3/VPB
+ VSUBS nbrhalf
Xnbrhalf_128_0 nbrhalf_128_0/unitcell_nbr_7/li_n384_n810# sky130_fd_sc_hd__inv_16_1/Y
+ nbrhalf_128_0/unitcell_nbr_10/li_n384_n810# nbrhalf_0/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B
+ nbrhalf_128_0/unitcell_nbr_2/li_n384_n810# nbrhalf_128_0/unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_5/B
+ VSUBS nbrhalf_128_0/unitcell_nbr_5/li_n384_n810# nbrhalf_128_0/unitcell_nbr_8/li_n384_n810#
+ nbrhalf_128_0/unitcell_nbr_cut_0/li_n384_n810# nbrhalf_128_0/unitcell_nbr_0/li_n384_n810#
+ sky130_fd_sc_hd__inv_16_1/Y VSUBS nbrhalf_128_0/unitcell_nbr_11/li_n384_n810# nbrhalf_128_0/unitcell_nbr_3/li_n384_n810#
+ VSUBS nbrhalf_0/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B nbrhalf_128_0/unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_4/B
+ nbrhalf_128_0/unitcell_nbr_6/li_n384_n810# sky130_fd_sc_hd__inv_16_3/VPB nbrhalf_128_0/unitcell_nbr_9/li_n384_n810#
+ nbrhalf_128_0/unitcell_nbr_cut_1/li_n384_n810# nbrhalf_128_0/unitcell_nbr_1/li_n384_n810#
+ nbrhalf_128_0/unitcell_nbr_12/li_n384_n810# VSUBS nbrhalf_128_0/unitcell_nbr_4/li_n384_n810#
+ VSUBS nbrhalf_128
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
.ends

.subckt NBR128 RESET C[0] C[1] C[2] C[3] C[4] C[5] C[7] C[8] C[9] C[10] C[11] C[12]
+ C[13] C[14] C[15] C[16] C[17] C[18] C[19] C[20] C[21] C[22] C[23] C[24] C[25] C[26]
+ C[27] C[28] C[29] C[30] C[6] C[31] C[32] C[33] C[34] C[35] C[36] C[37] C[38] C[39]
+ C[40] C[41] C[42] C[43] C[44] C[45] C[46] C[47] C[48] C[49] C[50] C[51] C[52] C[53]
+ C[54] C[55] C[56] C[57] C[58] C[59] C[60] C[61] C[62] C[95] C[96] C[97] C[98] C[99]
+ C[100] C[101] C[102] C[103] C[104] C[105] C[106] C[107] C[108] C[109] C[110] C[111]
+ C[112] C[113] C[114] C[115] C[116] C[117] C[118] C[119] C[120] C[121] C[122] C[123]
+ C[124] C[125] C[126] C[127] C[63] C[64] C[65] C[66] C[67] C[68] C[69] C[70] C[71]
+ C[72] C[73] C[74] C[75] C[76] C[77] C[78] C[79] C[80] C[81] C[82] C[83] C[84] C[85]
+ C[86] C[87] C[88] C[89] C[90] C[91] C[92] C[93] C[94] OUT VDD VSS
Xsky130_fd_sc_hd__inv_8_0 sky130_fd_sc_hd__inv_8_0/A sky130_fd_sc_hd__inv_8_0/Y VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__buf_2_0 VDD VSS sky130_fd_sc_hd__inv_8_0/A RESET VSS VDD sky130_fd_sc_hd__buf_2
Xunitcell_nbr_0 unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_0/m1_746_156# unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/Y unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/A
+ VDD C[127] unitcell_nbr_0/li_n176_n810# OUT VSS unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/a_27_47# unitcell_nbr
XNBR128half_0 C[99] unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/B C[110] C[122] C[98]
+ C[23] C[28] C[108] C[5] C[119] C[14] C[95] C[2] C[25] C[105] C[11] C[115] C[126]
+ C[113] C[124] sky130_fd_sc_hd__inv_16_1/Y C[101] C[21] C[30] C[8] C[17] C[102] C[121]
+ C[97] C[27] C[107] C[4] NBR128half_0/nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/A
+ C[15] unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/B
+ C[13] C[117] NBR128half_0/nbrhalf_3/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B
+ C[1] C[104] C[24] C[10] C[118] C[123] C[112] C[19] C[100] C[20] C[29] C[109] C[31]
+ C[6] NBR128half_0/nbrhalf_3/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B C[120] C[16]
+ C[3] C[96] unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/A C[26] C[106] C[7] C[12] C[116]
+ C[0] VDD C[114] C[125] C[103] C[22] unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A NBR128half_0/nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/A
+ C[9] VSS C[18] C[111] NBR128half
XNBR128half_bottom_0 C[74] C[45] C[54] C[59] C[84] C[93] C[71] C[81] C[42] C[34] C[56]
+ C[90] C[67] C[78] NBR128half_0/nbrhalf_3/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B
+ C[39] NBR128half_0/nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/A C[65]
+ C[76] sky130_fd_sc_hd__inv_16_1/Y C[52] C[46] C[61] C[87] C[35] C[48] C[73] C[44]
+ C[58] C[83] NBR128half_bottom_0/nbrhalf_2/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B
+ C[94] C[92] C[69] C[80] C[41] C[33] C[55] C[89] NBR128half_bottom_0/nbrhalf_2/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B
+ C[70] C[37] C[64] C[50] C[75] C[51] C[62] C[60] C[38] C[85] NBR128half_0/nbrhalf_3/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B
+ NBR128half_bottom_0/nbrhalf_2/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B C[47]
+ C[72] C[82] C[43] NBR128half_0/nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/A
+ C[57] C[86] C[91] C[68] C[79] C[40] C[32] C[66] C[77] C[53] NBR128half_bottom_0/nbrhalf_2/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B
+ C[88] VDD C[36] VSS C[63] C[49] NBR128half_bottom
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_8_0/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_8_0/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
.ends

.subckt nbrhalf_64 unitcell_nbr_7/li_n384_n810# unitcell_nbr_10/li_n384_n810# unitcell_nbr_2/li_n384_n810#
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A unitcell_nbr_13/li_n384_n810# unitcell_nbr_13/sky130_fd_sc_hd__nor2_1_4/B
+ sky130_fd_sc_hd__inv_16_2/VGND unitcell_nbr_5/li_n384_n810# unitcell_nbr_cut_0/li_n384_n810#
+ unitcell_nbr_8/li_n384_n810# unitcell_nbr_0/li_n384_n810# sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16_1/A unitcell_nbr_11/li_n384_n810# sky130_fd_sc_hd__inv_16_3/VGND
+ unitcell_nbr_3/li_n384_n810# sky130_fd_sc_hd__inv_16_0/VGND unitcell_nbr_6/li_n384_n810#
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_9/li_n384_n810# unitcell_nbr_1/li_n384_n810#
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell_nbr_13/sky130_fd_sc_hd__nor2_1_5/B unitcell_nbr_12/li_n384_n810#
+ unitcell_nbr_4/li_n384_n810# sky130_fd_sc_hd__inv_16_1/VGND VSUBS
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16_3/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell_nbr_10 unitcell_nbr_10/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_10/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_10/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_11/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_10/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_10/m1_746_156# unitcell_nbr_11/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_10/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_10/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_10/li_n384_n810# unitcell_nbr_10/li_n176_n810# unitcell_nbr_10/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_10/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_11 unitcell_nbr_11/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_11/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_11/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_12/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_11/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_11/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_11/m1_746_156# unitcell_nbr_12/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_11/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_11/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_11/li_n384_n810# unitcell_nbr_11/li_n176_n810# unitcell_nbr_11/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_11/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_11/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_13 unitcell_nbr_13/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_13/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_13/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_13/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_13/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_13/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_13/m1_746_156# unitcell_nbr_13/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_13/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_13/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_13/li_n384_n810# unitcell_nbr_13/li_n176_n810# unitcell_nbr_13/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_13/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_13/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_12 unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_12/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_13/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_12/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_12/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_12/m1_746_156# unitcell_nbr_13/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_12/li_n384_n810# unitcell_nbr_12/li_n176_n810# unitcell_nbr_12/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_12/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_12/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_0 unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_0/m1_746_156# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_0/li_n384_n810# unitcell_nbr_0/li_n176_n810# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_1 unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_1/m1_746_156# unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_1/li_n384_n810# unitcell_nbr_1/li_n176_n810# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_2 unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_2/m1_746_156# unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_2/li_n384_n810# unitcell_nbr_2/li_n176_n810# unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_3 unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_3/m1_746_156# unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_3/li_n384_n810# unitcell_nbr_3/li_n176_n810# unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_4 unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_4/m1_746_156# unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_4/li_n384_n810# unitcell_nbr_4/li_n176_n810# unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_5 unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_5/m1_746_156# unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_5/li_n384_n810# unitcell_nbr_5/li_n176_n810# unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_6 unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_6/m1_746_156# unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_6/li_n384_n810# unitcell_nbr_6/li_n176_n810# unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_cut_0 unitcell_nbr_cut_0/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_cut_0/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_cut_0/li_n176_n810#
+ unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/B unitcell_nbr_cut_0/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_cut_0/m1_746_156# sky130_fd_sc_hd__inv_16_3/VPB unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/A
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y unitcell_nbr_cut_0/li_n384_n810#
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_5/X VSUBS unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/B
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_5/a_27_47# unitcell_nbr_cut
Xunitcell_nbr_7 unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_7/m1_746_156# unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_7/li_n384_n810# unitcell_nbr_7/li_n176_n810# unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_8 unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_8/m1_746_156# unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_8/li_n384_n810# unitcell_nbr_8/li_n176_n810# unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_9 unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_9/m1_746_156# unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_9/li_n384_n810# unitcell_nbr_9/li_n176_n810# unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_0/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_1/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16_2/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
.ends

.subckt NBR64 OUT VDD RESET C[0] C[1] C[2] C[3] C[4] C[5] C[6] C[7] C[8] C[9] C[10]
+ C[11] C[12] C[13] C[14] C[15] C[16] C[17] C[18] C[19] C[20] C[21] C[22] C[23] C[24]
+ C[25] C[26] C[27] C[28] C[29] C[30] C[31] C[32] C[33] C[34] C[35] C[36] C[37] C[38]
+ C[39] C[40] C[41] C[42] C[43] C[44] C[45] C[46] C[47] C[48] C[49] C[50] C[51] C[52]
+ C[53] C[54] C[55] C[56] C[57] C[58] C[59] C[60] C[61] C[62] C[63] VSS
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__inv_16_4/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_4 sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__inv_16_4/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xnbrhalf_64_0 C[22] C[19] C[28] unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/B C[16] nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/A
+ VSS C[25] C[23] C[21] C[30] sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__inv_16_4/Y
+ C[18] VSS C[27] VSS C[24] unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/B C[20] C[29]
+ VDD nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/A C[17] C[26] VSS VSS
+ nbrhalf_64
Xsky130_fd_sc_hd__inv_4_0 sky130_fd_sc_hd__inv_4_0/Y RESET VDD VSS VSS VDD sky130_fd_sc_hd__inv_4
Xnbrhalf_0 C[6] sky130_fd_sc_hd__inv_16_2/Y C[3] nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_4/A
+ C[12] nbrhalf_0/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B VSS C[0] C[9] C[15]
+ C[5] C[14] nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/X VSS C[2] C[11]
+ VSS nbrhalf_0/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/A C[8] nbrhalf_0/sky130_fd_sc_hd__inv_16_7/Y
+ C[7] C[4] nbrhalf_0/sky130_fd_sc_hd__inv_16_5/Y C[13] nbrhalf_0/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B
+ C[1] sky130_fd_sc_hd__inv_16_2/Y VSS C[10] VDD VSS nbrhalf
Xnbrhalf_1 C[54] sky130_fd_sc_hd__inv_16_2/Y C[51] nbrhalf_0/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B
+ C[60] nbrhalf_1/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B VSS C[48] C[57] C[63]
+ C[53] C[62] OUT VSS C[50] C[59] VSS nbrhalf_0/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B
+ C[56] nbrhalf_1/sky130_fd_sc_hd__inv_16_7/Y C[55] C[52] nbrhalf_1/sky130_fd_sc_hd__inv_16_5/Y
+ C[61] nbrhalf_1/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B C[49] sky130_fd_sc_hd__inv_16_2/Y
+ VSS C[58] VDD VSS nbrhalf
Xnbrhalf_2 C[38] sky130_fd_sc_hd__inv_16_4/Y C[35] nbrhalf_1/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_5/B
+ C[44] unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A VSS C[32] C[41] C[47] C[37] C[46]
+ nbrhalf_2/unitcell_nbr_cut_2/sky130_fd_sc_hd__buf_1_5/X VSS C[34] C[43] VSS nbrhalf_1/unitcell_nbr_27/sky130_fd_sc_hd__nor2_1_4/B
+ C[40] nbrhalf_2/sky130_fd_sc_hd__inv_16_7/Y C[39] C[36] nbrhalf_2/sky130_fd_sc_hd__inv_16_5/Y
+ C[45] unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A C[33] sky130_fd_sc_hd__inv_16_4/Y
+ VSS C[42] VDD VSS nbrhalf
Xunitcell_nbr_0 unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_0/m1_746_156# unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/Y nbrhalf_2/sky130_fd_sc_hd__inv_16_7/Y
+ VDD C[31] unitcell_nbr_0/li_n176_n810# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/X
+ VSS unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_4_0/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__inv_16_4/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__inv_16_4/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
.ends

.subckt nbrhalf_32 unitcell_nbr_7/li_n384_n810# unitcell_nbr_10/li_n384_n810# unitcell_nbr_2/li_n384_n810#
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_4/A unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_5/X
+ unitcell_nbr_5/li_n384_n810# unitcell_nbr_cut_0/li_n384_n810# unitcell_nbr_8/li_n384_n810#
+ unitcell_nbr_0/li_n384_n810# unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_11/li_n384_n810# sky130_fd_sc_hd__inv_16_3/VGND unitcell_nbr_3/li_n384_n810#
+ sky130_fd_sc_hd__inv_16_3/A unitcell_nbr_6/li_n384_n810# sky130_fd_sc_hd__inv_16_3/Y
+ unitcell_nbr_9/li_n384_n810# unitcell_nbr_cut_1/li_n384_n810# unitcell_nbr_1/li_n384_n810#
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell_nbr_12/li_n384_n810# sky130_fd_sc_hd__inv_16_1/A
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_4/li_n384_n810# sky130_fd_sc_hd__inv_16_1/VGND
+ VSUBS
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16_3/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell_nbr_10 unitcell_nbr_10/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_10/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_10/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_11/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_10/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_10/m1_746_156# unitcell_nbr_11/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_10/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_10/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_10/li_n384_n810# unitcell_nbr_10/li_n176_n810# unitcell_nbr_10/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_10/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_11 unitcell_nbr_11/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_11/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_11/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_12/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_11/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_11/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_11/m1_746_156# unitcell_nbr_12/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_11/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_11/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_11/li_n384_n810# unitcell_nbr_11/li_n176_n810# unitcell_nbr_11/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_11/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_11/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_12 unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_12/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_12/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_12/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_12/m1_746_156# unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_12/li_n384_n810# unitcell_nbr_12/li_n176_n810# unitcell_nbr_12/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_12/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_12/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_0 unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_0/m1_746_156# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_0/li_n384_n810# unitcell_nbr_0/li_n176_n810# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_1 unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_1/m1_746_156# unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_1/li_n384_n810# unitcell_nbr_1/li_n176_n810# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_2 unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_2/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_2/m1_746_156# unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_2/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_2/li_n384_n810# unitcell_nbr_2/li_n176_n810# unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_2/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_3 unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_3/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_3/m1_746_156# unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_3/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_3/li_n384_n810# unitcell_nbr_3/li_n176_n810# unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_3/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_4 unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_4/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_4/m1_746_156# unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_4/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_4/li_n384_n810# unitcell_nbr_4/li_n176_n810# unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_4/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_5 unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_5/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_5/m1_746_156# unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_5/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_5/li_n384_n810# unitcell_nbr_5/li_n176_n810# unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_5/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_cut_0 unitcell_nbr_cut_0/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_cut_0/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_cut_0/li_n176_n810#
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_4/A unitcell_nbr_cut_0/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_cut_0/m1_746_156# sky130_fd_sc_hd__inv_16_3/VPB unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y unitcell_nbr_cut_0/li_n384_n810#
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_5/X VSUBS unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_5/A
+ unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_5/a_27_47# unitcell_nbr_cut
Xunitcell_nbr_6 unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_6/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_6/m1_746_156# unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_6/li_n384_n810# unitcell_nbr_6/li_n176_n810# unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_6/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_cut_1 unitcell_nbr_cut_1/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_cut_1/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_cut_1/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_cut_1/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_cut_1/li_n176_n810#
+ unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_5/B unitcell_nbr_cut_1/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_cut_1/m1_746_156# sky130_fd_sc_hd__inv_16_3/VPB unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/A
+ unitcell_nbr_cut_1/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y unitcell_nbr_cut_1/li_n384_n810#
+ unitcell_nbr_cut_1/sky130_fd_sc_hd__buf_1_5/X VSUBS unitcell_nbr_6/sky130_fd_sc_hd__nor2_1_4/B
+ unitcell_nbr_cut_1/sky130_fd_sc_hd__buf_1_5/a_27_47# unitcell_nbr_cut
Xunitcell_nbr_7 unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_7/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_7/m1_746_156# unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_7/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_7/li_n384_n810# unitcell_nbr_7/li_n176_n810# unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_7/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_8 unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_8/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_8/m1_746_156# unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_8/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_8/li_n384_n810# unitcell_nbr_8/li_n176_n810# unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_8/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_9 unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_9/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_9/m1_746_156# unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_9/sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell_nbr_9/li_n384_n810# unitcell_nbr_9/li_n176_n810# unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/X
+ VSUBS unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_9/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_1/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_1/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16_3/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
.ends

.subckt NBR32 C[31] C[30] C[29] C[28] C[27] C[26] C[25] C[24] C[23] C[22] C[21] C[20]
+ C[19] C[18] C[17] C[16] C[15] C[14] C[13] C[12] C[11] C[10] C[9] C[8] C[7] C[6]
+ C[5] C[4] C[3] C[2] C[1] C[0] RESET OUT VDD VSS
Xnbrhalf_32_0 C[5] C[2] C[11] unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/B nbrhalf_32_0/unitcell_nbr_cut_0/sky130_fd_sc_hd__buf_1_5/X
+ C[8] C[14] C[4] C[13] nbrhalf_32_0/unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_4/B nbrhalf_32_0/unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_5/B
+ C[1] VSS C[10] invcell_0/sky130_fd_sc_hd__inv_16_2/Y C[7] nbrhalf_32_0/sky130_fd_sc_hd__inv_16_3/Y
+ C[3] C[6] C[12] VDD C[0] invcell_0/sky130_fd_sc_hd__inv_16_3/Y unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/B
+ C[9] VSS VSS nbrhalf_32
Xnbrhalf_32_1 C[22] C[19] C[28] nbrhalf_32_0/unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_5/B
+ OUT C[25] C[31] C[21] C[30] unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/A
+ C[18] VSS C[27] invcell_0/sky130_fd_sc_hd__inv_16_3/Y C[24] nbrhalf_32_1/sky130_fd_sc_hd__inv_16_3/Y
+ C[20] C[23] C[29] VDD C[17] invcell_0/sky130_fd_sc_hd__inv_16_2/Y nbrhalf_32_0/unitcell_nbr_12/sky130_fd_sc_hd__nor2_1_4/B
+ C[26] VSS VSS nbrhalf_32
Xunitcell_nbr_0 unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/B
+ unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_0/m1_746_156# unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/B unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_0/sky130_fd_sc_hd__nor2_1_4/Y nbrhalf_32_1/sky130_fd_sc_hd__inv_16_3/Y
+ VDD C[15] unitcell_nbr_0/li_n176_n810# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/X
+ VSS unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xunitcell_nbr_1 unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_4/a_109_297# unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/X unitcell_nbr_0/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/a_27_47# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_4/A
+ unitcell_nbr_1/m1_746_156# unitcell_nbr_0/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_5/Y
+ unitcell_nbr_1/sky130_fd_sc_hd__nor2_1_4/Y nbrhalf_32_1/sky130_fd_sc_hd__inv_16_3/Y
+ VDD C[16] unitcell_nbr_1/li_n176_n810# unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/X
+ VSS unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/A unitcell_nbr_1/sky130_fd_sc_hd__buf_1_5/a_27_47#
+ unitcell_nbr
Xinvcell_0 VSS invcell_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD RESET invcell_0/sky130_fd_sc_hd__inv_16_2/Y
+ VSS invcell
.ends

.subckt brbufhalf_128 unitcell2bufcut_1/li_n460_n386# unitcell2buf_7/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/A unitcell2buf_2/li_n460_n386# unitcell2buf_11/m2_136_462#
+ sky130_fd_sc_hd__inv_16_2/VGND unitcell2buf_10/li_n460_n386# unitcell2buf_5/li_n460_n386#
+ unitcell2buf_8/li_n460_n386# unitcell2buf_0/li_n460_n386# sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_3/VGND unitcell2buf_3/li_n460_n386# unitcell2buf_11/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16_0/VGND unitcell2buf_6/li_n460_n386#
+ unitcell2bufcut_0/li_n460_n386# unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_9/li_n460_n386#
+ unitcell2buf_1/li_n460_n386# unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_1/VGND
+ VSUBS unitcell2buf_12/li_n460_n386#
Xunitcell2buf_1 unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_1/li_n460_n386# unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_1/li_80_172# unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_1/a_24_n198#
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16_3/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_2 unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_2/li_n460_n386# unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_2/li_80_172# unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_2/a_24_n198#
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_3 unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_3/li_n460_n386# unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_3/li_80_172# unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_3/a_24_n198#
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_4 unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_4/li_n460_n386# unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_4/li_80_172# unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_4/a_24_n198#
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_5 unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_5/li_n460_n386# unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_5/li_80_172# unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_5/a_24_n198#
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_6 unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_6/li_n460_n386# unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_6/li_80_172# unitcell2bufcut_1/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_6/a_24_n198#
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_7 unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_7/li_n460_n386# unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_7/li_80_172# unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_7/a_24_n198#
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_8 unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_8/li_n460_n386# unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_8/li_80_172# unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_8/a_24_n198#
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_9 unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_9/li_n460_n386# unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_9/li_80_172# unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_9/a_24_n198#
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_10 unitcell2buf_10/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_10/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_10/li_n460_n386# unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_10/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_10/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_10/li_80_172# unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_10/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_10/a_24_n198#
+ unitcell2buf_10/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_11 unitcell2buf_11/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_11/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_11/li_n460_n386# unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_11/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_11/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_11/li_80_172# unitcell2buf_11/m2_136_462# sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_11/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_11/a_24_n198#
+ unitcell2buf_11/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2buf_12 unitcell2buf_12/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_12/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_12/li_n460_n386# unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_12/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_12/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_12/li_80_172# unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_12/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_12/a_24_n198#
+ unitcell2buf_12/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xunitcell2bufcut_0 unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_2/B unitcell2bufcut_0/a_24_n198# unitcell2bufcut_0/li_n460_n386#
+ unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2bufcut_0/li_80_172# sky130_fd_sc_hd__inv_16_3/VPB unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/X
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_3/B VSUBS
+ unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_0/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2bufcut_1 unitcell2bufcut_1/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2bufcut_1/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2bufcut_1/sky130_fd_sc_hd__nor2_1_2/B unitcell2bufcut_1/a_24_n198# unitcell2bufcut_1/li_n460_n386#
+ unitcell2bufcut_1/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2bufcut_1/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2bufcut_1/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2bufcut_1/li_80_172# sky130_fd_sc_hd__inv_16_3/VPB unitcell2bufcut_1/sky130_fd_sc_hd__buf_1_1/X
+ sky130_fd_sc_hd__inv_16_3/Y unitcell2bufcut_1/sky130_fd_sc_hd__nor2_1_3/B VSUBS
+ unitcell2bufcut_1/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_1/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_0 unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_0/li_n460_n386# unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_0/li_80_172# unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_0/a_24_n198#
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16_2/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
.ends

.subckt BR128half_bottom brbufhalf_128_0/unitcell2bufcut_0/li_n460_n386# brbufhalf_2/unitcell2buf_4/li_n460_n386#
+ brbufhalf_0/unitcell2bufcut_3/li_n460_n386# brbufhalf_128_0/unitcell2buf_4/li_n460_n386#
+ brbufhalf_2/unitcell2buf_26/m2_136_462# brbufhalf_0/unitcell2buf_3/li_n460_n386#
+ brbufhalf_1/unitcell2buf_9/li_n460_n386# brbufhalf_2/unitcell2buf_26/li_n460_n386#
+ brbufhalf_2/unitcell2bufcut_2/li_n460_n386# brbufhalf_1/unitcell2buf_1/li_n460_n386#
+ brbufhalf_0/unitcell2buf_24/li_n460_n386# brbufhalf_2/unitcell2buf_7/li_n460_n386#
+ brbufhalf_128_0/unitcell2buf_7/li_n460_n386# brbufhalf_128_0/unitcell2buf_11/li_n460_n386#
+ brbufhalf_0/unitcell2buf_6/li_n460_n386# brbufhalf_0/unitcell2buf_27/li_n460_n386#
+ brbufhalf_1/unitcell2buf_4/li_n460_n386# brbufhalf_1/unitcell2buf_24/li_n460_n386#
+ brbufhalf_1/unitcell2bufcut_3/li_n460_n386# sky130_fd_sc_hd__inv_16_3/A brbufhalf_2/unitcell2buf_2/li_n460_n386#
+ brbufhalf_0/unitcell2buf_9/li_n460_n386# brbufhalf_128_0/unitcell2buf_11/m2_136_462#
+ brbufhalf_128_0/unitcell2buf_2/li_n460_n386# brbufhalf_0/unitcell2buf_1/li_n460_n386#
+ brbufhalf_1/unitcell2buf_7/li_n460_n386# brbufhalf_1/unitcell2buf_27/li_n460_n386#
+ brbufhalf_128_0/unitcell2bufcut_1/li_n460_n386# brbufhalf_2/unitcell2buf_24/li_n460_n386#
+ brbufhalf_2/unitcell2buf_5/li_n460_n386# brbufhalf_128_0/unitcell2buf_5/li_n460_n386#
+ brbufhalf_0/unitcell2buf_4/li_n460_n386# brbufhalf_0/unitcell2buf_25/li_n460_n386#
+ brbufhalf_2/unitcell2buf_27/li_n460_n386# brbufhalf_1/unitcell2buf_2/li_n460_n386#
+ brbufhalf_2/unitcell2bufcut_3/li_n460_n386# brbufhalf_2/unitcell2buf_8/li_n460_n386#
+ brbufhalf_128_0/unitcell2buf_8/li_n460_n386# brbufhalf_2/unitcell2buf_0/li_n460_n386#
+ brbufhalf_128_0/unitcell2buf_12/li_n460_n386# brbufhalf_0/unitcell2buf_7/li_n460_n386#
+ brbufhalf_128_0/unitcell2buf_0/li_n460_n386# brbufhalf_1/unitcell2buf_5/li_n460_n386#
+ brbufhalf_1/unitcell2buf_25/li_n460_n386# brbufhalf_2/unitcell2buf_3/li_n460_n386#
+ brbufhalf_0/unitcell2bufcut_2/li_n460_n386# brbufhalf_128_0/unitcell2buf_3/li_n460_n386#
+ brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A brbufhalf_0/unitcell2buf_2/li_n460_n386#
+ brbufhalf_1/unitcell2buf_8/li_n460_n386# brbufhalf_2/unitcell2buf_25/li_n460_n386#
+ brbufhalf_2/unitcell2buf_6/li_n460_n386# brbufhalf_1/unitcell2buf_0/li_n460_n386#
+ brbufhalf_128_0/unitcell2buf_6/li_n460_n386# brbufhalf_128_0/unitcell2buf_10/li_n460_n386#
+ brbufhalf_0/unitcell2buf_5/li_n460_n386# brbufhalf_0/unitcell2buf_26/li_n460_n386#
+ brbufhalf_1/unitcell2buf_3/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB brbufhalf_2/unitcell2buf_9/li_n460_n386#
+ brbufhalf_1/unitcell2bufcut_2/li_n460_n386# brbufhalf_128_0/unitcell2buf_9/li_n460_n386#
+ brbufhalf_2/unitcell2buf_1/li_n460_n386# brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_0/unitcell2buf_8/li_n460_n386# brbufhalf_128_0/unitcell2buf_1/li_n460_n386#
+ brbufhalf_0/unitcell2buf_0/li_n460_n386# brbufhalf_1/unitcell2buf_6/li_n460_n386#
+ VSUBS brbufhalf_1/unitcell2buf_26/li_n460_n386#
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xbrbufhalf_0 brbufhalf_0/unitcell2buf_7/li_n460_n386# brbufhalf_0/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_1/Y brbufhalf_0/unitcell2buf_2/li_n460_n386# brbufhalf_0/unitcell2buf_24/li_n460_n386#
+ VSUBS brbufhalf_0/unitcell2buf_5/li_n460_n386# brbufhalf_0/unitcell2buf_27/li_n460_n386#
+ brbufhalf_0/unitcell2buf_8/li_n460_n386# brbufhalf_0/unitcell2buf_0/li_n460_n386#
+ brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X brbufhalf_0/unitcell2buf_3/li_n460_n386#
+ VSUBS brbufhalf_0/unitcell2buf_25/li_n460_n386# brbufhalf_0/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_0/unitcell2buf_6/li_n460_n386# VSUBS brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_0/sky130_fd_sc_hd__inv_16_7/Y brbufhalf_0/unitcell2buf_9/li_n460_n386#
+ brbufhalf_0/unitcell2buf_1/li_n460_n386# brbufhalf_0/sky130_fd_sc_hd__inv_16_5/Y
+ brbufhalf_0/unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_1/Y brbufhalf_128_0/unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS VSUBS brbufhalf_0/unitcell2buf_26/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ brbufhalf
Xbrbufhalf_1 brbufhalf_1/unitcell2buf_7/li_n460_n386# brbufhalf_1/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/Y brbufhalf_1/unitcell2buf_2/li_n460_n386# brbufhalf_1/unitcell2buf_24/li_n460_n386#
+ VSUBS brbufhalf_1/unitcell2buf_5/li_n460_n386# brbufhalf_1/unitcell2buf_27/li_n460_n386#
+ brbufhalf_1/unitcell2buf_8/li_n460_n386# brbufhalf_1/unitcell2buf_0/li_n460_n386#
+ brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X brbufhalf_1/unitcell2buf_3/li_n460_n386#
+ VSUBS brbufhalf_1/unitcell2buf_25/li_n460_n386# brbufhalf_1/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_1/unitcell2buf_6/li_n460_n386# VSUBS brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_1/sky130_fd_sc_hd__inv_16_7/Y brbufhalf_1/unitcell2buf_9/li_n460_n386#
+ brbufhalf_1/unitcell2buf_1/li_n460_n386# brbufhalf_1/sky130_fd_sc_hd__inv_16_5/Y
+ brbufhalf_1/unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_3/Y brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS VSUBS brbufhalf_1/unitcell2buf_26/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ brbufhalf
Xbrbufhalf_2 brbufhalf_2/unitcell2buf_7/li_n460_n386# brbufhalf_2/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_1/Y brbufhalf_2/unitcell2buf_2/li_n460_n386# brbufhalf_2/unitcell2buf_24/li_n460_n386#
+ VSUBS brbufhalf_2/unitcell2buf_5/li_n460_n386# brbufhalf_2/unitcell2buf_27/li_n460_n386#
+ brbufhalf_2/unitcell2buf_8/li_n460_n386# brbufhalf_2/unitcell2buf_0/li_n460_n386#
+ brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X brbufhalf_2/unitcell2buf_3/li_n460_n386#
+ VSUBS brbufhalf_2/unitcell2buf_25/li_n460_n386# brbufhalf_2/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_2/unitcell2buf_6/li_n460_n386# VSUBS brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_2/sky130_fd_sc_hd__inv_16_7/Y brbufhalf_2/unitcell2buf_9/li_n460_n386#
+ brbufhalf_2/unitcell2buf_1/li_n460_n386# brbufhalf_2/sky130_fd_sc_hd__inv_16_5/Y
+ brbufhalf_2/unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_1/Y brbufhalf_2/unitcell2buf_26/m2_136_462#
+ VSUBS VSUBS brbufhalf_2/unitcell2buf_26/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ brbufhalf
Xbrbufhalf_128_0 brbufhalf_128_0/unitcell2bufcut_1/li_n460_n386# brbufhalf_128_0/unitcell2buf_7/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/Y brbufhalf_128_0/unitcell2buf_2/li_n460_n386# brbufhalf_128_0/unitcell2buf_11/m2_136_462#
+ VSUBS brbufhalf_128_0/unitcell2buf_10/li_n460_n386# brbufhalf_128_0/unitcell2buf_5/li_n460_n386#
+ brbufhalf_128_0/unitcell2buf_8/li_n460_n386# brbufhalf_128_0/unitcell2buf_0/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/Y VSUBS brbufhalf_128_0/unitcell2buf_3/li_n460_n386# brbufhalf_128_0/unitcell2buf_11/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/VPB VSUBS brbufhalf_128_0/unitcell2buf_6/li_n460_n386#
+ brbufhalf_128_0/unitcell2bufcut_0/li_n460_n386# brbufhalf_128_0/unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_128_0/unitcell2buf_9/li_n460_n386# brbufhalf_128_0/unitcell2buf_1/li_n460_n386#
+ brbufhalf_128_0/unitcell2buf_4/li_n460_n386# VSUBS VSUBS brbufhalf_128_0/unitcell2buf_12/li_n460_n386#
+ brbufhalf_128
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
.ends

.subckt BR128half brbufhalf_2/unitcell2buf_4/li_n460_n386# brbufhalf_0/unitcell2bufcut_3/li_n460_n386#
+ brbufhalf_0/unitcell2buf_3/li_n460_n386# brbufhalf_3/unitcell2buf_2/li_n460_n386#
+ brbufhalf_1/unitcell2buf_9/li_n460_n386# brbufhalf_2/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_2/unitcell2buf_26/li_n460_n386# brbufhalf_1/unitcell2buf_1/li_n460_n386#
+ brbufhalf_0/unitcell2buf_24/li_n460_n386# brbufhalf_2/unitcell2buf_7/li_n460_n386#
+ brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A brbufhalf_0/unitcell2buf_6/li_n460_n386#
+ brbufhalf_3/unitcell2buf_5/li_n460_n386# brbufhalf_1/unitcell2buf_4/li_n460_n386#
+ brbufhalf_0/unitcell2buf_27/li_n460_n386# brbufhalf_1/unitcell2buf_24/li_n460_n386#
+ brbufhalf_3/unitcell2buf_26/li_n460_n386# brbufhalf_1/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/A brbufhalf_1/unitcell2buf_26/m2_136_462# brbufhalf_2/unitcell2buf_2/li_n460_n386#
+ brbufhalf_0/unitcell2buf_9/li_n460_n386# brbufhalf_3/unitcell2buf_8/li_n460_n386#
+ brbufhalf_3/unitcell2buf_0/li_n460_n386# brbufhalf_0/unitcell2buf_1/li_n460_n386#
+ brbufhalf_3/unitcell2bufcut_2/li_n460_n386# brbufhalf_1/unitcell2buf_7/li_n460_n386#
+ brbufhalf_1/unitcell2buf_27/li_n460_n386# brbufhalf_2/unitcell2buf_24/li_n460_n386#
+ brbufhalf_2/unitcell2buf_5/li_n460_n386# brbufhalf_0/unitcell2buf_4/li_n460_n386#
+ brbufhalf_3/unitcell2buf_3/li_n460_n386# brbufhalf_2/unitcell2bufcut_3/li_n460_n386#
+ brbufhalf_2/unitcell2buf_27/li_n460_n386# brbufhalf_0/unitcell2buf_25/li_n460_n386#
+ brbufhalf_1/unitcell2buf_2/li_n460_n386# brbufhalf_2/unitcell2buf_8/li_n460_n386#
+ brbufhalf_3/unitcell2buf_24/li_n460_n386# brbufhalf_2/unitcell2buf_0/li_n460_n386#
+ brbufhalf_3/unitcell2buf_6/li_n460_n386# brbufhalf_0/unitcell2buf_7/li_n460_n386#
+ brbufhalf_1/unitcell2buf_5/li_n460_n386# brbufhalf_3/unitcell2buf_27/li_n460_n386#
+ brbufhalf_1/unitcell2buf_25/li_n460_n386# brbufhalf_3/unitcell2buf_9/li_n460_n386#
+ brbufhalf_2/unitcell2buf_3/li_n460_n386# brbufhalf_0/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A brbufhalf_0/unitcell2buf_2/li_n460_n386#
+ brbufhalf_3/unitcell2buf_1/li_n460_n386# brbufhalf_1/unitcell2buf_8/li_n460_n386#
+ brbufhalf_3/unitcell2bufcut_3/li_n460_n386# brbufhalf_2/unitcell2buf_25/li_n460_n386#
+ brbufhalf_2/unitcell2buf_6/li_n460_n386# brbufhalf_1/unitcell2buf_0/li_n460_n386#
+ brbufhalf_0/unitcell2buf_5/li_n460_n386# brbufhalf_3/unitcell2buf_4/li_n460_n386#
+ brbufhalf_2/sky130_fd_sc_hd__inv_16_5/Y brbufhalf_3/unitcell2buf_26/m2_136_462#
+ brbufhalf_0/unitcell2buf_26/li_n460_n386# brbufhalf_1/unitcell2buf_3/li_n460_n386#
+ brbufhalf_2/unitcell2buf_9/li_n460_n386# brbufhalf_3/unitcell2buf_25/li_n460_n386#
+ brbufhalf_1/unitcell2bufcut_2/li_n460_n386# brbufhalf_2/unitcell2buf_1/li_n460_n386#
+ brbufhalf_3/unitcell2buf_7/li_n460_n386# brbufhalf_0/unitcell2buf_8/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/VPB brbufhalf_0/unitcell2buf_0/li_n460_n386# brbufhalf_1/unitcell2buf_6/li_n460_n386#
+ VSUBS brbufhalf_1/unitcell2buf_26/li_n460_n386#
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xbrbufhalf_0 brbufhalf_0/unitcell2buf_7/li_n460_n386# brbufhalf_0/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_1/Y brbufhalf_0/unitcell2buf_2/li_n460_n386# brbufhalf_0/unitcell2buf_24/li_n460_n386#
+ VSUBS brbufhalf_0/unitcell2buf_5/li_n460_n386# brbufhalf_0/unitcell2buf_27/li_n460_n386#
+ brbufhalf_0/unitcell2buf_8/li_n460_n386# brbufhalf_0/unitcell2buf_0/li_n460_n386#
+ brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X brbufhalf_0/unitcell2buf_3/li_n460_n386#
+ VSUBS brbufhalf_0/unitcell2buf_25/li_n460_n386# brbufhalf_0/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_0/unitcell2buf_6/li_n460_n386# VSUBS brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_0/sky130_fd_sc_hd__inv_16_7/Y brbufhalf_0/unitcell2buf_9/li_n460_n386#
+ brbufhalf_0/unitcell2buf_1/li_n460_n386# brbufhalf_0/sky130_fd_sc_hd__inv_16_5/Y
+ brbufhalf_0/unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_1/Y brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS VSUBS brbufhalf_0/unitcell2buf_26/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ brbufhalf
Xbrbufhalf_1 brbufhalf_1/unitcell2buf_7/li_n460_n386# brbufhalf_1/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/Y brbufhalf_1/unitcell2buf_2/li_n460_n386# brbufhalf_1/unitcell2buf_24/li_n460_n386#
+ VSUBS brbufhalf_1/unitcell2buf_5/li_n460_n386# brbufhalf_1/unitcell2buf_27/li_n460_n386#
+ brbufhalf_1/unitcell2buf_8/li_n460_n386# brbufhalf_1/unitcell2buf_0/li_n460_n386#
+ brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X brbufhalf_1/unitcell2buf_3/li_n460_n386#
+ VSUBS brbufhalf_1/unitcell2buf_25/li_n460_n386# brbufhalf_1/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_1/unitcell2buf_6/li_n460_n386# VSUBS brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_1/sky130_fd_sc_hd__inv_16_7/Y brbufhalf_1/unitcell2buf_9/li_n460_n386#
+ brbufhalf_1/unitcell2buf_1/li_n460_n386# brbufhalf_1/sky130_fd_sc_hd__inv_16_5/Y
+ brbufhalf_1/unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_3/Y brbufhalf_1/unitcell2buf_26/m2_136_462#
+ VSUBS VSUBS brbufhalf_1/unitcell2buf_26/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ brbufhalf
Xbrbufhalf_2 brbufhalf_2/unitcell2buf_7/li_n460_n386# brbufhalf_2/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/Y brbufhalf_2/unitcell2buf_2/li_n460_n386# brbufhalf_2/unitcell2buf_24/li_n460_n386#
+ VSUBS brbufhalf_2/unitcell2buf_5/li_n460_n386# brbufhalf_2/unitcell2buf_27/li_n460_n386#
+ brbufhalf_2/unitcell2buf_8/li_n460_n386# brbufhalf_2/unitcell2buf_0/li_n460_n386#
+ brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X brbufhalf_2/unitcell2buf_3/li_n460_n386#
+ VSUBS brbufhalf_2/unitcell2buf_25/li_n460_n386# brbufhalf_2/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_2/unitcell2buf_6/li_n460_n386# VSUBS brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_2/sky130_fd_sc_hd__inv_16_7/Y brbufhalf_2/unitcell2buf_9/li_n460_n386#
+ brbufhalf_2/unitcell2buf_1/li_n460_n386# brbufhalf_2/sky130_fd_sc_hd__inv_16_5/Y
+ brbufhalf_2/unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_3/Y brbufhalf_3/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS VSUBS brbufhalf_2/unitcell2buf_26/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ brbufhalf
Xbrbufhalf_3 brbufhalf_3/unitcell2buf_7/li_n460_n386# brbufhalf_3/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_1/Y brbufhalf_3/unitcell2buf_2/li_n460_n386# brbufhalf_3/unitcell2buf_24/li_n460_n386#
+ VSUBS brbufhalf_3/unitcell2buf_5/li_n460_n386# brbufhalf_3/unitcell2buf_27/li_n460_n386#
+ brbufhalf_3/unitcell2buf_8/li_n460_n386# brbufhalf_3/unitcell2buf_0/li_n460_n386#
+ brbufhalf_3/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X brbufhalf_3/unitcell2buf_3/li_n460_n386#
+ VSUBS brbufhalf_3/unitcell2buf_25/li_n460_n386# brbufhalf_3/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_3/unitcell2buf_6/li_n460_n386# VSUBS brbufhalf_3/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_3/sky130_fd_sc_hd__inv_16_7/Y brbufhalf_3/unitcell2buf_9/li_n460_n386#
+ brbufhalf_3/unitcell2buf_1/li_n460_n386# brbufhalf_3/sky130_fd_sc_hd__inv_16_5/Y
+ brbufhalf_3/unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_1/Y brbufhalf_3/unitcell2buf_26/m2_136_462#
+ VSUBS VSUBS brbufhalf_3/unitcell2buf_26/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ brbufhalf
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
.ends

.subckt BR128 RESET VDD C[0] C[1] C[2] C[3] C[4] C[5] C[7] C[8] C[9] C[10] C[11] C[12]
+ C[13] C[14] C[15] C[16] C[17] C[18] C[19] C[20] C[21] C[22] C[23] C[24] C[25] C[26]
+ C[27] C[28] C[29] C[30] C[6] C[31] C[32] C[33] C[34] C[35] C[36] C[37] C[38] C[39]
+ C[40] C[41] C[42] C[43] C[44] C[45] C[46] C[47] C[48] C[49] C[50] C[51] C[52] C[53]
+ C[54] C[55] C[56] C[57] C[58] C[59] C[60] C[61] C[62] C[95] C[96] C[97] C[98] C[99]
+ C[100] C[101] C[102] C[103] C[104] C[105] C[106] C[107] C[108] C[109] C[110] C[111]
+ C[112] C[113] C[114] C[115] C[116] C[117] C[118] C[119] C[120] C[121] C[122] C[123]
+ C[124] C[125] C[126] C[127] C[63] C[64] C[65] C[66] C[67] C[68] C[69] C[70] C[71]
+ C[72] C[73] C[74] C[75] C[76] C[77] C[78] C[79] C[80] C[81] C[82] C[83] C[84] C[85]
+ C[86] C[87] C[88] C[89] C[90] C[91] C[92] C[93] C[94] OUT VSS
XBR128half_bottom_0 C[46] C[73] C[54] C[41] BR128half_bottom_0/brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ C[58] C[83] C[63] C[78] C[92] C[50] C[69] C[37] C[32] C[55] C[48] C[89] C[82] C[86]
+ sky130_fd_sc_hd__inv_16_1/Y C[75] C[51] BR128half_0/brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ C[43] C[60] C[85] C[80] C[38] C[66] C[72] C[40] C[57] C[49] C[64] C[91] C[70] C[68]
+ C[36] C[77] C[33] C[53] C[45] C[88] C[81] C[74] C[62] C[42] BR128half_bottom_0/brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ C[59] C[84] C[65] C[71] C[93] C[39] C[34] C[56] C[47] C[90] VDD C[67] C[94] C[35]
+ C[76] BR128half_bottom_0/brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ C[52] C[44] C[61] C[87] VSS C[79] BR128half_bottom
Xsky130_fd_sc_hd__inv_8_0 sky130_fd_sc_hd__inv_8_0/A sky130_fd_sc_hd__inv_8_0/Y VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__buf_2_0 VDD VSS sky130_fd_sc_hd__inv_8_0/A RESET VSS VDD sky130_fd_sc_hd__buf_2
XBR128half_0 C[121] C[23] C[27] C[107] C[4] C[126] C[111] C[13] C[19] C[117] BR128half_0/brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ C[24] C[104] C[10] C[17] C[3] C[95] C[7] sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ C[123] C[20] C[100] C[109] C[29] C[110] C[6] C[1] C[114] C[120] C[26] C[106] C[118]
+ C[112] C[18] C[12] C[116] C[98] C[125] C[103] C[22] C[9] C[96] C[2] C[99] C[122]
+ C[31] BR128half_0/brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A C[28]
+ C[108] C[5] C[102] C[113] C[119] C[14] C[25] C[105] unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/A
+ BR128half_bottom_0/brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A C[16]
+ C[11] C[115] C[97] C[15] C[124] C[101] C[21] VDD C[30] C[8] VSS C[0] BR128half
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_8_0/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_8_0/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xunitcell2buf_0 unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/a_109_297#
+ OUT C[127] unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_0/li_80_172# BR128half_0/brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ VDD unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/A
+ unitcell2buf_0/a_24_n198# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/B unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ VSS unitcell2buf
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=5.36e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__buf_12 A X VGND VPWR VNB VPB
X0 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__nand2b_1 Y A_N B VGND VPWR VNB VPB
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__o21ai_2 B1 Y A2 A1 VGND VPWR VNB VPB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_0 VGND VPWR Y B1 A2 A1 VNB VPB
X0 a_120_369# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 Y A2 a_120_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt puf_super reset clk si rstn puf_sel1 puf_sel0 length1 length0 out so vccd1
+ vssd1
Xsky130_fd_sc_hd__decap_12_2470 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2481 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2492 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1780 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1791 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_7 vssd1 vccd1 BR128_1/C[113] BR128_0/C[113] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_7 sky130_fd_sc_hd__clkinv_4_2/A NBR32_1/C[12] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1010 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1021 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1032 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1043 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1054 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1065 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1076 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1087 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1098 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5309 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4608 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4619 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3907 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3918 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3929 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5106 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5117 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5128 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5139 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4405 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4416 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4427 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4438 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3704 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4449 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3715 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3726 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3737 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3748 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3759 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5640 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4950 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4961 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4972 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4983 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4994 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1609 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_9 sky130_fd_sc_hd__nand2_1_9/Y BR128_0/OUT sky130_fd_sc_hd__nor2_1_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_4202 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4213 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4224 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4235 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3501 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4246 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3512 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4257 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3523 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4268 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3534 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4279 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2800 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3545 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2811 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3556 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3567 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2822 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3578 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2833 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2844 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3589 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2855 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2866 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2877 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2888 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2899 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_10 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_21 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_32 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_43 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_54 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_65 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5470 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_76 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5481 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_87 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5492 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_98 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4780 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4791 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_10 vccd1 vssd1 BR128_1/C[84] sky130_fd_sc_hd__buf_6_10/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__decap_12_407 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_418 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_429 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2107 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2118 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2129 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1406 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1417 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1428 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1439 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_930 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_941 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_952 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_963 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_974 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4010 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_985 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4021 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_996 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4032 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4043 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4054 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3320 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4065 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3331 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4076 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3342 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4087 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4098 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3353 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3364 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3375 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2630 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3386 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2652 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3397 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2663 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2674 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1940 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1951 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2696 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1962 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1973 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1984 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1995 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_8_1 BR64_1/C[9] sky130_fd_sc_hd__clkbuf_8_1/A vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__decap_12_204 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_215 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_226 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_237 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_248 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_259 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1203 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1214 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1225 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1236 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1247 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1258 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1269 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_1 sky130_fd_sc_hd__clkinv_8_3/A sky130_fd_sc_hd__clkinv_8_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_760 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_771 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_782 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_793 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3150 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3161 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3172 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3183 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3194 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2460 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2471 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2482 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2493 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1770 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1781 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1792 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_8 vssd1 vccd1 BR128_1/C[123] BR128_0/C[123] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_8 sky130_fd_sc_hd__clkinv_4_3/A BR32_0/C[5] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1000 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1011 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1022 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1033 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1044 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1055 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1066 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1077 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1088 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1099 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_590 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2290 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4609 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3908 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3919 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5107 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5118 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5129 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4406 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4417 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4428 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4439 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3705 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3716 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3727 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3738 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3749 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5630 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4940 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4951 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4962 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4973 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4984 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4995 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4203 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4214 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4225 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4236 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3502 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4247 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4258 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3513 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3524 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4269 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3535 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2801 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3546 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2812 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2823 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3568 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2834 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3579 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2845 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2856 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2867 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2878 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2889 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_11 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_22 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_33 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_44 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_55 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5460 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_66 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5471 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_77 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5482 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_88 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5493 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_99 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4770 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4781 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4792 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_408 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_419 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2108 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2119 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1407 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1418 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1429 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_920 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_931 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_942 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_953 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_964 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4000 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_975 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4011 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_986 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4022 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_997 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4033 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4044 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3310 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4055 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3321 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4066 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4077 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3332 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3343 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4088 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3354 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4099 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2620 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3365 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2631 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3376 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2642 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3387 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2653 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3398 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2664 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1930 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2675 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1941 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2686 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1952 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1963 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1974 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1985 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1996 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5290 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_8_2 BR64_1/C[7] sky130_fd_sc_hd__clkbuf_8_2/A vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__decap_12_205 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_216 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_227 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_238 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_249 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1204 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1215 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1226 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1237 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1248 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1259 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_2 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__clkinv_8_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_750 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_761 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_772 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_783 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_794 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3140 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3151 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3162 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3173 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3184 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2450 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3195 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2461 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2472 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2483 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2494 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1760 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1771 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1782 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1793 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_9 vssd1 vccd1 BR128_1/C[121] BR128_0/C[121] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_9 sky130_fd_sc_hd__clkinv_4_4/A BR32_0/C[3] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1001 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1012 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1023 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1034 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1045 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1056 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1067 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1078 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1089 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_580 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_591 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2280 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2291 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1590 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3909 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5108 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5119 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4407 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4418 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4429 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3706 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3717 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3728 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3739 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_10 sky130_fd_sc_hd__clkinv_4_5/A sky130_fd_sc_hd__dfrtp_2_125/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_5620 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5631 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4930 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4941 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4952 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4963 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4974 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4985 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4996 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4204 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4215 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4226 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4237 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3503 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4248 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3514 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4259 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3525 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3536 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2802 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3547 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2813 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3558 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3569 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2824 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2835 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2846 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2857 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2868 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2879 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_12 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_23 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_34 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_45 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5450 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_56 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5461 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_67 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5472 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_78 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5483 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_89 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5494 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4760 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4771 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4782 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4793 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_409 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2109 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1408 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1419 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_910 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_921 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_932 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_943 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_954 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_965 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4001 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_976 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4012 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_987 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4023 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_998 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4034 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3300 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4045 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3311 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4056 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3322 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4067 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3333 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4078 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3344 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4089 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2610 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3355 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2621 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3366 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2632 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3377 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2643 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3388 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2654 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3399 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1920 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2665 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1931 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2676 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1942 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2687 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1953 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2698 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1964 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1975 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1986 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1997 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5280 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5291 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4590 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_8_3 BR64_1/C[6] sky130_fd_sc_hd__clkbuf_8_3/A vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__decap_12_206 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_217 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_228 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_239 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_90 NBR64_0/C[37] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[36]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1205 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1216 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1227 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1238 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1249 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_3 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__clkinv_8_3/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_740 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_751 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_762 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_773 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_784 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_795 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3130 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3141 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3152 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3163 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3174 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3185 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2440 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3196 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2451 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2462 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2473 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2484 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1750 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2495 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1761 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1772 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1783 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1794 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1002 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1013 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1024 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1035 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1046 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1057 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1068 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1079 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_570 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_581 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_592 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2270 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2281 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2292 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1580 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1591 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5109 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4408 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4419 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3707 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3718 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3729 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5610 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5621 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5632 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4920 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4931 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4942 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4953 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4964 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4975 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4986 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4997 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4205 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4216 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4227 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4238 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4249 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3504 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3515 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3526 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3537 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2803 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3548 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2814 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3559 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2825 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2836 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2847 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2858 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2869 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_13 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_24 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_35 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5440 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_46 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5451 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_57 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5462 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_68 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5473 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_79 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5484 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4750 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5495 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4761 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4772 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4783 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4794 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1409 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_900 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_911 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_922 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_933 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_944 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_955 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_966 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4002 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_977 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4013 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_988 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4024 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_999 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4035 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3301 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4046 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3312 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4057 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3323 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4068 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3334 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4079 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2600 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3345 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2611 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3356 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2622 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3367 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2633 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3378 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2644 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3389 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1910 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2655 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1921 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2666 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1932 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2677 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1943 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2688 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1954 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2699 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1965 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1976 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1987 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1998 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5270 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5281 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5292 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4580 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4591 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3890 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_8_4 BR64_1/C[4] sky130_fd_sc_hd__clkbuf_8_4/A vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__decap_12_207 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_218 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_229 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_80 NBR64_1/C[47] sky130_fd_sc_hd__clkbuf_4_1/X NBR64_1/C[46]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_91 NBR64_1/C[36] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[35]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1206 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1217 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1228 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1239 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_4 sky130_fd_sc_hd__clkinv_8_7/A sky130_fd_sc_hd__clkinv_8_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_730 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_741 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_752 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_763 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_774 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_785 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_796 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3120 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3131 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3142 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3153 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3164 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2430 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3175 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2441 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3186 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2452 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3197 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2463 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2474 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1740 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2485 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1751 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2496 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1762 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1773 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1784 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1795 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1003 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1014 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1025 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1036 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1047 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1058 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1069 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_560 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_571 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_582 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_593 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2260 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2271 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2282 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2293 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1570 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1581 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1592 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_390 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2090 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4409 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3708 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3719 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5600 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5611 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5622 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5633 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4910 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4921 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4932 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4943 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4954 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4965 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4976 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4987 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4998 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4206 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4217 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4228 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4239 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3505 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3516 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3527 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3538 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2804 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3549 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2815 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2826 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2837 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2848 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2859 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_14 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_25 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5430 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_36 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5441 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_47 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5452 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_58 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5463 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_69 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5474 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4740 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5485 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4751 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5496 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4762 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4773 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4784 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4795 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_901 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_912 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_923 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_934 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_945 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_956 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_967 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4003 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_978 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4014 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_989 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4025 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4036 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3302 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4047 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3313 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4058 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3324 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4069 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3335 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3346 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2612 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3357 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3368 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2623 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2634 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3379 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1900 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1911 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2656 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1922 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2667 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1933 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2678 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1944 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2689 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1955 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1966 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1977 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1988 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1999 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5260 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5271 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5282 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5293 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4570 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4581 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4592 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3880 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3891 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_8_5 BR64_1/C[13] NBR32_1/C[13] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__decap_12_208 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_219 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_70 NBR64_1/C[57] sky130_fd_sc_hd__clkbuf_4_1/X NBR64_1/C[56]
+ sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_81 NBR64_1/C[46] sky130_fd_sc_hd__clkbuf_4_1/A NBR64_1/C[45]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_92 NBR64_1/C[35] sky130_fd_sc_hd__clkbuf_4_1/A NBR64_1/C[34]
+ sky130_fd_sc_hd__clkinv_8_5/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1207 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1218 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1229 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_5 sky130_fd_sc_hd__clkinv_8_5/Y sky130_fd_sc_hd__clkinv_8_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_720 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_731 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_742 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_753 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_764 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_775 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_786 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_797 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3110 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3121 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3132 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3143 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3154 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2420 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3165 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3176 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2431 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3187 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2442 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2453 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3198 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2464 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1730 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2475 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1741 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2486 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1752 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2497 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1763 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1774 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1785 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1796 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5090 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1004 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1015 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1026 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1037 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1048 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1059 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_550 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_561 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_572 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_583 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_594 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2250 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2261 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2272 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2283 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2294 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1560 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1571 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1582 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1593 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_380 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_391 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2080 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2091 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1390 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3709 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5612 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5623 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5634 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4900 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4911 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4922 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4933 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4944 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4955 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4966 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4977 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4988 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4999 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4207 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4218 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4229 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3506 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3517 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3528 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3539 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2805 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2816 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2827 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2838 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2849 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_15 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5420 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_26 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5431 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_37 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5442 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_48 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5453 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_59 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5464 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4730 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5475 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4741 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5486 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4752 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5497 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4763 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4774 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4785 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4796 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2_1_0 reset sky130_fd_sc_hd__nor2_1_0/Y puf_sel1 vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_902 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_913 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_924 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_935 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_946 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_957 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_968 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4004 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_979 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4015 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4026 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4037 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3303 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4048 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3314 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4059 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3325 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3336 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2602 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3347 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3358 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2624 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3369 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2635 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1901 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2646 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1912 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1923 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2668 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1934 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2679 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1945 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1956 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1967 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1978 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1989 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5250 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5261 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5272 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5283 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5294 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4560 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4571 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4582 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4593 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3870 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3881 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3892 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_60 BR128_0/C[67] sky130_fd_sc_hd__clkbuf_4_1/X BR128_0/C[66]
+ sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_71 NBR64_1/C[56] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[55]
+ sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_82 NBR64_1/C[45] sky130_fd_sc_hd__clkbuf_4_1/A NBR64_1/C[44]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_93 NBR64_1/C[34] sky130_fd_sc_hd__clkbuf_4_1/A NBR64_1/C[33]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1208 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1219 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_6 sky130_fd_sc_hd__clkinv_8_6/Y sky130_fd_sc_hd__clkinv_8_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_710 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_721 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_732 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_743 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_754 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_765 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_776 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_787 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_798 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3100 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3111 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3122 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3133 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3144 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2410 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3155 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2421 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3166 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2432 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3177 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2443 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3188 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2454 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3199 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1720 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2465 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1731 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2476 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1742 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2487 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1753 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2498 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1764 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1775 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1786 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1797 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5080 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5091 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4390 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1005 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1016 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1027 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1038 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1049 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_540 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_551 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_562 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_573 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_584 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_595 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2240 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2251 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2262 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2273 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2284 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2295 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1550 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1561 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1572 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1583 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1594 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_0 sky130_fd_sc_hd__clkbuf_4_1/A rstn vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_4_0 clk sky130_fd_sc_hd__clkinv_8_0/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_370 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_381 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_392 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2070 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2081 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2092 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1380 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1391 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5602 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5624 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5635 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4901 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4912 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4923 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4934 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4945 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4956 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4967 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4978 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4989 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4208 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4219 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3507 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3518 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3529 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2806 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2817 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2828 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2839 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5410 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_16 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5421 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_27 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5432 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_38 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5443 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_49 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5454 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4720 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5465 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5476 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4731 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_0 vccd1 vssd1 BR64_1/C[47] NBR64_1/C[47] vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__decap_12_4742 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5487 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4753 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5498 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4764 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4775 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4786 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4797 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_1/B sky130_fd_sc_hd__nor2_1_1/Y
+ reset vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_1/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_903 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_914 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_925 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_936 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_947 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_958 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_969 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4005 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4016 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4027 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4038 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3304 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4049 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3315 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3326 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3337 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2603 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3348 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2614 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3359 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2625 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2636 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2647 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1902 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1913 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2658 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1924 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1935 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1946 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1957 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1968 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1979 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5240 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5251 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5262 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5273 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5284 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4550 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5295 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4561 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4572 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4583 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4594 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3860 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3871 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3882 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3893 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_50 NBR128_0/C[77] sky130_fd_sc_hd__clkbuf_4_1/X NBR128_0/C[76]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_61 BR128_0/C[66] sky130_fd_sc_hd__clkbuf_4_1/X NBR128_1/C[65]
+ sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_72 NBR64_1/C[55] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[54]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_83 NBR64_1/C[44] sky130_fd_sc_hd__clkbuf_4_1/A NBR64_1/C[43]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_94 NBR64_1/C[33] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[32]
+ sky130_fd_sc_hd__clkinv_8_5/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_7 sky130_fd_sc_hd__clkinv_8_7/Y sky130_fd_sc_hd__clkinv_8_7/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_700 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_711 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_722 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_733 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_744 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_755 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_766 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_777 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_788 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_799 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3101 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3112 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3123 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3134 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2400 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3145 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2411 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3156 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3167 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2422 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3178 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2433 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2444 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3189 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1710 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2455 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1721 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2466 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1732 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2477 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1743 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2488 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1754 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2499 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1765 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1776 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1787 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1798 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5070 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5081 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5092 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4380 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4391 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3690 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1006 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1017 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1028 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1039 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_530 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_541 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_552 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_563 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_574 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_585 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_596 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2230 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2241 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2252 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2263 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2274 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1540 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2285 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1551 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2296 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1562 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1573 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1584 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1595 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_1 sky130_fd_sc_hd__clkbuf_4_1/X sky130_fd_sc_hd__clkbuf_4_1/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_4_1 sky130_fd_sc_hd__clkinv_4_1/A BR64_1/C[30] vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_360 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_371 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_382 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_393 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2060 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2071 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2082 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2093 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1370 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1381 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1392 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5603 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5614 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5625 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5636 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4902 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4913 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4924 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4935 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4946 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4957 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4968 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4979 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_190 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3508 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3519 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2807 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2818 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2829 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR64_0 BR64_0/OUT vccd1 BR64_0/RESET BR64_1/C[0] BR64_1/C[1] BR64_1/C[2] BR64_1/C[3]
+ BR64_1/C[4] BR64_1/C[5] BR64_1/C[6] BR64_1/C[7] BR64_1/C[8] BR64_1/C[9] BR64_1/C[10]
+ BR64_1/C[11] BR64_1/C[12] BR64_1/C[13] BR64_1/C[14] BR64_1/C[15] BR64_1/C[16] BR64_1/C[17]
+ BR64_1/C[18] BR64_1/C[19] BR64_1/C[20] BR64_1/C[21] BR64_1/C[22] BR64_1/C[23] BR64_1/C[24]
+ BR64_1/C[25] BR64_1/C[26] BR64_1/C[27] BR64_1/C[28] BR64_1/C[29] BR64_1/C[30] BR64_1/C[31]
+ BR64_1/C[32] BR64_1/C[33] BR64_1/C[34] BR64_1/C[35] BR64_1/C[36] BR64_1/C[37] BR64_1/C[38]
+ BR64_1/C[39] BR64_1/C[40] BR64_1/C[41] BR64_1/C[42] BR64_1/C[43] BR64_1/C[44] BR64_1/C[45]
+ BR64_1/C[46] BR64_1/C[47] BR64_1/C[48] BR64_1/C[49] BR64_1/C[50] BR64_1/C[51] BR64_1/C[52]
+ BR64_1/C[53] BR64_1/C[54] BR64_1/C[55] BR64_1/C[56] BR64_1/C[57] BR64_1/C[58] BR64_1/C[59]
+ BR64_1/C[60] BR64_1/C[61] BR64_1/C[62] BR64_1/C[63] vssd1 BR64
Xsky130_fd_sc_hd__decap_12_5400 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_17 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5411 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5422 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_28 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5433 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_39 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5444 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4710 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5455 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4721 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5466 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4732 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5477 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_1 vccd1 vssd1 BR64_1/C[28] sky130_fd_sc_hd__buf_6_1/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__decap_12_4743 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5488 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4754 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5499 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4765 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4776 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4787 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4798 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2_1_2 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__nor2_1_2/Y
+ length1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_2/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_904 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_915 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_926 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_937 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_948 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_959 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4006 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4017 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4028 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4039 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3305 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3316 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3327 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3338 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2604 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3349 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2615 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2626 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2637 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1903 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2648 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1914 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2659 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1925 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1936 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1947 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1958 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1969 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5230 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5241 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5252 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5263 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5274 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4540 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5285 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4551 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5296 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4562 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4573 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4584 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3850 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4595 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3861 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3872 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3883 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3894 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_40 NBR128_0/C[87] sky130_fd_sc_hd__clkbuf_4_1/A NBR128_0/C[86]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_51 NBR128_0/C[76] sky130_fd_sc_hd__clkbuf_4_1/X BR128_1/C[75]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_62 NBR128_1/C[65] sky130_fd_sc_hd__clkbuf_4_1/X NBR128_1/C[64]
+ sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_73 NBR64_1/C[54] sky130_fd_sc_hd__clkbuf_4_1/X NBR64_1/C[53]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_84 NBR64_1/C[43] sky130_fd_sc_hd__clkbuf_4_1/A NBR64_1/C[42]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_95 NBR64_1/C[32] sky130_fd_sc_hd__clkbuf_4_1/A NBR64_1/C[31]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkinv_8_8 sky130_fd_sc_hd__clkinv_8_9/A sky130_fd_sc_hd__clkinv_8_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_701 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_712 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_723 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_734 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_745 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_756 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_767 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_778 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_789 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3102 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3113 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3124 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3135 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3146 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2401 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2412 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3157 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2423 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3168 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2434 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3179 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1700 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2445 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1711 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2456 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1722 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2467 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2478 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1733 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1744 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2489 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1755 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1766 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1777 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1788 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_2_0 sky130_fd_sc_hd__nor2_1_2/B puf_sel0 sky130_fd_sc_hd__nor2_1_1/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__decap_12_1799 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5060 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5071 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5082 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5093 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4370 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4381 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4392 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3680 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3691 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2990 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1007 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1018 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1029 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_520 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_531 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_542 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_553 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_564 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_575 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_586 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_597 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2220 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2231 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2242 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2253 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2264 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1530 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2275 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1541 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2286 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2297 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1552 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1563 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1574 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1585 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1596 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_2 BR128_1/C[107] NBR128_0/C[107] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_4_2 sky130_fd_sc_hd__clkinv_4_2/A BR64_1/C[12] vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_350 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_361 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_372 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_383 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_394 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2050 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2061 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2072 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2083 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2094 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1360 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1371 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1382 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1393 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5604 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5615 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5626 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5637 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4903 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4914 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4925 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4936 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4947 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4958 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4969 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_180 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_10 BR32_0/RESET sky130_fd_sc_hd__o22ai_1_5/B1 sky130_fd_sc_hd__nor2_1_4/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_191 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1190 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3509 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2808 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2819 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR64_1 BR64_1/OUT vccd1 BR64_1/RESET BR64_1/C[0] BR64_1/C[1] BR64_1/C[2] BR64_1/C[3]
+ BR64_1/C[4] BR64_1/C[5] BR64_1/C[6] BR64_1/C[7] BR64_1/C[8] BR64_1/C[9] BR64_1/C[10]
+ BR64_1/C[11] BR64_1/C[12] BR64_1/C[13] BR64_1/C[14] BR64_1/C[15] BR64_1/C[16] BR64_1/C[17]
+ BR64_1/C[18] BR64_1/C[19] BR64_1/C[20] BR64_1/C[21] BR64_1/C[22] BR64_1/C[23] BR64_1/C[24]
+ BR64_1/C[25] BR64_1/C[26] BR64_1/C[27] BR64_1/C[28] BR64_1/C[29] BR64_1/C[30] BR64_1/C[31]
+ BR64_1/C[32] BR64_1/C[33] BR64_1/C[34] BR64_1/C[35] BR64_1/C[36] BR64_1/C[37] BR64_1/C[38]
+ BR64_1/C[39] BR64_1/C[40] BR64_1/C[41] BR64_1/C[42] BR64_1/C[43] BR64_1/C[44] BR64_1/C[45]
+ BR64_1/C[46] BR64_1/C[47] BR64_1/C[48] BR64_1/C[49] BR64_1/C[50] BR64_1/C[51] BR64_1/C[52]
+ BR64_1/C[53] BR64_1/C[54] BR64_1/C[55] BR64_1/C[56] BR64_1/C[57] BR64_1/C[58] BR64_1/C[59]
+ BR64_1/C[60] BR64_1/C[61] BR64_1/C[62] BR64_1/C[63] vssd1 BR64
Xsky130_fd_sc_hd__decap_12_5401 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5412 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_18 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5423 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_29 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5434 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4700 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5445 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4711 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5456 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5467 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4722 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5478 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4733 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_2 vccd1 vssd1 BR64_1/C[27] sky130_fd_sc_hd__buf_6_2/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__decap_12_4744 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5489 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4755 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4766 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4777 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4788 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4799 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2_1_3 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__nor2_1_5/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_3/a_109_297#
+ sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_3_0 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_12_905 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_916 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_927 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_938 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_949 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4007 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4018 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4029 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3306 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3317 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3328 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3339 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2605 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2616 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2627 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2638 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1904 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2649 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1915 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1926 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1937 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1948 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1959 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5220 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5231 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5242 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5253 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5264 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4530 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5275 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4541 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5286 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4552 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5297 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4563 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4574 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3840 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4585 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3851 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4596 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3862 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3873 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3884 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3895 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_30 NBR128_1/C[97] rstn NBR128_1/C[96] sky130_fd_sc_hd__clkinv_8_5/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_41 NBR128_0/C[86] sky130_fd_sc_hd__clkbuf_4_1/A BR128_1/C[85]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_52 sky130_fd_sc_hd__buf_6_7/A sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_1/C[74] sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_63 NBR128_1/C[64] sky130_fd_sc_hd__clkbuf_4_1/X NBR64_1/C[63]
+ sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_74 NBR64_1/C[53] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[52]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_85 NBR64_1/C[42] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[41]
+ sky130_fd_sc_hd__clkinv_8_5/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_96 BR32_0/C[31] sky130_fd_sc_hd__clkbuf_4_1/A sky130_fd_sc_hd__dfrtp_2_97/Q
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkinv_8_9 sky130_fd_sc_hd__clkinv_8_9/Y sky130_fd_sc_hd__clkinv_8_9/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_702 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_713 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_724 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_735 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_746 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_757 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_120 sky130_fd_sc_hd__clkbuf_8_2/A sky130_fd_sc_hd__clkbuf_4_1/X
+ BR64_1/C[6] sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_768 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_779 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3103 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3114 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3125 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3136 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2402 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3147 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2413 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3158 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3169 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2424 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2435 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1701 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2446 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1712 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2457 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1723 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2468 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1734 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2479 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1745 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1756 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1767 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1778 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1789 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5050 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5061 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5072 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5083 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5094 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4360 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4371 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4382 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4393 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3670 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3681 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3692 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2980 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2991 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1008 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1019 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_510 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_521 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_532 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_543 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_554 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_565 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_576 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_587 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_598 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2210 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2232 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2243 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2254 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1520 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2265 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1531 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2276 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1542 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2287 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1553 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2298 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1564 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1575 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1586 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1597 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4190 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_3 BR64_1/C[59] NBR64_1/C[59] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_4_3 sky130_fd_sc_hd__clkinv_4_3/A BR64_1/C[5] vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_340 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_351 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_362 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_373 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_384 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_395 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2040 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2051 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2062 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2073 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2084 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1350 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2095 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1361 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1372 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1383 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1394 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5605 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5616 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5627 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5638 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4904 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4915 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4926 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4937 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4948 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4959 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_170 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_181 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_11 BR64_0/RESET sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__nand2_1_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_192 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1180 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1191 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2809 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5402 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_19 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5413 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5424 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5435 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4701 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5446 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4712 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5457 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4723 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5468 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4734 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5479 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_3 vccd1 vssd1 BR64_1/C[26] sky130_fd_sc_hd__buf_6_3/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__decap_12_4745 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4756 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4767 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4778 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4789 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2_1_4 sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__nor2_1_4/Y
+ sky130_fd_sc_hd__nor2_1_5/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_4/a_109_297#
+ sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_3_1 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_12_906 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_917 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_928 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_939 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4008 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4019 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3307 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3318 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3329 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2606 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2628 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2639 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1905 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1916 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1927 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1938 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1949 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5210 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5232 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5243 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5254 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4520 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5265 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4531 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5276 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4542 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5287 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4553 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5298 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4564 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3830 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4575 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4586 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3841 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4597 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3852 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3863 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3874 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3885 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3896 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_20 NBR128_0/C[107] sky130_fd_sc_hd__clkbuf_4_1/A NBR128_1/C[106]
+ sky130_fd_sc_hd__clkinv_8_5/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_31 NBR128_1/C[96] sky130_fd_sc_hd__clkbuf_4_1/A NBR128_1/C[95]
+ sky130_fd_sc_hd__clkinv_8_5/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_42 NBR128_0/C[85] sky130_fd_sc_hd__clkbuf_4_1/A sky130_fd_sc_hd__buf_6_10/A
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_53 sky130_fd_sc_hd__buf_6_9/A sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_1/C[73] sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_64 NBR64_1/C[63] sky130_fd_sc_hd__clkbuf_4_1/X NBR64_1/C[62]
+ sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_75 NBR64_1/C[52] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[51]
+ sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_86 NBR64_1/C[41] sky130_fd_sc_hd__clkbuf_4_1/A NBR64_1/C[40]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_97 sky130_fd_sc_hd__dfrtp_2_97/Q sky130_fd_sc_hd__clkbuf_4_1/A
+ BR64_1/C[29] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_703 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_714 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_725 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_736 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_747 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_110 NBR64_1/C[17] sky130_fd_sc_hd__clkbuf_4_1/A BR32_0/C[16]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_758 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_121 sky130_fd_sc_hd__clkbuf_8_3/A sky130_fd_sc_hd__clkbuf_4_1/X
+ BR32_0/C[5] sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_769 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3104 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3115 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3126 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3137 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2403 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3148 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2414 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3159 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2425 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2436 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1702 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2447 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1713 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2458 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1724 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2469 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1735 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1746 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1757 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1768 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1779 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5040 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5051 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5062 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5073 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5084 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4350 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5095 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4361 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4372 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4383 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4394 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3660 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3671 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3682 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3693 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2970 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2981 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2992 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1009 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR32_0 BR32_0/C[31] BR64_1/C[30] BR64_1/C[29] BR64_1/C[28] BR64_1/C[27] BR64_1/C[26]
+ BR64_1/C[25] BR64_1/C[24] BR64_1/C[23] BR64_1/C[22] BR64_1/C[21] BR64_1/C[20] BR64_1/C[19]
+ BR64_1/C[18] BR64_1/C[17] BR32_0/C[16] BR32_0/C[15] BR32_0/C[14] BR32_1/C[13] BR64_1/C[12]
+ BR64_1/C[11] BR64_1/C[10] BR64_1/C[9] BR64_1/C[8] BR64_1/C[7] BR64_1/C[6] BR32_0/C[5]
+ BR64_1/C[4] BR32_0/C[3] BR64_1/C[2] BR64_1/C[1] BR64_1/C[0] vssd1 vccd1 BR32_0/RESET
+ BR32_0/OUT BR32
Xsky130_fd_sc_hd__decap_12_500 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_511 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_522 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_533 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_544 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_555 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_566 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_577 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_588 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_599 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2200 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2211 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2222 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2233 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2244 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1510 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2255 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1521 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2266 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1532 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2277 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1543 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2288 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2299 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1554 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1565 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1576 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1587 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1598 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4180 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4191 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3490 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_4 BR64_1/C[58] NBR64_1/C[58] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_4_4 sky130_fd_sc_hd__clkinv_4_4/A BR64_1/C[3] vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_330 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_341 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_352 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_363 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_374 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_385 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_396 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2030 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2041 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2052 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2063 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2074 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1340 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2085 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1351 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2096 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1362 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1373 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1384 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1395 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5606 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5628 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5639 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4905 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4916 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4927 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4938 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4949 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_160 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_171 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_12 sky130_fd_sc_hd__o21ai_1_1/B1 BR128_1/OUT sky130_fd_sc_hd__nor2_1_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_182 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_193 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1170 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1181 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1192 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5403 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5414 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5425 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5436 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4702 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5447 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5458 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4713 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5469 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4724 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4735 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_4 vccd1 vssd1 BR64_1/C[24] sky130_fd_sc_hd__buf_6_4/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__decap_12_4746 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4757 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4768 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4779 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2_1_5 sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__nor2_1_5/Y
+ sky130_fd_sc_hd__nor2_1_5/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_3_2 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_12_907 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_918 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_929 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4009 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3308 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3319 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2607 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2618 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1906 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1917 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1928 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1939 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5200 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5211 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5222 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5233 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5244 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4510 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5255 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4521 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5266 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4532 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5277 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4543 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5288 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4554 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5299 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3820 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4565 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3831 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4576 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3842 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4587 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3853 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4598 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3864 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3875 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3886 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3897 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_10 NBR128_0/C[117] sky130_fd_sc_hd__clkbuf_4_1/X NBR128_0/C[116]
+ sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_21 NBR128_1/C[106] rstn NBR128_1/C[105] sky130_fd_sc_hd__clkinv_8_5/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_32 NBR128_1/C[95] sky130_fd_sc_hd__clkbuf_4_1/A NBR128_1/C[94]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_43 sky130_fd_sc_hd__buf_6_10/A sky130_fd_sc_hd__clkbuf_4_1/A
+ BR128_1/C[83] sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_54 sky130_fd_sc_hd__dfrtp_2_54/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_1/C[72] sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_65 NBR64_1/C[62] sky130_fd_sc_hd__clkbuf_4_1/X NBR64_1/C[61]
+ sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_76 NBR64_1/C[51] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[50]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_87 NBR64_1/C[40] sky130_fd_sc_hd__clkbuf_4_1/A NBR64_1/C[39]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_98 NBR64_1/C[29] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[28]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_704 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_715 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_726 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_737 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_100 sky130_fd_sc_hd__buf_6_2/A sky130_fd_sc_hd__clkbuf_4_1/A
+ BR64_1/C[26] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_748 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_111 BR32_0/C[16] sky130_fd_sc_hd__clkbuf_4_1/A BR32_0/C[15]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_759 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_122 BR32_0/C[5] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[4]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_3105 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3116 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3127 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3138 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2404 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3149 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2415 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2426 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2437 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1703 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2448 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1714 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2459 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1725 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1736 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1747 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1758 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1769 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5030 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5041 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5052 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5063 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5074 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4340 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5085 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4351 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5096 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4362 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4373 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4384 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3650 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4395 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3661 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3672 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3683 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3694 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2960 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2971 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2982 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2993 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR32_1 BR64_1/C[31] BR64_1/C[30] BR64_1/C[29] BR64_1/C[28] BR64_1/C[27] BR64_1/C[26]
+ BR64_1/C[25] BR64_1/C[24] BR64_1/C[23] BR64_1/C[22] BR64_1/C[21] BR64_1/C[20] BR64_1/C[19]
+ BR64_1/C[18] BR64_1/C[17] BR64_1/C[16] BR64_1/C[15] BR32_1/C[14] BR32_1/C[13] BR64_1/C[12]
+ BR64_1/C[11] BR64_1/C[10] BR64_1/C[9] BR64_1/C[8] BR64_1/C[7] BR64_1/C[6] BR64_1/C[5]
+ BR64_1/C[4] BR64_1/C[3] BR64_1/C[2] BR64_1/C[1] BR64_1/C[0] vssd1 vccd1 BR32_1/RESET
+ BR32_1/OUT BR32
Xsky130_fd_sc_hd__decap_12_501 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_512 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_523 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_534 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_545 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_556 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_567 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_578 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_589 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2201 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2212 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2223 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2234 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1500 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2245 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1511 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2256 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1522 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2267 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1533 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2278 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1544 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2289 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1555 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1566 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1577 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1588 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1599 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o22ai_1_0 sky130_fd_sc_hd__o22ai_1_2/Y sky130_fd_sc_hd__nor2_1_1/B
+ sky130_fd_sc_hd__o22ai_1_0/Y puf_sel1 sky130_fd_sc_hd__o22ai_1_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__decap_12_4170 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4181 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4192 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3480 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3491 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2790 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_5 BR64_1/C[55] NBR64_1/C[55] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_4_5 sky130_fd_sc_hd__clkinv_4_5/A BR64_1/C[2] vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_320 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_331 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_342 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_353 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_364 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_375 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_386 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_397 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2020 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2031 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2042 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2053 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2064 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1330 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2075 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1341 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2086 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1352 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2097 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1363 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1374 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1385 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1396 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5607 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5618 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4906 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4917 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4928 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4939 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_150 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_161 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_172 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_183 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_13 BR32_1/RESET sky130_fd_sc_hd__o22ai_1_6/B1 sky130_fd_sc_hd__nor2_1_5/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_194 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1160 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1171 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1182 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1193 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5404 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5415 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5426 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5437 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4703 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5448 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4714 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5459 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4725 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4736 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_5 vccd1 vssd1 BR64_1/C[1] NBR32_1/C[1] vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__decap_12_4747 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4758 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4769 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_3_3 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_12_908 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_919 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3309 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2608 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2619 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1907 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1918 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1929 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5201 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5212 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5223 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5234 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4500 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5245 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4511 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5256 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4522 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5267 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4533 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5278 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4544 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5289 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3810 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4555 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3821 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4566 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3832 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4577 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4588 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3843 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3854 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4599 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3865 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3876 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3887 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3898 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_11 NBR128_0/C[116] sky130_fd_sc_hd__clkbuf_4_1/X BR128_1/C[115]
+ sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_22 NBR128_1/C[105] rstn NBR128_1/C[104] sky130_fd_sc_hd__clkinv_8_5/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_33 NBR128_1/C[94] sky130_fd_sc_hd__clkbuf_4_1/A NBR128_1/C[93]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_44 NBR128_0/C[83] sky130_fd_sc_hd__clkbuf_4_1/X BR128_1/C[82]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_55 sky130_fd_sc_hd__dfrtp_2_55/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_1/C[71] sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_66 NBR64_1/C[61] sky130_fd_sc_hd__clkbuf_4_1/X NBR64_1/C[60]
+ sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_77 NBR64_1/C[50] sky130_fd_sc_hd__clkbuf_4_1/X NBR64_1/C[49]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_88 NBR64_1/C[39] sky130_fd_sc_hd__clkbuf_4_1/A NBR64_1/C[38]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_99 sky130_fd_sc_hd__buf_6_1/A sky130_fd_sc_hd__clkbuf_4_1/A
+ BR64_1/C[27] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_705 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_716 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_727 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_738 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_101 sky130_fd_sc_hd__buf_6_3/A sky130_fd_sc_hd__clkbuf_4_1/A
+ BR64_1/C[25] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_749 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_112 BR32_0/C[15] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[14]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_123 sky130_fd_sc_hd__clkbuf_8_4/A sky130_fd_sc_hd__clkbuf_4_1/X
+ BR32_0/C[3] sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_3106 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3117 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3128 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3139 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2405 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2416 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2427 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2438 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1704 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2449 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1715 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1726 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1737 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1748 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1759 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5020 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5031 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5042 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5053 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5064 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4330 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5075 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4341 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5086 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4352 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5097 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4363 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4374 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3640 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4385 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3651 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4396 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3662 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3684 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2950 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3695 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2961 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2972 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2983 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2994 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_502 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_513 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_524 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_535 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_546 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_568 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_579 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2202 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2213 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2224 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2235 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1501 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2246 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1512 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2257 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1523 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2268 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1534 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2279 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1545 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1556 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1567 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1578 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1589 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o22ai_1_1 sky130_fd_sc_hd__o22ai_1_1/A2 sky130_fd_sc_hd__nand2_1_2/B
+ sky130_fd_sc_hd__o22ai_1_1/Y puf_sel0 sky130_fd_sc_hd__o22ai_1_1/B2 vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__decap_12_4160 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4171 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4182 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4193 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3470 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3481 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3492 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2780 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2791 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_6 BR64_1/C[54] NBR64_1/C[54] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_310 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_321 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_332 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_343 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_354 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_365 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_376 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_387 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_398 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2010 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2021 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2032 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2043 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2054 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1320 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2065 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1331 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2076 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1342 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2087 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1353 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2098 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1364 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1375 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1386 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1397 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5608 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5619 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4907 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4918 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4929 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_0 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_5/A sky130_fd_sc_hd__o22ai_1_5/Y
+ sky130_fd_sc_hd__nand2_1_9/Y sky130_fd_sc_hd__o21ai_1_0/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_140 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_151 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_162 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_173 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_14 BR64_1/RESET sky130_fd_sc_hd__nor2_1_5/Y sky130_fd_sc_hd__nand2_1_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_184 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_195 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1150 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1161 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1172 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1183 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1194 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5405 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5416 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5427 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5438 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4704 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5449 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4715 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4726 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4737 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_6 vccd1 vssd1 BR64_1/C[0] sky130_fd_sc_hd__buf_6_6/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__decap_12_4748 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4759 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_909 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2609 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1908 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1919 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5202 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5213 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5224 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5235 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4501 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5246 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4512 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5257 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4523 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5268 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4534 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5279 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4545 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3800 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3811 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4556 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3822 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4567 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3833 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4578 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3844 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4589 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3855 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3866 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3877 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3888 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3899 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_12 sky130_fd_sc_hd__dfrtp_2_12/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_0/C[114] sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_23 NBR128_1/C[104] rstn NBR128_1/C[103] sky130_fd_sc_hd__clkinv_8_5/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_34 NBR128_1/C[93] sky130_fd_sc_hd__clkbuf_4_1/A NBR128_1/C[92]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_45 NBR128_0/C[82] sky130_fd_sc_hd__clkbuf_4_1/X NBR128_0/C[81]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_56 sky130_fd_sc_hd__dfrtp_2_56/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_1/C[70] sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_67 NBR64_1/C[60] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[59]
+ sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_78 NBR64_1/C[49] sky130_fd_sc_hd__clkbuf_4_1/X NBR64_1/C[48]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_89 NBR64_1/C[38] sky130_fd_sc_hd__clkbuf_4_1/A NBR64_0/C[37]
+ sky130_fd_sc_hd__clkinv_8_5/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_706 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_717 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_728 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_739 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_102 NBR64_1/C[25] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[24]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_113 BR32_0/C[14] sky130_fd_sc_hd__clkbuf_4_1/A NBR32_1/C[13]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_124 BR32_0/C[3] sky130_fd_sc_hd__clkbuf_4_1/X sky130_fd_sc_hd__dfrtp_2_125/Q
+ sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_3107 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3118 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3129 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2406 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2417 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2428 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2439 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1705 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1716 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1727 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1738 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1749 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5010 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5021 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5032 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5043 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5054 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4320 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5065 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4331 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5076 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_0 vccd1 vssd1 NBR64_0/C[16] BR32_0/C[16] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_4342 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5087 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4353 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5098 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4364 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3630 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4375 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4386 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3652 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4397 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3663 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3674 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2940 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3696 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2951 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2962 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2973 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2984 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2995 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_503 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_514 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_525 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_536 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_547 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_558 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_569 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2203 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2214 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2225 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2236 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1502 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2247 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1513 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2258 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1524 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2269 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1535 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1546 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1568 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1579 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o22ai_1_2 sky130_fd_sc_hd__o21ai_1_1/Y sky130_fd_sc_hd__nand2_1_2/B
+ sky130_fd_sc_hd__o22ai_1_2/Y puf_sel0 sky130_fd_sc_hd__o21ai_1_0/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__decap_12_4150 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4161 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4172 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4183 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4194 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3460 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3471 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3482 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3493 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2770 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2781 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2792 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_7 BR64_1/C[52] NBR64_1/C[52] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_300 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_311 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_322 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_333 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_344 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_355 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_366 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_377 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_388 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_399 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2000 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2011 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2022 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2033 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2044 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2055 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1310 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1321 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2066 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1332 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2077 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1343 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2088 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1354 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2099 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1365 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1376 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1387 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1398 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3290 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5609 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4908 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4919 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_5/A sky130_fd_sc_hd__o22ai_1_6/Y
+ sky130_fd_sc_hd__o21ai_1_1/B1 sky130_fd_sc_hd__o21ai_1_1/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_130 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_141 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_152 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_163 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_174 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_185 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_196 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1140 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1151 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1162 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1173 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1184 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1195 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5406 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5417 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5428 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5439 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4705 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4716 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4727 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4738 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_7 vccd1 vssd1 BR128_1/C[75] sky130_fd_sc_hd__buf_6_7/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__decap_12_4749 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1909 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5203 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5214 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5225 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5236 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4502 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5247 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4513 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5258 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4524 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5269 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4535 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3801 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4546 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3812 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3823 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4568 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3834 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4579 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3845 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3856 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3867 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3878 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3889 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_13 BR128_0/C[114] sky130_fd_sc_hd__clkbuf_4_1/X BR128_0/C[113]
+ sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_24 NBR128_1/C[103] rstn NBR128_1/C[102] sky130_fd_sc_hd__clkinv_8_5/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_35 NBR128_1/C[92] sky130_fd_sc_hd__clkbuf_4_1/A BR128_1/C[91]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_46 NBR128_0/C[81] sky130_fd_sc_hd__clkbuf_4_1/X BR128_1/C[80]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_57 sky130_fd_sc_hd__dfrtp_2_57/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_1/C[69] sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_68 NBR64_1/C[59] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[58]
+ sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_79 NBR64_1/C[48] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[47]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkbuf_4_60 BR64_1/C[16] BR32_0/C[16] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_707 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_718 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_729 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_103 sky130_fd_sc_hd__buf_6_4/A sky130_fd_sc_hd__clkbuf_4_1/A
+ NBR64_1/C[23] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_114 NBR32_1/C[13] sky130_fd_sc_hd__clkbuf_4_1/A NBR32_1/C[12]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_125 sky130_fd_sc_hd__dfrtp_2_125/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR64_1/C[1] sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_3108 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3119 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2407 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2418 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2429 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1706 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1717 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1728 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1739 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5000 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5011 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5022 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5033 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5044 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4310 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5055 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4321 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5066 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4332 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5077 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_1 vccd1 vssd1 BR128_1/C[68] BR128_0/C[68] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_4343 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5088 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4354 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5099 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3620 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4365 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3631 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4376 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3642 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4387 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3653 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4398 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3664 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2930 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3675 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2941 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3686 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2952 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2963 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2974 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2985 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2996 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_504 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_515 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_526 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_537 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_548 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_559 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2204 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2215 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2226 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2237 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1503 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2248 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1514 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2259 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1525 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1536 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1547 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1558 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1569 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o22ai_1_3 NBR32_0/OUT sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__o22ai_1_3/Y
+ length0 NBR64_0/OUT vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__decap_12_4140 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4151 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4162 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4173 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4184 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3450 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4195 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3461 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3472 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3483 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3494 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2760 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2771 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2782 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2793 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_8 BR64_1/C[51] NBR64_1/C[51] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_301 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_312 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_323 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_334 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_345 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_356 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_367 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_378 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_389 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2001 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2012 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2023 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2034 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1300 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2045 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1311 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2056 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1322 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2067 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1333 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2078 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1344 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2089 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1355 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1366 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1377 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1388 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1399 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_890 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3280 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3291 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2590 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4909 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_120 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_131 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_142 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_153 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_164 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_175 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_186 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_197 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1130 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1141 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1152 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1163 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1174 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1185 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1196 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5407 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5418 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5429 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4706 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4717 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4728 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4739 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_8 vccd1 vssd1 BR128_1/C[88] sky130_fd_sc_hd__buf_6_8/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__decap_12_5204 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5215 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5226 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5237 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4503 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5248 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4514 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5259 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4525 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4536 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4547 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3802 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3813 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4558 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3824 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4569 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3835 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3846 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3857 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3868 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3879 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_14 BR128_0/C[113] sky130_fd_sc_hd__clkbuf_4_1/X BR128_1/C[112]
+ sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_25 NBR128_1/C[102] rstn NBR128_1/C[101] sky130_fd_sc_hd__clkinv_8_5/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_36 sky130_fd_sc_hd__dfrtp_2_36/Q sky130_fd_sc_hd__clkbuf_4_1/A
+ BR128_1/C[90] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_47 NBR128_0/C[80] sky130_fd_sc_hd__clkbuf_4_1/X NBR128_0/C[79]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_58 sky130_fd_sc_hd__dfrtp_2_58/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ NBR128_1/C[68] sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_69 NBR64_1/C[58] sky130_fd_sc_hd__clkbuf_4_1/X NBR64_1/C[57]
+ sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkbuf_4_50 BR64_1/C[39] NBR64_1/C[39] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_61 NBR64_1/C[15] BR32_0/C[15] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_708 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_719 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_104 NBR64_1/C[23] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[22]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_115 NBR32_1/C[12] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[11]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_126 NBR32_1/C[1] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[0]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_3109 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2408 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2419 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1707 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1718 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1729 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5001 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5012 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5023 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5034 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4300 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5045 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4311 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5056 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4322 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5067 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4333 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5078 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_2 vccd1 vssd1 NBR64_1/C[31] BR32_0/C[31] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_4344 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5089 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4355 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3610 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3621 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4366 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3632 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4377 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3643 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4388 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3654 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4399 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2920 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3665 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2931 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3676 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2942 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3687 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3698 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2953 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2964 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2975 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2986 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2997 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5590 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_505 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_516 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_527 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_538 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_549 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2205 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2216 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2227 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2238 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1504 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2249 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1515 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1526 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1537 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1548 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1559 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o22ai_1_4 NBR32_1/OUT sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__o22ai_1_4/Y
+ sky130_fd_sc_hd__nand2_1_8/A NBR64_1/OUT vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__decap_12_4130 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4141 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4152 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4163 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4174 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3440 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4185 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3451 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4196 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3462 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3473 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3484 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2750 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3495 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2761 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2772 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2783 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2794 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_9 BR64_1/C[50] NBR64_1/C[50] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_302 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_313 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_324 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_335 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_346 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_357 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_368 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_379 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2002 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2013 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2024 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2035 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2046 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1301 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2057 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1312 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1323 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2068 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1334 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2079 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1345 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1356 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1367 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1378 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1389 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_880 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_891 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3270 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3281 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3292 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2580 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2591 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1890 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_110 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_121 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_132 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_143 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_154 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_165 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_176 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_187 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_198 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1120 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1131 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1142 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1153 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1164 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1175 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XNBR128_0 NBR128_0/RESET BR64_1/C[0] BR64_1/C[1] BR64_1/C[2] BR64_1/C[3] BR64_1/C[4]
+ BR64_1/C[5] BR64_1/C[7] BR64_1/C[8] BR64_1/C[9] BR64_1/C[10] BR64_1/C[11] BR64_1/C[12]
+ BR64_1/C[13] BR64_1/C[14] NBR64_1/C[15] NBR64_0/C[16] NBR64_0/C[17] NBR64_0/C[18]
+ NBR64_1/C[19] NBR64_1/C[20] NBR64_1/C[21] NBR64_1/C[22] NBR64_1/C[23] BR64_1/C[24]
+ NBR64_1/C[25] BR64_1/C[26] BR64_1/C[27] BR64_1/C[28] NBR64_1/C[29] BR64_1/C[30]
+ BR64_1/C[6] NBR64_1/C[31] NBR64_1/C[32] NBR64_1/C[33] NBR64_1/C[34] NBR64_1/C[35]
+ NBR64_1/C[36] NBR64_0/C[37] NBR64_1/C[38] NBR64_1/C[39] NBR64_1/C[40] NBR64_1/C[41]
+ NBR64_1/C[42] NBR64_1/C[43] NBR64_1/C[44] NBR64_1/C[45] NBR64_1/C[46] NBR64_1/C[47]
+ NBR64_1/C[48] NBR64_1/C[49] NBR64_1/C[50] NBR64_1/C[51] NBR64_1/C[52] NBR64_1/C[53]
+ NBR64_1/C[54] NBR64_1/C[55] NBR64_1/C[56] NBR64_1/C[57] NBR64_1/C[58] NBR64_1/C[59]
+ NBR64_1/C[60] NBR64_1/C[61] NBR64_1/C[62] NBR128_1/C[95] NBR128_1/C[96] NBR128_1/C[97]
+ NBR128_1/C[98] NBR128_1/C[99] NBR128_1/C[100] NBR128_1/C[101] NBR128_1/C[102] NBR128_1/C[103]
+ NBR128_1/C[104] NBR128_1/C[105] NBR128_1/C[106] NBR128_0/C[107] NBR128_1/C[108]
+ NBR128_1/C[109] NBR128_1/C[110] NBR128_0/C[111] BR128_1/C[112] BR128_0/C[113] BR128_0/C[114]
+ BR128_1/C[115] NBR128_0/C[116] NBR128_0/C[117] BR128_1/C[118] BR128_1/C[119] BR128_0/C[120]
+ BR128_0/C[121] BR128_1/C[122] BR128_0/C[123] BR128_0/C[124] BR128_0/C[125] BR128_0/C[126]
+ NBR128_1/C[127] NBR64_1/C[63] NBR128_1/C[64] NBR128_1/C[65] BR128_0/C[66] BR128_0/C[67]
+ NBR128_1/C[68] BR128_1/C[69] BR128_1/C[70] BR128_1/C[71] BR128_1/C[72] BR128_1/C[73]
+ BR128_1/C[74] BR128_1/C[75] NBR128_0/C[76] NBR128_0/C[77] NBR128_0/C[78] NBR128_0/C[79]
+ NBR128_0/C[80] NBR128_0/C[81] NBR128_0/C[82] NBR128_0/C[83] BR128_1/C[84] NBR128_0/C[85]
+ NBR128_0/C[86] NBR128_0/C[87] BR128_1/C[88] BR128_1/C[89] BR128_1/C[90] BR128_1/C[91]
+ NBR128_1/C[92] NBR128_1/C[93] NBR128_1/C[94] NBR128_0/OUT vccd1 vssd1 NBR128
Xsky130_fd_sc_hd__decap_12_1186 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1197 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5408 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5419 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_0 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4707 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4718 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4729 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_9 vccd1 vssd1 BR128_1/C[74] sky130_fd_sc_hd__buf_6_9/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
XNBR64_0 NBR64_0/OUT vccd1 NBR64_0/RESET BR64_1/C[0] BR64_1/C[1] BR64_1/C[2] BR64_1/C[3]
+ BR64_1/C[4] BR64_1/C[5] BR64_1/C[6] BR64_1/C[7] BR64_1/C[8] BR64_1/C[9] BR64_1/C[10]
+ BR64_1/C[11] BR64_1/C[12] BR64_1/C[13] BR64_1/C[14] NBR64_1/C[15] NBR64_0/C[16]
+ NBR64_0/C[17] NBR64_0/C[18] NBR64_1/C[19] NBR64_1/C[20] NBR64_1/C[21] NBR64_1/C[22]
+ NBR64_1/C[23] BR64_1/C[24] NBR64_1/C[25] BR64_1/C[26] BR64_1/C[27] BR64_1/C[28]
+ NBR64_1/C[29] BR64_1/C[30] NBR64_1/C[31] NBR64_1/C[32] NBR64_1/C[33] NBR64_1/C[34]
+ NBR64_1/C[35] NBR64_1/C[36] NBR64_0/C[37] NBR64_1/C[38] NBR64_1/C[39] NBR64_1/C[40]
+ NBR64_1/C[41] NBR64_1/C[42] NBR64_1/C[43] NBR64_1/C[44] NBR64_1/C[45] NBR64_1/C[46]
+ NBR64_1/C[47] NBR64_1/C[48] NBR64_1/C[49] NBR64_1/C[50] NBR64_1/C[51] NBR64_1/C[52]
+ NBR64_1/C[53] NBR64_1/C[54] NBR64_1/C[55] NBR64_1/C[56] NBR64_1/C[57] NBR64_1/C[58]
+ NBR64_1/C[59] NBR64_1/C[60] NBR64_1/C[61] NBR64_1/C[62] NBR64_1/C[63] vssd1 NBR64
Xsky130_fd_sc_hd__decap_12_5205 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5216 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5227 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5238 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4504 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5249 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4515 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4526 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4537 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3803 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4548 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3814 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4559 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3825 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3836 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3847 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3858 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3869 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_15 sky130_fd_sc_hd__dfrtp_2_15/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ NBR128_0/C[111] sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_26 NBR128_1/C[101] rstn NBR128_1/C[100] sky130_fd_sc_hd__clkinv_8_5/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_37 sky130_fd_sc_hd__dfrtp_2_37/Q sky130_fd_sc_hd__clkbuf_4_1/A
+ BR128_1/C[89] sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_48 NBR128_0/C[79] sky130_fd_sc_hd__clkbuf_4_1/X NBR128_0/C[78]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_59 NBR128_1/C[68] sky130_fd_sc_hd__clkbuf_4_1/X BR128_0/C[67]
+ sky130_fd_sc_hd__clkinv_8_10/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkbuf_4_40 BR64_1/C[56] NBR64_1/C[56] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_51 BR64_1/C[38] NBR64_1/C[38] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_62 BR64_1/C[15] BR32_0/C[15] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_709 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_105 NBR64_1/C[22] sky130_fd_sc_hd__clkbuf_4_1/A NBR64_1/C[21]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_116 sky130_fd_sc_hd__buf_12_0/A sky130_fd_sc_hd__clkbuf_4_1/A
+ BR64_1/C[10] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_127 sky130_fd_sc_hd__buf_6_6/A sky130_fd_sc_hd__clkbuf_4_1/X
+ si sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_2409 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1708 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1719 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_10 sky130_fd_sc_hd__clkinv_8_10/Y sky130_fd_sc_hd__clkinv_8_9/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_5002 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5013 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5024 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5035 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4301 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5046 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4312 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5057 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4323 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5068 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4334 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5079 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_3 vccd1 vssd1 so NBR128_1/C[127] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_3600 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4345 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3611 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4356 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3622 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4367 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3633 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4378 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3644 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4389 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3655 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2910 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2921 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3666 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2932 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3677 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2943 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3688 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2954 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3699 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2965 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2976 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2987 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2998 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5580 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5591 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4890 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_506 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_517 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_528 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_539 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2206 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2217 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2228 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2239 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1505 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1516 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1527 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1538 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1549 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o22ai_1_5 BR32_0/OUT sky130_fd_sc_hd__o22ai_1_5/B1 sky130_fd_sc_hd__o22ai_1_5/Y
+ sky130_fd_sc_hd__nand2_1_8/A BR64_0/OUT vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__decap_12_4120 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4131 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4142 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4153 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4164 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3430 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4175 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3441 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4186 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3452 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4197 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3463 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3474 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2740 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3485 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2751 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3496 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2762 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2773 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2784 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2795 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_303 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_314 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_325 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_336 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_347 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_358 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_369 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2003 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2014 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2025 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2036 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1302 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2047 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1313 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2058 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1324 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2069 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1335 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1346 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1357 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1368 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1379 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_870 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_881 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_892 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3260 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3271 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3282 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3293 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2570 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2581 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2592 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1880 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1891 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_100 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_111 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_122 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_133 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_144 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_155 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_166 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_177 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_188 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_199 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1110 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1121 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1132 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1143 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1154 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1165 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1176 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XNBR128_1 NBR128_1/RESET BR64_1/C[0] BR64_1/C[1] BR64_1/C[2] BR64_1/C[3] BR64_1/C[4]
+ BR64_1/C[5] BR64_1/C[7] BR64_1/C[8] BR64_1/C[9] BR64_1/C[10] BR64_1/C[11] BR64_1/C[12]
+ BR64_1/C[13] BR64_1/C[14] BR32_0/C[15] BR32_0/C[16] NBR64_1/C[17] NBR128_1/C[18]
+ NBR64_1/C[19] NBR64_1/C[20] NBR64_1/C[21] BR64_1/C[22] BR64_1/C[23] BR64_1/C[24]
+ BR64_1/C[25] BR64_1/C[26] BR64_1/C[27] BR64_1/C[28] BR64_1/C[29] BR64_1/C[30] BR64_1/C[6]
+ BR32_0/C[31] BR64_1/C[32] NBR64_1/C[33] BR64_1/C[34] BR64_1/C[35] BR64_1/C[36] BR64_1/C[37]
+ BR64_1/C[38] BR64_1/C[39] BR64_1/C[40] BR64_1/C[41] BR64_1/C[42] BR64_1/C[43] BR64_1/C[44]
+ BR64_1/C[45] BR64_1/C[46] BR64_1/C[47] NBR128_1/C[48] BR64_1/C[49] BR64_1/C[50]
+ BR64_1/C[51] BR64_1/C[52] BR64_1/C[53] BR64_1/C[54] BR64_1/C[55] BR64_1/C[56] BR64_1/C[57]
+ BR64_1/C[58] BR64_1/C[59] NBR64_1/C[60] NBR64_1/C[61] NBR64_1/C[62] NBR128_1/C[95]
+ NBR128_1/C[96] NBR128_1/C[97] NBR128_1/C[98] NBR128_1/C[99] NBR128_1/C[100] NBR128_1/C[101]
+ NBR128_1/C[102] NBR128_1/C[103] NBR128_1/C[104] NBR128_1/C[105] NBR128_1/C[106]
+ BR128_1/C[107] NBR128_1/C[108] NBR128_1/C[109] NBR128_1/C[110] BR128_1/C[111] BR128_1/C[112]
+ BR128_0/C[113] BR128_0/C[114] BR128_1/C[115] BR128_1/C[116] BR128_1/C[117] BR128_1/C[118]
+ BR128_1/C[119] BR128_0/C[120] BR128_0/C[121] BR128_1/C[122] BR128_0/C[123] BR128_0/C[124]
+ BR128_0/C[125] BR128_0/C[126] NBR128_1/C[127] NBR64_1/C[63] NBR128_1/C[64] NBR128_1/C[65]
+ BR128_0/C[66] BR128_0/C[67] NBR128_1/C[68] BR128_1/C[69] BR128_1/C[70] BR128_1/C[71]
+ BR128_1/C[72] BR128_1/C[73] BR128_1/C[74] BR128_1/C[75] BR128_1/C[76] BR128_1/C[77]
+ BR128_1/C[78] BR128_1/C[79] BR128_1/C[80] BR128_1/C[81] BR128_1/C[82] BR128_1/C[83]
+ BR128_1/C[84] BR128_1/C[85] BR128_1/C[86] BR128_1/C[87] BR128_1/C[88] BR128_1/C[89]
+ BR128_1/C[90] BR128_1/C[91] NBR128_1/C[92] NBR128_1/C[93] NBR128_1/C[94] NBR128_1/OUT
+ vccd1 vssd1 NBR128
Xsky130_fd_sc_hd__decap_12_1187 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1198 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3090 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5409 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4708 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4719 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XNBR64_1 NBR64_1/OUT vccd1 NBR64_1/RESET BR64_1/C[0] BR64_1/C[1] BR64_1/C[2] BR64_1/C[3]
+ BR64_1/C[4] BR64_1/C[5] BR64_1/C[6] BR64_1/C[7] BR64_1/C[8] BR64_1/C[9] BR64_1/C[10]
+ BR64_1/C[11] BR64_1/C[12] BR64_1/C[13] BR64_1/C[14] NBR64_1/C[15] BR32_0/C[16] NBR64_1/C[17]
+ NBR64_1/C[18] NBR64_1/C[19] NBR64_1/C[20] NBR64_1/C[21] NBR64_1/C[22] NBR64_1/C[23]
+ BR64_1/C[24] NBR64_1/C[25] BR64_1/C[26] BR64_1/C[27] BR64_1/C[28] NBR64_1/C[29]
+ BR64_1/C[30] NBR64_1/C[31] NBR64_1/C[32] NBR64_1/C[33] NBR64_1/C[34] NBR64_1/C[35]
+ NBR64_1/C[36] BR64_1/C[37] NBR64_1/C[38] NBR64_1/C[39] NBR64_1/C[40] NBR64_1/C[41]
+ NBR64_1/C[42] NBR64_1/C[43] NBR64_1/C[44] NBR64_1/C[45] NBR64_1/C[46] NBR64_1/C[47]
+ NBR64_1/C[48] NBR64_1/C[49] NBR64_1/C[50] NBR64_1/C[51] NBR64_1/C[52] NBR64_1/C[53]
+ NBR64_1/C[54] NBR64_1/C[55] NBR64_1/C[56] NBR64_1/C[57] NBR64_1/C[58] NBR64_1/C[59]
+ NBR64_1/C[60] NBR64_1/C[61] NBR64_1/C[62] NBR64_1/C[63] vssd1 NBR64
Xsky130_fd_sc_hd__decap_12_5206 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5217 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5228 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5239 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4505 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4516 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4527 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4538 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3804 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4549 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3815 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3826 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3837 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3848 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3859 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_16 NBR128_0/C[111] sky130_fd_sc_hd__clkbuf_4_1/X NBR128_1/C[110]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_27 NBR128_1/C[100] rstn NBR128_1/C[99] sky130_fd_sc_hd__clkinv_8_5/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_38 sky130_fd_sc_hd__dfrtp_2_38/Q sky130_fd_sc_hd__clkbuf_4_1/A
+ BR128_1/C[88] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_49 NBR128_0/C[78] sky130_fd_sc_hd__clkbuf_4_1/X BR128_1/C[77]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkbuf_4_30 BR128_1/C[69] sky130_fd_sc_hd__dfrtp_2_58/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_41 BR64_1/C[53] NBR64_1/C[53] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_52 BR64_1/C[37] NBR64_0/C[37] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_63 sky130_fd_sc_hd__o22ai_1_1/B2 sky130_fd_sc_hd__o21ai_0_0/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__dfrtp_2_106 NBR64_1/C[21] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[20]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_117 sky130_fd_sc_hd__buf_12_1/A sky130_fd_sc_hd__clkbuf_4_1/A
+ BR64_1/C[9] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1709 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5003 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5014 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5025 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5036 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4302 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5047 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5058 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4313 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4324 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5069 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4335 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_4 vccd1 vssd1 BR128_1/C[117] NBR128_0/C[117] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_4346 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3612 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4357 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3623 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4368 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3634 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4379 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2900 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2911 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3656 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2922 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3667 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2933 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3678 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3689 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2944 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2955 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2966 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2977 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2988 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2999 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5570 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5581 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5592 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4880 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4891 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_507 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_518 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_529 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2207 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2218 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2229 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1506 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1517 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1528 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1539 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o22ai_1_6 BR32_1/OUT sky130_fd_sc_hd__o22ai_1_6/B1 sky130_fd_sc_hd__o22ai_1_6/Y
+ sky130_fd_sc_hd__nand2_1_8/A BR64_1/OUT vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__decap_12_4110 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4121 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4132 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4143 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4154 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3420 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4165 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3431 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4176 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3442 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4187 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3453 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4198 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3464 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2730 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3475 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2741 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3486 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3497 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2752 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2763 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2774 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2785 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2796 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_304 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_315 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_326 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_337 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_348 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_359 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2004 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2015 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2026 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2037 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2048 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1303 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1314 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2059 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1325 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1336 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1347 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1358 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1369 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_860 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_871 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_882 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_893 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3250 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3261 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3272 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3283 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3294 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2560 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2571 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2582 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2593 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1870 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1881 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1892 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_101 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_112 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_123 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_134 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_145 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_156 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_167 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_178 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_189 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1100 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1111 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1122 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1133 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1144 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1155 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1166 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1177 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1188 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1199 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_690 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3080 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3091 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2390 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4709 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5207 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5218 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5229 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4506 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4517 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4528 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4539 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3805 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3816 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3827 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3838 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3849 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_17 NBR128_1/C[110] sky130_fd_sc_hd__clkbuf_4_1/A NBR128_1/C[109]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_28 NBR128_1/C[99] rstn NBR128_1/C[98] sky130_fd_sc_hd__clkinv_8_5/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_39 sky130_fd_sc_hd__buf_6_8/A sky130_fd_sc_hd__clkbuf_4_1/A
+ NBR128_0/C[87] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkbuf_4_20 BR128_1/C[85] NBR128_0/C[85] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_31 NBR64_1/C[19] sky130_fd_sc_hd__dfrtp_2_108/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_42 BR64_1/C[49] NBR64_1/C[49] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_53 BR64_1/C[34] NBR64_1/C[34] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_64 BR128_1/C[79] NBR128_0/C[79] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__dfrtp_2_107 NBR64_1/C[20] sky130_fd_sc_hd__clkbuf_4_1/A NBR64_1/C[19]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_118 sky130_fd_sc_hd__clkbuf_8_1/A sky130_fd_sc_hd__clkbuf_4_1/A
+ BR64_1/C[8] sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_5004 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5015 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5026 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5037 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4303 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5048 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4314 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5059 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4325 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4336 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_5 vccd1 vssd1 BR128_1/C[116] NBR128_0/C[116] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_3602 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4347 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4358 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3624 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4369 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3635 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3646 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2901 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2912 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2923 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3668 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2934 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3679 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2945 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2956 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2967 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2978 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2989 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5560 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5571 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5582 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5593 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4870 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4881 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4892 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_508 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_519 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2208 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2219 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1507 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1518 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1529 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XNBR32_0 NBR64_1/C[31] BR64_1/C[30] NBR64_1/C[29] BR64_1/C[28] BR64_1/C[27] BR64_1/C[26]
+ NBR64_1/C[25] BR64_1/C[24] NBR64_1/C[23] NBR64_1/C[22] NBR64_1/C[21] NBR64_1/C[20]
+ NBR64_1/C[19] NBR64_0/C[18] NBR64_0/C[17] NBR64_0/C[16] NBR64_1/C[15] BR64_1/C[14]
+ NBR32_1/C[13] NBR32_1/C[12] BR64_1/C[11] BR64_1/C[10] BR64_1/C[9] BR64_1/C[8] BR64_1/C[7]
+ BR64_1/C[6] BR64_1/C[5] BR64_1/C[4] BR64_1/C[3] BR64_1/C[2] BR64_1/C[1] BR64_1/C[0]
+ NBR32_0/RESET NBR32_0/OUT vccd1 vssd1 NBR32
Xsky130_fd_sc_hd__decap_12_4100 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4111 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4122 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4133 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4144 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3410 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4155 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3421 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4166 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3432 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4177 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3443 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4188 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3454 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4199 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2720 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3465 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2731 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3476 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2742 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3487 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2753 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3498 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2764 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2775 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2786 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2797 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_10 vssd1 vccd1 BR128_1/C[124] BR128_0/C[124] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_5390 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_305 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_316 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_327 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_338 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_349 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2005 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2016 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2027 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2038 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1304 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2049 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1315 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1326 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1337 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1348 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1359 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_850 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_861 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_872 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_883 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_894 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3240 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3251 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3262 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3273 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3284 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2550 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3295 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2561 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2572 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2583 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2594 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1860 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1871 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1882 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1893 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_102 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_113 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_124 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_135 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_146 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_157 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_168 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_179 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1101 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1112 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1123 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1134 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1145 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1156 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1167 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1178 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1189 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_680 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_691 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3070 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3081 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3092 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2380 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2391 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR128_0 BR128_0/RESET vccd1 BR64_1/C[0] BR64_1/C[1] BR64_1/C[2] BR64_1/C[3] BR64_1/C[4]
+ BR64_1/C[5] BR64_1/C[7] BR64_1/C[8] BR64_1/C[9] BR64_1/C[10] BR64_1/C[11] BR64_1/C[12]
+ BR64_1/C[13] BR64_1/C[14] BR64_1/C[15] BR64_1/C[16] BR64_1/C[17] BR64_1/C[18] BR64_1/C[19]
+ BR64_1/C[20] BR64_1/C[21] BR64_1/C[22] BR64_1/C[23] BR64_1/C[24] BR64_1/C[25] BR64_1/C[26]
+ BR64_1/C[27] BR64_1/C[28] BR64_1/C[29] BR64_1/C[30] BR64_1/C[6] BR64_1/C[31] BR64_1/C[32]
+ BR64_1/C[33] BR64_1/C[34] BR64_1/C[35] BR64_1/C[36] BR64_1/C[37] BR64_1/C[38] BR64_1/C[39]
+ BR64_1/C[40] BR64_1/C[41] BR64_1/C[42] BR64_1/C[43] BR64_1/C[44] BR64_1/C[45] BR64_1/C[46]
+ BR64_1/C[47] BR64_1/C[48] BR64_1/C[49] BR64_1/C[50] BR64_1/C[51] BR64_1/C[52] BR64_1/C[53]
+ BR64_1/C[54] BR64_1/C[55] BR64_1/C[56] BR64_1/C[57] BR64_1/C[58] BR64_1/C[59] BR64_1/C[60]
+ BR64_1/C[61] BR64_1/C[62] BR128_1/C[95] BR128_1/C[96] BR128_1/C[97] BR128_1/C[98]
+ BR128_1/C[99] BR128_1/C[100] BR128_1/C[101] BR128_1/C[102] BR128_1/C[103] BR128_1/C[104]
+ BR128_1/C[105] BR128_1/C[106] BR128_1/C[107] BR128_1/C[108] BR128_1/C[109] BR128_1/C[110]
+ BR128_1/C[111] BR128_1/C[112] BR128_0/C[113] BR128_0/C[114] BR128_1/C[115] BR128_1/C[116]
+ BR128_1/C[117] BR128_1/C[118] BR128_1/C[119] BR128_0/C[120] BR128_0/C[121] BR128_1/C[122]
+ BR128_0/C[123] BR128_0/C[124] BR128_0/C[125] BR128_0/C[126] so BR64_1/C[63] BR128_1/C[64]
+ BR128_1/C[65] BR128_0/C[66] BR128_0/C[67] BR128_0/C[68] BR128_1/C[69] BR128_1/C[70]
+ BR128_1/C[71] BR128_1/C[72] BR128_1/C[73] BR128_1/C[74] BR128_1/C[75] BR128_1/C[76]
+ BR128_1/C[77] BR128_1/C[78] BR128_1/C[79] BR128_1/C[80] BR128_1/C[81] BR128_1/C[82]
+ BR128_1/C[83] BR128_1/C[84] BR128_1/C[85] BR128_1/C[86] BR128_1/C[87] BR128_1/C[88]
+ BR128_1/C[89] BR128_1/C[90] BR128_1/C[91] BR128_1/C[92] BR128_1/C[93] BR128_1/C[94]
+ BR128_0/OUT vssd1 BR128
Xsky130_fd_sc_hd__decap_12_1690 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5208 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5219 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4507 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4518 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4529 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3806 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3817 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3828 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3839 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__diode_2_0 BR32_0/C[14] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__dfrtp_2_18 NBR128_1/C[109] sky130_fd_sc_hd__clkbuf_4_1/A NBR128_1/C[108]
+ sky130_fd_sc_hd__clkinv_8_5/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_29 NBR128_1/C[98] rstn NBR128_1/C[97] sky130_fd_sc_hd__clkinv_8_5/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkbuf_4_10 BR64_1/C[41] NBR64_1/C[41] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_21 BR128_1/C[80] NBR128_0/C[80] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_32 BR128_1/C[112] sky130_fd_sc_hd__dfrtp_2_15/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_43 BR64_1/C[48] NBR128_1/C[48] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_54 BR64_1/C[31] BR32_0/C[31] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_65 BR128_1/C[81] NBR128_0/C[81] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__dfrtp_2_108 sky130_fd_sc_hd__dfrtp_2_108/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ NBR64_1/C[18] sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_119 sky130_fd_sc_hd__buf_12_2/A sky130_fd_sc_hd__clkbuf_4_1/X
+ BR64_1/C[7] sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_5005 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5016 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5027 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5038 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4304 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5049 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4315 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4326 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4337 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_6 vccd1 vssd1 BR128_1/C[111] NBR128_0/C[111] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_4348 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3603 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3614 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4359 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3625 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3636 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2902 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3647 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2913 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3658 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2924 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2935 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2946 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2957 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2968 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2979 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5550 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5561 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5572 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5583 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5594 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4860 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4871 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4882 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4893 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_509 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1508 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1519 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XNBR32_1 BR32_0/C[31] BR64_1/C[30] NBR64_1/C[29] BR64_1/C[28] BR64_1/C[27] BR64_1/C[26]
+ NBR64_1/C[25] BR64_1/C[24] NBR64_1/C[23] NBR64_1/C[22] NBR64_1/C[21] NBR64_1/C[20]
+ NBR64_1/C[19] NBR64_1/C[18] NBR64_1/C[17] BR32_0/C[16] NBR64_1/C[15] BR32_0/C[14]
+ NBR32_1/C[13] NBR32_1/C[12] BR64_1/C[11] BR64_1/C[10] BR64_1/C[9] BR64_1/C[8] BR64_1/C[7]
+ BR64_1/C[6] BR32_0/C[5] BR64_1/C[4] BR32_0/C[3] BR64_1/C[2] NBR32_1/C[1] BR64_1/C[0]
+ NBR32_1/RESET NBR32_1/OUT vccd1 vssd1 NBR32
Xsky130_fd_sc_hd__decap_12_4101 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4112 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4123 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4134 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4145 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3400 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3411 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4156 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3422 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4167 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3433 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4178 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3444 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4189 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2710 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3455 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2721 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3466 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2732 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3477 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3488 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2743 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3499 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2754 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2765 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2776 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2787 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2798 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_11 vssd1 vccd1 BR128_1/C[114] BR128_0/C[114] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_5380 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5391 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4690 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_0 sky130_fd_sc_hd__buf_12_0/A BR64_1/C[11] vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_306 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_317 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_328 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_339 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2006 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2017 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2028 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2039 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1305 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1316 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1327 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1338 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1349 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_840 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_851 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_862 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_873 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_884 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_895 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3230 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3241 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3252 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3263 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3274 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2540 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3285 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2551 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3296 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2562 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2573 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2584 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1850 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2595 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1861 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1872 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1883 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1894 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_103 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_114 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_125 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_136 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_147 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_158 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_169 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1102 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1113 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1124 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1135 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1146 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1157 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1168 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1179 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_670 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_681 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_692 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3060 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3071 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3082 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3093 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2370 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2381 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2392 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR128_1 BR128_1/RESET vccd1 BR64_1/C[0] BR64_1/C[1] BR64_1/C[2] BR64_1/C[3] BR64_1/C[4]
+ BR64_1/C[5] BR64_1/C[7] BR64_1/C[8] BR64_1/C[9] BR64_1/C[10] BR64_1/C[11] BR64_1/C[12]
+ BR64_1/C[13] BR64_1/C[14] BR64_1/C[15] BR64_1/C[16] BR64_1/C[17] BR64_1/C[18] BR64_1/C[19]
+ BR64_1/C[20] BR64_1/C[21] BR64_1/C[22] BR64_1/C[23] BR64_1/C[24] BR64_1/C[25] BR64_1/C[26]
+ BR64_1/C[27] BR64_1/C[28] BR64_1/C[29] BR64_1/C[30] BR64_1/C[6] BR64_1/C[31] BR64_1/C[32]
+ BR64_1/C[33] BR64_1/C[34] BR64_1/C[35] BR64_1/C[36] BR64_1/C[37] BR64_1/C[38] BR64_1/C[39]
+ BR64_1/C[40] BR64_1/C[41] BR64_1/C[42] BR64_1/C[43] BR64_1/C[44] BR64_1/C[45] BR64_1/C[46]
+ BR64_1/C[47] BR64_1/C[48] BR64_1/C[49] BR64_1/C[50] BR64_1/C[51] BR64_1/C[52] BR64_1/C[53]
+ BR64_1/C[54] BR64_1/C[55] BR64_1/C[56] BR64_1/C[57] BR64_1/C[58] BR64_1/C[59] BR64_1/C[60]
+ BR64_1/C[61] BR64_1/C[62] BR128_1/C[95] BR128_1/C[96] BR128_1/C[97] BR128_1/C[98]
+ BR128_1/C[99] BR128_1/C[100] BR128_1/C[101] BR128_1/C[102] BR128_1/C[103] BR128_1/C[104]
+ BR128_1/C[105] BR128_1/C[106] BR128_1/C[107] BR128_1/C[108] BR128_1/C[109] BR128_1/C[110]
+ BR128_1/C[111] BR128_1/C[112] BR128_1/C[113] BR128_1/C[114] BR128_1/C[115] BR128_1/C[116]
+ BR128_1/C[117] BR128_1/C[118] BR128_1/C[119] BR128_1/C[120] BR128_1/C[121] BR128_1/C[122]
+ BR128_1/C[123] BR128_1/C[124] BR128_1/C[125] BR128_1/C[126] so BR64_1/C[63] BR128_1/C[64]
+ BR128_1/C[65] BR128_1/C[66] BR128_1/C[67] BR128_1/C[68] BR128_1/C[69] BR128_1/C[70]
+ BR128_1/C[71] BR128_1/C[72] BR128_1/C[73] BR128_1/C[74] BR128_1/C[75] BR128_1/C[76]
+ BR128_1/C[77] BR128_1/C[78] BR128_1/C[79] BR128_1/C[80] BR128_1/C[81] BR128_1/C[82]
+ BR128_1/C[83] BR128_1/C[84] BR128_1/C[85] BR128_1/C[86] BR128_1/C[87] BR128_1/C[88]
+ BR128_1/C[89] BR128_1/C[90] BR128_1/C[91] BR128_1/C[92] BR128_1/C[93] BR128_1/C[94]
+ BR128_1/OUT vssd1 BR128
Xsky130_fd_sc_hd__decap_12_1680 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1691 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4508 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4519 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3807 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3818 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3829 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__diode_2_1 BR128_0/C[120] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__dfrtp_2_19 NBR128_1/C[108] sky130_fd_sc_hd__clkbuf_4_1/A BR128_1/C[107]
+ sky130_fd_sc_hd__clkinv_8_5/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkbuf_4_11 BR64_1/C[36] NBR64_1/C[36] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_22 BR128_1/C[77] NBR128_0/C[77] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_33 BR128_1/C[118] sky130_fd_sc_hd__dfrtp_2_9/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_44 BR64_1/C[46] NBR64_1/C[46] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_55 BR64_1/C[23] NBR64_1/C[23] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_66 BR128_1/C[78] NBR128_0/C[78] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__dfrtp_2_109 NBR64_1/C[18] sky130_fd_sc_hd__clkbuf_4_1/X NBR64_1/C[17]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_5006 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5017 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5028 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5039 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4305 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4316 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4327 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4338 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_7 vccd1 vssd1 BR128_1/C[110] NBR128_1/C[110] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_3604 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4349 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3615 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3626 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3637 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3648 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2903 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2914 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3659 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2925 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2936 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2947 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2958 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2969 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5540 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5551 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5562 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5573 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5584 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4850 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5595 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4861 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4872 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4883 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4894 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1509 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4102 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4113 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4124 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4135 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3401 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4146 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3412 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4157 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3423 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4168 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3434 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4179 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2700 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3445 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3456 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2711 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2722 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3467 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2733 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3478 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2744 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3489 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2755 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2766 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2777 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2788 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2799 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_12 vssd1 vccd1 BR128_1/C[126] BR128_0/C[126] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_5370 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5381 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5392 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4680 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4691 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3990 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_1 sky130_fd_sc_hd__buf_12_1/A BR64_1/C[10] vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_307 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_318 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_329 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2007 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2018 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2029 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1306 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1317 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1328 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1339 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_830 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_841 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_852 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_863 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_874 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_885 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_896 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3220 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3231 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3242 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3253 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3264 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2530 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3275 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2541 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3286 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2552 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3297 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2563 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2574 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1840 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2585 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1851 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2596 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1862 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1873 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1884 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1895 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_0 NBR128_1/C[127] sky130_fd_sc_hd__clkbuf_4_1/X BR128_0/C[126]
+ sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_104 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_115 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_126 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_137 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_148 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_159 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1103 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1114 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1125 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1136 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1147 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1158 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1169 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_660 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_671 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_682 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_693 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3050 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3061 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3072 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3083 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3094 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2360 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2371 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2382 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2393 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1670 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1681 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1692 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_490 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2190 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4509 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3808 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3819 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_12 BR64_1/C[35] NBR64_1/C[35] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_23 BR128_1/C[89] sky130_fd_sc_hd__dfrtp_2_38/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_34 BR128_1/C[122] sky130_fd_sc_hd__dfrtp_2_5/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_45 BR64_1/C[45] NBR64_1/C[45] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_56 BR64_1/C[21] NBR64_1/C[21] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_67 BR128_1/C[86] NBR128_0/C[86] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_5007 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5018 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5029 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4306 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4317 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4328 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4339 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_8 vccd1 vssd1 BR128_1/C[109] NBR128_1/C[109] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_3605 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3616 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3627 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3638 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2904 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3649 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2915 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2926 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2937 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2948 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2959 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5530 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5541 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5552 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5563 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5574 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4840 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5585 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4851 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5596 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4862 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4873 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4884 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4895 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4103 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4114 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4125 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4136 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4147 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3402 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3413 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4158 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3424 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4169 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3435 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2701 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3446 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2712 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3457 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2723 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3468 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2734 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3479 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2745 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2756 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2767 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2778 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2789 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_13 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_1/A2 sky130_fd_sc_hd__o21ai_2_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_5360 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5371 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5382 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5393 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4670 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4681 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4692 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3980 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3991 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_12_2 sky130_fd_sc_hd__buf_12_2/A BR64_1/C[8] vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_308 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_319 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2008 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2019 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1307 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1318 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1329 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_820 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_831 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_842 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_853 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_864 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_875 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_886 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_897 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3210 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3232 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3243 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3254 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2520 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3265 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2531 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3276 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2542 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3287 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2553 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3298 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2564 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1830 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2575 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1841 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2586 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1852 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2597 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1863 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1874 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1885 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1896 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5190 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_1 BR128_0/C[126] sky130_fd_sc_hd__clkbuf_4_1/X BR128_0/C[125]
+ sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_105 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_116 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_127 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_138 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_149 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1104 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1115 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1126 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1137 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1148 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1159 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_650 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_661 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_672 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_683 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_694 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3040 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3051 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3062 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3073 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3084 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2350 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3095 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2361 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2372 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2383 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2394 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1660 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1671 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1682 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1693 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_6 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_480 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_491 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2180 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2191 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1490 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_30 vccd1 vssd1 BR64_1/C[60] NBR64_1/C[60] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_3809 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_13 BR64_1/C[32] NBR64_1/C[32] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_24 BR128_1/C[90] sky130_fd_sc_hd__dfrtp_2_37/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_35 BR128_1/C[119] sky130_fd_sc_hd__dfrtp_2_8/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_46 BR64_1/C[44] NBR64_1/C[44] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_57 BR64_1/C[19] NBR64_1/C[19] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_68 BR128_1/C[87] NBR128_0/C[87] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_6_0 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_12_5008 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5019 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4307 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4318 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4329 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_9 vccd1 vssd1 BR128_1/C[108] NBR128_1/C[108] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_3606 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3628 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3639 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2905 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2916 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2927 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2938 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2949 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5520 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5531 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5542 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5553 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5564 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4830 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5575 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4841 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5586 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4852 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5597 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4863 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4874 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4885 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4896 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4104 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4115 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4126 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4137 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3403 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4148 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3414 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4159 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3425 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3436 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3447 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2702 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3458 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2713 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2724 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3469 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2735 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2746 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2757 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2768 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2779 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_14 vssd1 vccd1 out sky130_fd_sc_hd__o22ai_1_0/Y vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_5350 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5361 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5372 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5383 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5394 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4660 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4671 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4682 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4693 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3970 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3981 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3992 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_309 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2009 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1308 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1319 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_810 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_821 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_832 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_843 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_854 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_865 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_876 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_887 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_898 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3200 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3211 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3222 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3233 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3244 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3255 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2510 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2521 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3266 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2532 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3277 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2543 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3288 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2554 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3299 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1820 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2565 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1831 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2576 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1842 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2587 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1853 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2598 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1864 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1875 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1886 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1897 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5180 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5191 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4490 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_2 BR128_0/C[125] sky130_fd_sc_hd__clkbuf_4_1/X BR128_0/C[124]
+ sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_106 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_117 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_128 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_139 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1105 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1116 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1127 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1138 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1149 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_640 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_651 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_662 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_684 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_695 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3030 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3041 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3052 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3063 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3074 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2340 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3085 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2351 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3096 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2362 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2373 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2384 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1650 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2395 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1661 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1672 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1683 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1694 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_7 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_470 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_481 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_492 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2170 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2181 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2192 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1480 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1491 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_20 vccd1 vssd1 BR128_1/C[96] NBR128_1/C[96] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_31 vccd1 vssd1 BR64_1/C[33] NBR64_1/C[33] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__clkbuf_4_14 BR64_1/C[29] NBR64_1/C[29] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_25 BR128_1/C[73] sky130_fd_sc_hd__dfrtp_2_54/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_36 BR128_1/C[115] sky130_fd_sc_hd__dfrtp_2_12/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_47 BR64_1/C[43] NBR64_1/C[43] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_58 BR64_1/C[18] NBR128_1/C[18] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_69 BR128_1/C[76] NBR128_0/C[76] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_5009 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4308 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4319 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3607 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3618 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2906 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2917 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2928 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2939 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5510 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5521 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5532 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5543 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5554 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4820 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5565 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4831 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5576 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4842 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5587 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4853 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5598 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4864 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4875 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4886 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4897 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4105 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4116 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4127 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4138 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3404 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4149 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3415 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3426 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3437 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2703 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3448 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2714 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3459 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2725 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2736 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2747 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2758 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2769 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_15 vssd1 vccd1 NBR128_1/C[18] NBR64_1/C[18] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_5340 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5351 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5362 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5373 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5384 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4650 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5395 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4661 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4672 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4683 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4694 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3960 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3971 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3982 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3993 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1309 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_800 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_811 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_822 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_833 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_844 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_855 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_866 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_877 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_888 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_899 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3201 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3212 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3223 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3234 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2500 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3245 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2511 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3256 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2522 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3267 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2533 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3278 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2544 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3289 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1810 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2555 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2566 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1821 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1832 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2577 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1843 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2588 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1854 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2599 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1865 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1876 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1887 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1898 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5170 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5181 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5192 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4480 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4491 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3790 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_3 BR128_0/C[124] sky130_fd_sc_hd__clkbuf_4_1/X BR128_0/C[123]
+ sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_107 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_118 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_129 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1106 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1117 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1128 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1139 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_630 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_652 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_663 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_674 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_696 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3020 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3031 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3042 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3053 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3064 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2330 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3075 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2341 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3086 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3097 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2352 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2363 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2374 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2385 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1640 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1651 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2396 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1662 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1684 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1695 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_8 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_460 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_471 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_482 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_493 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2160 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2171 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2182 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2193 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1470 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1481 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1492 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_10 vccd1 vssd1 BR128_1/C[106] NBR128_1/C[106] vssd1 vccd1
+ sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_21 vccd1 vssd1 BR128_1/C[95] NBR128_1/C[95] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_32 vccd1 vssd1 BR32_1/C[13] NBR32_1/C[13] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__clkbuf_4_15 BR64_1/C[25] NBR64_1/C[25] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_26 BR128_1/C[72] sky130_fd_sc_hd__dfrtp_2_55/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_37 sky130_fd_sc_hd__nor2_1_5/A length1 vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_48 BR64_1/C[42] NBR64_1/C[42] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_59 BR64_1/C[17] NBR64_1/C[17] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_290 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4309 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3608 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3619 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2907 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2918 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2929 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5500 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5511 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5522 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5533 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5544 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4810 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5555 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4821 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5566 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4832 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5577 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4843 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5588 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4854 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5599 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4865 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4876 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4887 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4898 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4106 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4117 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4128 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4139 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3405 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3416 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3427 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3438 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3449 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2704 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2715 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2726 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2737 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2748 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2759 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_16 vssd1 vccd1 NBR128_1/C[48] NBR64_1/C[48] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_5330 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5341 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5352 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5363 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5374 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4640 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5385 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4651 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5396 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4662 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4684 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3950 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4695 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3961 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3972 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3983 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3994 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_801 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_812 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_823 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_834 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_845 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_856 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_867 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_878 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_889 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3202 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3213 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3224 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3235 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3246 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2501 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3257 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2512 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2523 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3268 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2534 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3279 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1800 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2545 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1811 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2556 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1822 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2567 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1833 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2578 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1844 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2589 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1855 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1866 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1877 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1888 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1899 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5160 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5171 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5182 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5193 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4470 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4481 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4492 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3780 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3791 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_4 BR128_0/C[123] sky130_fd_sc_hd__clkbuf_4_1/X BR128_1/C[122]
+ sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_108 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_119 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1107 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1118 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1129 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_620 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_631 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_642 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_653 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_664 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_675 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_686 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3010 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3021 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3032 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3043 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3054 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2320 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3065 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2331 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3076 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2342 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3087 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2353 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3098 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2364 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1630 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2375 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2386 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1652 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2397 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1663 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1674 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1696 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_450 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_461 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_472 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_483 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_494 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2150 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2161 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2172 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2183 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2194 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1460 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1471 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1482 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1493 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_11 vccd1 vssd1 BR128_1/C[105] NBR128_1/C[105] vssd1 vccd1
+ sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_22 vccd1 vssd1 BR128_1/C[94] NBR128_1/C[94] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__clkbuf_4_16 BR64_1/C[22] NBR64_1/C[22] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_27 BR128_1/C[91] sky130_fd_sc_hd__dfrtp_2_36/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_38 sky130_fd_sc_hd__nand2_1_8/A length0 vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_49 BR64_1/C[40] NBR64_1/C[40] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_280 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_291 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1290 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3609 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2b_1_0 NBR128_0/RESET sky130_fd_sc_hd__nor2_1_2/B length1 vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__decap_12_2908 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2919 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5501 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5512 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5523 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5534 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4800 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5545 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4811 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5556 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4822 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5567 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4833 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5578 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4844 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5589 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4855 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4866 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4877 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4888 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4899 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_0 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_4107 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4118 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4129 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3406 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3417 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3428 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3439 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2705 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2716 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2727 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2738 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2749 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_17 vssd1 vccd1 BR128_0/C[68] NBR128_1/C[68] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_5320 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5331 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5342 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5353 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5364 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4630 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5375 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5386 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4652 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5397 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4663 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4674 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3940 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3951 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4696 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3962 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3973 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3984 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3995 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_802 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_813 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_824 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_835 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_846 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_857 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_868 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_879 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3203 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3214 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3225 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3236 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2502 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3247 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2513 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3258 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2524 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3269 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2535 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1801 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2546 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1812 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1823 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2568 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1834 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2579 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1845 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1856 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1867 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1878 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1889 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5150 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5161 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5172 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5183 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5194 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4460 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4471 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4482 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4493 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3770 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3781 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3792 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_5 sky130_fd_sc_hd__dfrtp_2_5/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_0/C[121] sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_109 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1108 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1119 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_610 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_621 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_632 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_643 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_654 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_665 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_676 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_687 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_698 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3000 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3011 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3022 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3033 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3044 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2310 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3055 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2321 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3066 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2332 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3077 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3088 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2343 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3099 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2354 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1620 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2365 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1631 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2376 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1642 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2387 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1653 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2398 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1664 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1675 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1686 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4290 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_440 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_451 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_462 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_473 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_484 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_495 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2140 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2151 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2162 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2173 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2184 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1450 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2195 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1461 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1472 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1483 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1494 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_12 vccd1 vssd1 BR128_1/C[104] NBR128_1/C[104] vssd1 vccd1
+ sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_23 vccd1 vssd1 BR128_1/C[93] NBR128_1/C[93] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__clkbuf_4_17 BR64_1/C[20] NBR64_1/C[20] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_28 BR128_1/C[70] sky130_fd_sc_hd__dfrtp_2_57/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_39 BR64_1/C[57] NBR64_1/C[57] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_270 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_281 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_292 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1280 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1291 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2b_1_1 NBR128_1/RESET sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__decap_12_2909 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5502 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5513 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5524 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5535 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4801 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5546 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4812 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4823 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5568 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4834 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5579 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4845 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4856 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4867 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4878 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4889 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4108 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4119 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3407 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3418 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3429 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2706 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2717 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2728 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2739 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5310 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5321 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5332 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5343 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5354 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4620 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5365 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4631 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5376 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4642 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5387 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4653 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5398 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4664 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3930 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4675 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3941 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4686 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3952 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3963 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3974 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3985 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3996 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_803 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_814 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_825 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_836 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_847 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_858 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_869 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3204 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3215 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3226 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3237 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3248 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2503 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3259 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2514 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2525 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2536 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1802 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2547 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1813 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2558 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1824 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2569 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1835 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1846 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1857 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1868 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1879 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5140 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5151 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5162 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5173 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5184 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4450 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5195 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4461 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4472 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4483 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4494 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3760 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3771 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3782 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3793 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_6 BR128_0/C[121] sky130_fd_sc_hd__clkbuf_4_1/X BR128_0/C[120]
+ sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1109 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_600 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_611 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_622 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_633 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_644 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_655 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_666 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_677 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_688 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_699 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3001 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3012 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3023 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3034 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2300 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3045 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3056 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2311 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2322 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3067 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2333 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3078 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2344 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3089 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1610 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2355 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1621 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2366 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1632 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2377 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1643 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2388 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1654 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2399 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1665 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1676 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1687 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1698 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4280 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4291 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3590 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_430 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_441 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_452 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_463 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_474 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_485 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_496 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2130 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2141 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2152 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2163 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2174 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1440 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2185 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1451 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2196 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1462 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1473 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1484 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1495 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_13 vccd1 vssd1 BR128_1/C[103] NBR128_1/C[103] vssd1 vccd1
+ sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_24 vccd1 vssd1 BR128_1/C[92] NBR128_1/C[92] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__clkbuf_4_18 BR128_1/C[82] NBR128_0/C[82] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_29 BR128_1/C[71] sky130_fd_sc_hd__dfrtp_2_56/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_260 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_271 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_282 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_293 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1270 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1281 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1292 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2b_1_2 BR128_0/RESET sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__nor2_1_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__decap_12_5503 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5514 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5525 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5536 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4802 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5547 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4813 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5558 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4824 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5569 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4835 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4846 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4857 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4868 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4879 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4109 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3408 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3419 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2707 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2718 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2729 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5300 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5311 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5322 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5333 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5344 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4610 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5355 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4621 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5366 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4632 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5377 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4643 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5388 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4654 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5399 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3920 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4665 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4676 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3931 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3942 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4687 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3953 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4698 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3964 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3975 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3986 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3997 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_804 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_815 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_826 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_837 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_848 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_859 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3205 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3216 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3227 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3238 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2504 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3249 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2515 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2526 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2537 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1803 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2548 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2559 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1814 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1825 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1836 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1847 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1858 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1869 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5130 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5141 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5152 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5163 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5174 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4440 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5185 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5196 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4451 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4462 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4473 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4484 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3750 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4495 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3761 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3772 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3783 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3794 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_7 BR128_0/C[120] sky130_fd_sc_hd__clkbuf_4_1/X BR128_1/C[119]
+ sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_612 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_623 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_634 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_656 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_667 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_678 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_689 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3002 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3013 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3024 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3035 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2301 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3046 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2312 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3057 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2323 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3068 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2334 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3079 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1600 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2345 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1611 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2356 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1622 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2367 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1633 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2378 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1644 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2389 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1655 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1666 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1677 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1688 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_0 sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__nand2_1_2/B
+ sky130_fd_sc_hd__nor2_1_0/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1699 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4270 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4281 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4292 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3580 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3591 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2890 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_420 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_431 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_442 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_453 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_464 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_475 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_486 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_497 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2120 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2131 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2142 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2153 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2164 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1430 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2175 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1441 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2186 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1452 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2197 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1463 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1474 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1485 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1496 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_14 vccd1 vssd1 BR128_1/C[102] NBR128_1/C[102] vssd1 vccd1
+ sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_25 vccd1 vssd1 BR128_1/C[65] NBR128_1/C[65] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__clkbuf_4_19 BR128_1/C[83] NBR128_0/C[83] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_250 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_261 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_272 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_283 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_294 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1260 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1271 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1282 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1293 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2b_1_3 BR128_1/RESET sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__nor2_1_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__decap_12_5504 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5515 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5526 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5537 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4803 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5548 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4814 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5559 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4825 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4836 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4847 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4858 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4869 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1090 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3409 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2708 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2719 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5301 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5312 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5323 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5334 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5345 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4600 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5356 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4611 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4622 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5367 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4633 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5378 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4644 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5389 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3910 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4655 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3921 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4666 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3932 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4677 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3943 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4688 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4699 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3954 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3965 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3976 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3987 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3998 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_805 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_816 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_827 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_838 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_849 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3206 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3217 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3228 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3239 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2505 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2516 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2527 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2538 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1804 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2549 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1815 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1826 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1837 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1848 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1859 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5120 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5131 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5142 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5153 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5164 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4430 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5175 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4441 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5186 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4452 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5197 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4463 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4474 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3740 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4485 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3751 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4496 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3762 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3773 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3784 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3795 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_8 sky130_fd_sc_hd__dfrtp_2_8/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_1/C[118] sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_602 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_624 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_635 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_646 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_668 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_679 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3003 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3014 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3025 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3036 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2302 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3047 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3058 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2313 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2324 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3069 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2335 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2346 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1612 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2357 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1623 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2368 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1634 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2379 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1656 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1667 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1678 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1689 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_1 sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__nor2_1_0/Y
+ puf_sel0 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_4260 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4271 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4282 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4293 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3570 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3581 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3592 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2880 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2891 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_90 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_410 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_421 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_432 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_443 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_454 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_465 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_476 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_487 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_498 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2110 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2121 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2132 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2143 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2154 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1420 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2165 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1431 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2176 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1442 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2187 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1453 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2198 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1464 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1475 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1486 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1497 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_15 vccd1 vssd1 BR128_1/C[101] NBR128_1/C[101] vssd1 vccd1
+ sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_26 vccd1 vssd1 BR128_1/C[64] NBR128_1/C[64] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_4090 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_2_0 sky130_fd_sc_hd__nand2_1_6/Y sky130_fd_sc_hd__o21ai_2_0/Y
+ sky130_fd_sc_hd__nor2_1_5/A sky130_fd_sc_hd__o22ai_1_4/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__decap_12_240 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_251 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_262 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_273 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_284 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_295 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1250 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1261 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1272 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1283 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1294 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_0 vssd1 vccd1 NBR64_0/C[18] NBR64_1/C[18] vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_5505 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5516 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5527 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5538 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4804 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5549 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4815 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4826 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4837 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4848 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4859 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_0 sky130_fd_sc_hd__nand2_1_2/B puf_sel0 vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1080 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1091 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2709 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5302 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5313 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5324 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5335 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5346 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4612 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5357 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4623 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5368 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4634 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5379 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3900 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3911 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4656 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3922 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4667 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3933 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4678 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3944 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4689 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3955 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3966 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3977 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3988 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3999 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_806 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_817 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_828 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_839 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3207 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3218 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3229 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2506 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2517 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2528 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2539 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1805 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1816 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1827 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1838 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1849 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5110 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5121 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5132 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5143 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5154 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4420 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5165 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4431 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5176 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4442 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5187 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5198 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4453 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4464 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4475 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3730 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3741 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4486 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3752 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4497 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3763 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3774 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3785 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3796 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_9 sky130_fd_sc_hd__dfrtp_2_9/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ NBR128_0/C[117] sky130_fd_sc_hd__clkinv_8_9/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_603 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_614 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_625 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_636 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_647 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_658 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3004 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3015 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3026 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3037 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2303 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3048 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2314 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3059 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2325 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2336 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1602 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2347 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2358 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1624 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2369 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1635 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1646 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1668 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1679 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_2 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nand2_1_2/B
+ sky130_fd_sc_hd__nor2_1_1/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_4250 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4261 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4272 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4283 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4294 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3560 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3571 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3582 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3593 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2870 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2881 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2892 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_80 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_91 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_400 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_411 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_422 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_433 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_444 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_455 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_466 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_477 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_488 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_499 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2100 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2111 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2122 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2133 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2144 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1410 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2155 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1421 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2166 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1432 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2177 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1443 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2188 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1454 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2199 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1465 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1476 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1487 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1498 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_16 vccd1 vssd1 BR128_1/C[100] NBR128_1/C[100] vssd1 vccd1
+ sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_27 vccd1 vssd1 BR64_1/C[63] NBR64_1/C[63] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_4080 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4091 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3390 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_230 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_241 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_252 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_263 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_274 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_285 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_296 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1240 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1251 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1262 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1273 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1284 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1295 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_1 vssd1 vccd1 NBR64_0/C[17] NBR64_1/C[17] vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_5506 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5517 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5528 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5539 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4805 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4816 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4827 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4838 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4849 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_1 sky130_fd_sc_hd__nor2_1_1/B puf_sel1 vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1070 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1081 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1092 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5303 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5314 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5325 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5336 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5347 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4602 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5358 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4624 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5369 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4635 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3901 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4646 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3912 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3923 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4668 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3934 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4679 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3945 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3956 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3967 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3978 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3989 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_807 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_818 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_829 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3208 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3219 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2507 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2518 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2529 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1806 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1817 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1828 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1839 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5100 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5111 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5122 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5133 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5144 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5155 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4410 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5166 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4421 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4432 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5177 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4443 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5188 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4454 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5199 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3720 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4465 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3731 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4476 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3742 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4487 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3753 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4498 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3764 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3775 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3786 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3797 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_604 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_615 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_626 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_637 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_648 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_659 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3005 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3016 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3027 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3038 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2304 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3049 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2315 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2326 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2337 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1603 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2348 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1614 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2359 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1625 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1636 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1647 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1658 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_3 sky130_fd_sc_hd__nand2_1_3/Y NBR128_0/OUT length1 vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_4240 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4251 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4262 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4273 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4284 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3550 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4295 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3561 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3572 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3583 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3594 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2860 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2871 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2882 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2893 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_70 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_81 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_92 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_401 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_412 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_423 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_434 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_445 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_456 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_467 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_478 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_489 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2101 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2112 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2123 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2134 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1400 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2145 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1411 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2156 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1422 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2167 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1433 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2178 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1444 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2189 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1455 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1466 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1477 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1488 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1499 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_17 vccd1 vssd1 BR128_1/C[99] NBR128_1/C[99] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_28 vccd1 vssd1 BR64_1/C[62] NBR64_1/C[62] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_990 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4070 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4081 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4092 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3380 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3391 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2690 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_220 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_231 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_242 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_253 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_264 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_275 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_286 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_297 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1230 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1241 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1252 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1263 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1274 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1285 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1296 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_2 vssd1 vccd1 BR128_1/C[67] BR128_0/C[67] vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_5507 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5518 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5529 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4806 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4817 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4828 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4839 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_2 sky130_fd_sc_hd__nand2_1_4/B length0 vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1060 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1071 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1082 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1093 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5304 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5315 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5326 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5337 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4603 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5348 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4614 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5359 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4625 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4636 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3902 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4647 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3913 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4658 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3924 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3935 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3946 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3957 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3968 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3979 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_808 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_819 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2508 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2519 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1807 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1818 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1829 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5101 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5112 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5123 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5134 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4400 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5145 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4411 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5156 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4422 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5167 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4433 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5178 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5189 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4444 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3710 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4455 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3721 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4466 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4477 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3732 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3743 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4488 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3754 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4499 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3765 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3776 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3787 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3798 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_605 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_616 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_627 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_638 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_649 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3006 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3017 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3028 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3039 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2305 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2316 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2327 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2338 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1604 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2349 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1615 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1626 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1637 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1648 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1659 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_4 NBR32_0/RESET sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nor2_1_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_4230 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4241 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4252 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4263 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4274 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4285 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3540 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3551 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4296 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3562 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3573 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3584 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2850 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3595 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2861 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2872 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2883 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2894 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_60 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_71 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_82 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_93 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_402 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_413 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_424 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_435 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_446 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_457 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_468 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_479 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2102 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2113 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2124 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2135 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1401 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2146 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1412 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2157 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1423 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2168 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1434 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2179 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1445 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1456 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1467 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1478 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1489 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_18 vccd1 vssd1 BR128_1/C[98] NBR128_1/C[98] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_29 vccd1 vssd1 BR64_1/C[61] NBR64_1/C[61] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_980 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_991 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4060 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4071 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4082 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4093 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3370 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3381 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3392 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2680 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2691 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1990 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_210 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_232 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_243 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_254 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_265 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_276 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_287 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_298 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1220 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1231 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1242 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1253 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1264 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1275 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1286 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1297 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_3 vssd1 vccd1 BR128_1/C[66] BR128_0/C[66] vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_5508 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5519 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4807 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4818 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4829 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_0_0 vssd1 vccd1 sky130_fd_sc_hd__o21ai_0_0/Y sky130_fd_sc_hd__nand2_1_3/Y
+ length1 sky130_fd_sc_hd__o22ai_1_3/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_0
Xsky130_fd_sc_hd__clkinv_1_3 sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__nand2_1_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1050 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1061 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1072 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1083 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1094 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5305 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5316 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5327 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5338 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5349 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4604 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4615 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4626 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4637 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3903 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4648 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3914 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4659 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3925 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3936 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3947 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3958 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3969 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_809 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2509 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1808 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1819 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5102 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5113 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5124 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5135 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4401 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5146 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5157 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4412 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4423 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5168 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4434 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5179 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3700 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4445 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3711 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4456 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3722 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4467 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3733 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4478 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3744 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4489 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3755 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3766 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3777 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3788 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3799 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4990 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_606 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_628 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_639 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3007 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3018 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3029 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2306 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2317 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2328 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2339 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1605 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1616 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1627 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1638 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1649 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_5 NBR64_0/RESET sky130_fd_sc_hd__nor2_1_2/Y length0 vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_4220 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4231 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4242 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4253 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4264 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3530 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4275 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3541 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4286 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3552 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4297 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3563 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3574 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3585 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2840 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2851 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3596 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2862 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2873 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2884 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2895 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_50 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_61 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_72 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_83 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_94 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_403 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_414 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_425 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_436 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_447 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_458 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_469 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2103 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2114 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2125 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2136 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1402 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2147 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1413 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2158 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1424 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2169 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1435 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1446 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1457 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1468 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1479 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_19 vccd1 vssd1 BR128_1/C[97] NBR128_1/C[97] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_970 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_981 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_992 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4050 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4061 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4072 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4083 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4094 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3360 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3371 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3382 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3393 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2670 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2681 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2692 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1980 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1991 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_200 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_211 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_222 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_233 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_244 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_255 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_266 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_277 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_288 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_299 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1210 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1232 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1243 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1254 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1265 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1276 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1287 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1298 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3190 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_4 vssd1 vccd1 BR32_1/C[14] BR32_0/C[14] vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_5509 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4808 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4819 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_4 sky130_fd_sc_hd__o22ai_1_5/B1 sky130_fd_sc_hd__nand2_1_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1040 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1051 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1062 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1073 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1084 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1095 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5306 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5317 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5328 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5339 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4605 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4616 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4627 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4638 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3904 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4649 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3915 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3926 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3937 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3948 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3959 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1809 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5103 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5114 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5125 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5136 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4402 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5147 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4413 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5158 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4424 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5169 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4435 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3701 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4446 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3712 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4457 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3723 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4468 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3734 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4479 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3745 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3756 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3767 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3778 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3789 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4980 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4991 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_607 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_618 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3008 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3019 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2307 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2318 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2329 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1606 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1628 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1639 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_6 sky130_fd_sc_hd__nand2_1_6/Y NBR128_1/OUT sky130_fd_sc_hd__nor2_1_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_4210 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4232 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4243 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4254 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3520 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4265 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4276 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3531 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3542 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4287 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3553 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4298 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3564 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2830 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3575 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2841 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3586 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2852 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3597 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2863 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2874 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2885 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2896 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_40 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_51 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_62 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_73 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_84 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_95 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_404 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_415 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_426 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_437 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_448 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_459 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2104 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2115 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2126 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2137 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1403 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2148 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1414 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2159 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1425 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1436 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1447 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1458 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1469 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_960 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_971 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_982 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_993 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4040 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4051 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4062 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4073 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4084 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3350 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4095 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3361 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3372 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3383 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3394 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2660 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2671 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2682 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2693 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1970 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1981 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1992 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_201 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_212 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_223 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_234 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_245 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_256 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_267 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_278 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_289 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1200 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1211 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1222 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1233 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1244 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1255 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1266 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1277 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1288 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1299 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_790 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3180 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3191 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2490 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_5 vssd1 vccd1 BR128_1/C[120] BR128_0/C[120] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_4809 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_5 sky130_fd_sc_hd__o22ai_1_6/B1 sky130_fd_sc_hd__nand2_1_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1030 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1041 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1052 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1063 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1074 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1085 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1096 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5307 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5318 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5329 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4606 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4628 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4639 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3905 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3916 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3927 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3938 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3949 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5104 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5115 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5126 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5137 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4403 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5148 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4414 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5159 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4425 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4436 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3702 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4447 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3713 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4458 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3724 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4469 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3735 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3746 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3757 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3768 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3779 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4970 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4981 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4992 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_608 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_619 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3009 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2308 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2319 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1607 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1618 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_7 NBR32_1/RESET sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__nor2_1_3/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_4200 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4211 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4222 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4233 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4244 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3510 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4255 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3521 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4266 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3532 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4277 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3543 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4288 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4299 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3554 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2820 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3565 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3576 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2831 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3587 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2842 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2853 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3598 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2864 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2875 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2886 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2897 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_30 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_41 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_52 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_63 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_74 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_85 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5490 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_96 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_405 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_416 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_427 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_438 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_449 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2105 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2116 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2127 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2138 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1404 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2149 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1415 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1426 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1437 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1448 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1459 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_950 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_961 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_972 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_983 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_994 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4030 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4041 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4052 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4063 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4074 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3340 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4085 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3351 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4096 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3362 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3373 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3384 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2650 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3395 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2661 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2672 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2683 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2694 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1960 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1971 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1982 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1993 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_202 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_213 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_224 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_235 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_246 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_257 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_268 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_279 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1201 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1212 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1223 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1234 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1245 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1256 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1267 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1278 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1289 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_780 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_791 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3170 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3181 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3192 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2480 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2491 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1790 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_6 vssd1 vccd1 BR128_1/C[125] BR128_0/C[125] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_6 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__dfrtp_2_97/Q
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1020 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1031 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1042 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1053 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1064 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1075 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1086 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1097 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5308 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5319 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4607 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4618 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3906 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3917 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3928 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3939 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5105 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5116 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5127 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5138 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4404 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5149 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4415 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4426 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4437 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4448 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3703 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3714 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4459 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3725 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3736 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3747 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3758 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3769 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4960 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4971 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4982 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4993 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_609 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2309 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1608 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1619 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_8 NBR64_1/RESET sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__nand2_1_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_4201 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4212 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4223 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4234 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3500 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4245 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4256 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3511 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3522 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4267 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3533 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4278 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3544 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4289 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2810 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3555 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2821 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3566 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2832 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3577 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2843 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3588 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2854 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3599 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2865 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2876 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2887 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2898 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_20 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_31 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_42 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_53 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_64 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_75 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5480 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_86 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5491 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_97 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4790 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_406 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_417 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_428 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_439 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2106 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2117 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2128 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2139 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1405 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1416 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1427 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1438 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1449 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_940 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_951 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_962 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_973 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_984 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4020 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_995 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4031 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4042 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4053 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4064 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4075 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3330 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3341 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4086 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3352 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4097 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3363 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3374 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2640 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3385 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2651 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3396 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2662 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2684 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1950 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2695 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1961 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1972 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1983 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1994 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_8_0 BR64_1/C[14] BR32_0/C[14] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__decap_12_203 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_214 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_225 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_236 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_247 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_258 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_269 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1202 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1213 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1224 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1235 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1246 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1257 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1268 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1279 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_0 sky130_fd_sc_hd__clkinv_8_8/A sky130_fd_sc_hd__clkinv_8_0/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_770 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_781 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_792 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3160 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3171 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3182 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3193 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
.ends

.subckt sky130_fd_pr__res_generic_m1_DBNWX4 m1_n500_n557# m1_n500_500#
R0 m1_n500_n557# m1_n500_500# sky130_fd_pr__res_generic_m1 w=5e+06u l=5e+06u
.ends

.subckt puf_top m1_44147_10052# puf_super_0/si puf_super_0/length0 puf_super_0/out
+ puf_super_0/clk puf_super_0/reset puf_super_0/puf_sel0 puf_super_0/length1 puf_super_0/puf_sel1
+ puf_super_0/vccd1 puf_super_0/so m1_40740_16650# VSUBS puf_super_0/rstn
Xpuf_super_0 puf_super_0/reset puf_super_0/clk puf_super_0/si puf_super_0/rstn puf_super_0/puf_sel1
+ puf_super_0/puf_sel0 puf_super_0/length1 puf_super_0/length0 puf_super_0/out puf_super_0/so
+ puf_super_0/vccd1 VSUBS puf_super
Xsky130_fd_pr__res_generic_m1_DBNWX4_0 puf_super_0/so m1_40740_16650# sky130_fd_pr__res_generic_m1_DBNWX4
Xsky130_fd_pr__res_generic_m1_DBNWX4_1 puf_super_0/out m1_44147_10052# sky130_fd_pr__res_generic_m1_DBNWX4
.ends

.subckt nmos_flat VPWR SOURCE DRAIN GATE VGND
X0 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X2 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X3 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X4 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X5 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X6 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X7 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X8 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X9 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X10 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X11 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X12 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X13 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X14 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X15 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X16 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X17 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X18 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X19 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__res_generic_m4_LS59QM m4_n4500_n3057# m4_n4500_3000#
R0 m4_n4500_n3057# m4_n4500_3000# sky130_fd_pr__res_generic_m4 w=4.5e+07u l=3e+07u
.ends

.subckt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 Emitter Collector Base m=1
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
.ends

.subckt bandgaptop_flat_io bandgaptop_flat_0/porst bandgaptop_flat_0/VDD bandgaptop_flat_0/GND
+ bandgaptop_flat_0/bandgapcorev3_0/Vbg
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|0] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|0] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|0] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|0] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|0] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5|0] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|0] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|0] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|1] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|1] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|1] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|1] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|1] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5|1] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|1] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|1] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|3] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|3] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|3] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|3] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|3] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5|3] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|3] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|3] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|4] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|4] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|4] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|4] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|4] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5|4] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter
+ bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
X0 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X4 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.156e+13p ps=1.36e+07u w=3.87e+07u l=2e+06u
X5 bandgaptop_flat_0/bandgapcorev3_0/Vb bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X6 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X7 a_463132_642452# bandgaptop_flat_0/bandgapcorev3_0/VbEnd bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X8 bandgaptop_flat_0/amplifier_0/Vx bandgaptop_flat_0/GND bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.5632e+14p ps=1.424e+09u w=2e+06u l=2e+06u
X9 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X10 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X11 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X12 bandgaptop_flat_0/GND bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X13 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X14 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X15 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X16 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X17 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X18 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X19 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X20 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X21 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X22 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X23 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X24 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X25 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X26 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X27 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X28 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X29 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X30 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X31 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X32 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X33 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X34 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X35 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X36 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X37 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X38 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X39 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X40 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X41 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X42 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X43 bandgaptop_flat_0/bandgapcorev3_0/VbgEnd a_463950_649188# bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X44 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X46 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/bandgapcorev3_0/Vb bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X47 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X48 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X49 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X50 bandgaptop_flat_0/GND bandgaptop_flat_0/bandgapcorev3_0/VaEnd bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=2.15e+07u
X51 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X52 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X53 bandgaptop_flat_0/GND bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=2.15e+07u
X54 bandgaptop_flat_0/bandgapcorev3_0/Vb bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X55 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X56 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X57 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X58 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X60 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X61 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X63 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X64 a_468858_642452# a_466404_649188# bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X65 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X66 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X67 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X68 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X69 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X70 bandgaptop_flat_0/GND bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=1.662e+07u
X71 bandgaptop_flat_0/bandgapcorev3_0/Vb a_471312_649188# bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X72 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X73 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X74 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X75 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X76 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X77 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X78 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X79 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X80 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X81 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X82 bandgaptop_flat_0/bandgapcorev3_0/Vb bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X83 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X84 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X85 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X86 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X87 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X88 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X89 a_463132_642452# a_466404_649188# bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X90 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X91 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X92 a_462314_642452# a_464768_649188# bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X93 bandgaptop_flat_0/bandgapcorev3_0/Vbg bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X94 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X95 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X96 bandgaptop_flat_0/bandgapcorev3_0/Vbg bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X97 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X98 a_468858_642452# a_471312_649188# bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X99 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X101 bandgaptop_flat_0/bandgapcorev3_0/Vbg bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X102 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X103 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X104 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X105 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X106 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X107 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X108 bandgaptop_flat_0/amplifier_0/Vq bandgaptop_flat_0/bandgapcorev3_0/Vb bandgaptop_flat_0/amplifier_0/vg bandgaptop_flat_0/GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=9e+06u l=2e+06u
X109 bandgaptop_flat_0/amplifier_0/Vq sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=9e+06u l=2e+06u
X110 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X111 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X115 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X116 bandgaptop_flat_0/GND bandgaptop_flat_0/amplifier_0/Vx bandgaptop_flat_0/amplifier_0/Vq bandgaptop_flat_0/GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X117 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X118 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X119 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X120 bandgaptop_flat_0/GND bandgaptop_flat_0/GND bandgaptop_flat_0/amplifier_0/Vx bandgaptop_flat_0/GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X121 bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X122 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X123 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7|4]/Emitter bandgaptop_flat_0/bandgapcorev3_0/Vb bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X124 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X125 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X126 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X127 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X128 a_462314_642452# bandgaptop_flat_0/bandgapcorev3_0/VaEnd bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X129 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X130 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/amplifier_0/Vx bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.29e+07u l=2e+06u
X131 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X132 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X133 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X134 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X135 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X136 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X137 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/amplifier_0/Vx bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.29e+07u l=2e+06u
X138 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X139 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X140 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X141 bandgaptop_flat_0/amplifier_0/Vq sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=9e+06u l=2e+06u
X142 bandgaptop_flat_0/GND bandgaptop_flat_0/GND bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=9e+06u l=2e+06u
X143 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X144 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X145 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X146 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X147 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X148 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/bandgapcorev3_0/Vbg bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X149 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X150 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X151 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X152 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X153 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X154 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X155 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X156 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X157 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X158 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X159 bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.29e+07u l=2e+06u
X160 bandgaptop_flat_0/amplifier_0/Vq sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=9e+06u l=2e+06u
X161 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X162 bandgaptop_flat_0/amplifier_0/Vq bandgaptop_flat_0/bandgapcorev3_0/Vb bandgaptop_flat_0/amplifier_0/vg bandgaptop_flat_0/GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=9e+06u l=2e+06u
X163 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X164 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X165 bandgaptop_flat_0/amplifier_0/Vx bandgaptop_flat_0/amplifier_0/Vx bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X166 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/bandgapcorev3_0/Vb bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X167 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X168 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X169 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X170 bandgaptop_flat_0/GND bandgaptop_flat_0/bandgapcorev3_0/VbEnd bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=2.15e+07u
X171 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X172 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X173 bandgaptop_flat_0/VDD bandgaptop_flat_0/amplifier_0/vg bandgaptop_flat_0/amplifier_0/vg bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.29e+07u l=2e+06u
X174 bandgaptop_flat_0/VDD bandgaptop_flat_0/amplifier_0/vg bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.29e+07u l=2e+06u
X175 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X176 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X177 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X178 bandgaptop_flat_0/GND bandgaptop_flat_0/GND bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=9e+06u l=2e+06u
X179 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/bandgapcorev3_0/Vbg bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X180 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X181 bandgaptop_flat_0/bandgapcorev3_0/Vbg bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X182 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X183 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X184 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X185 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X186 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X187 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X188 bandgaptop_flat_0/bandgapcorev3_0/Vbg bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X189 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X190 bandgaptop_flat_0/amplifier_0/Vq bandgaptop_flat_0/amplifier_0/Vx bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X191 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X192 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X193 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X194 bandgaptop_flat_0/VDD bandgaptop_flat_0/amplifier_0/vg bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.29e+07u l=2e+06u
X195 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/amplifier_0/Vx bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.29e+07u l=2e+06u
X196 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X197 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X198 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X199 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter a_470494_649188# bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X200 bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.29e+07u l=2e+06u
X201 bandgaptop_flat_0/GND bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=2.15e+07u
X202 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X203 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X204 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X205 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X206 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X207 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X208 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X209 bandgaptop_flat_0/GND bandgaptop_flat_0/porst bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.7e+07u l=2e+06u
X210 bandgaptop_flat_0/GND bandgaptop_flat_0/amplifier_0/Vx bandgaptop_flat_0/amplifier_0/Vx bandgaptop_flat_0/GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=2e+06u
X211 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X212 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X213 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X214 bandgaptop_flat_0/amplifier_0/Vq bandgaptop_flat_0/bandgapcorev3_0/Vb bandgaptop_flat_0/amplifier_0/vg bandgaptop_flat_0/GND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=9e+06u l=2e+06u
X215 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X216 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X217 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X218 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X219 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X220 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X221 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X222 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X223 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X224 a_465586_642452# a_469676_649188# bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X225 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/amplifier_0/Vx bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.29e+07u l=2e+06u
X226 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/amplifier_0/Vx bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.29e+07u l=2e+06u
X227 bandgaptop_flat_0/VDD bandgaptop_flat_0/amplifier_0/vg bandgaptop_flat_0/amplifier_0/vg bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.29e+07u l=2e+06u
X228 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X229 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X230 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X231 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X232 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X233 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X234 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X235 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X236 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X237 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X238 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X239 bandgaptop_flat_0/GND bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X240 bandgaptop_flat_0/bandgapcorev3_0/VbgEnd bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=1.662e+07u
X241 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X242 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X243 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/bandgapcorev3_0/Vb bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X244 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X245 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X246 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X247 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/bandgapcorev3_0/Vbg bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X248 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X249 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/bandgapcorev3_0/Vb bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X250 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X251 bandgaptop_flat_0/bandgapcorev3_0/Vb bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X252 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/amplifier_0/Vx bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.29e+07u l=2e+06u
X253 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X254 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X255 bandgaptop_flat_0/bandgapcorev3_0/Vb bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X256 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X257 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X258 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X259 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X260 a_467222_642452# a_464768_649188# bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X261 bandgaptop_flat_0/VDD bandgaptop_flat_0/amplifier_0/vg bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.29e+07u l=2e+06u
X262 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X263 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X264 a_465586_642452# a_463950_649188# bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X265 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X266 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X267 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X268 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/bandgapcorev3_0/Vb bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X269 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X270 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X271 bandgaptop_flat_0/bandgapcorev3_0/Vbg a_469676_649188# bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X272 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/bandgapcorev3_0/Vbg bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X273 a_467222_642452# a_470494_649188# bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=3.152e+07u
X274 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X275 bandgaptop_flat_0/VDD bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/bandgapcorev3_0/Vbg bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.87e+07u l=2e+06u
X276 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X277 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X278 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X279 bandgaptop_flat_0/GND bandgaptop_flat_0/GND bandgaptop_flat_0/GND sky130_fd_pr__res_xhigh_po_2p85 l=1.662e+07u
X280 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X281 bandgaptop_flat_0/currentmirror_0/Vgate bandgaptop_flat_0/VDD sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X282 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X283 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Emitter bandgaptop_flat_0/GND sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
X284 bandgaptop_flat_0/VDD bandgaptop_flat_0/amplifier_0/vg bandgaptop_flat_0/amplifier_0/vg bandgaptop_flat_0/VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.29e+07u l=2e+06u
.ends

.subckt sky130_asc_res_xhigh_po_2p85_1 Rin Rout VPWR VGND
X0 Rin a_2148_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X1 Rout a_2148_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
.ends

.subckt sky130_asc_pfet_01v8_lvt_60 GATE SOURCE DRAIN VGND VPWR
X0 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X1 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X6 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X7 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X8 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X9 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X10 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X11 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X12 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X13 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X14 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X15 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X16 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X17 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X18 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X19 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X20 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X21 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X22 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X23 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X24 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X25 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X26 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X27 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X28 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X29 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X30 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X31 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X32 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X33 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X34 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X35 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X36 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X37 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X38 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X39 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X40 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X41 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X42 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X43 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X44 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X45 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X46 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X47 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X48 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X49 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X50 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X51 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X52 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X53 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X54 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X55 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X56 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X57 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X58 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X59 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
.ends

.subckt sky130_asc_pnp_05v5_W3p40L3p40_7 Emitter Base Collector VPWR VGND
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X1 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X2 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X3 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X4 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X5 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X6 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
.ends

.subckt sky130_asc_res_xhigh_po_2p85_2 Rin Rout VPWR VGND
X0 Rout a_2723_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
X1 Rin a_2723_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
.ends

.subckt sky130_asc_pfet_01v8_lvt_12 GATE SOURCE DRAIN VGND VPWR
X0 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X1 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X6 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X7 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X8 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X9 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X10 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X11 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
.ends

.subckt sky130_asc_nfet_01v8_lvt_9 GATE SOURCE DRAIN VPWR VGND
X0 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X1 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X8 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
.ends

.subckt sky130_asc_pfet_01v8_lvt_6 GATE SOURCE DRAIN VGND VPWR
X0 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X1 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
.ends

.subckt sky130_asc_pnp_05v5_W3p40L3p40_1 Emitter Base Collector VPWR VGND
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
.ends

.subckt sky130_asc_cap_mim_m3_1 Cin Cout VPWR VGND
X0 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X8 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X9 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X10 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X11 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X12 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X13 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X14 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X15 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X16 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X17 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X18 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X19 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
.ends

.subckt sky130_asc_pnp_05v5_W3p40L3p40_8 Emitter Base Collector VPWR VGND
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X1 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X2 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X3 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X4 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X5 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X6 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X7 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
.ends

.subckt sky130_asc_nfet_01v8_lvt_1 GATE SOURCE DRAIN VPWR VGND
X0 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
.ends

.subckt bgr_gen7 porst vbg VSS VDD
Xsky130_asc_res_xhigh_po_2p85_1_7 vbg sky130_asc_res_xhigh_po_2p85_1_2/Rin VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_8 sky130_asc_res_xhigh_po_2p85_1_8/Rin sky130_asc_res_xhigh_po_2p85_1_1/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_9 sky130_asc_cap_mim_m3_1_9/Cin sky130_asc_res_xhigh_po_2p85_1_9/Rout
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_60_0 sky130_asc_cap_mim_m3_1_4/Cout VDD vbg VSS VDD sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_pfet_01v8_lvt_60_1 sky130_asc_cap_mim_m3_1_4/Cout VDD sky130_asc_nfet_01v8_lvt_9_1/GATE
+ VSS VDD sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_pfet_01v8_lvt_60_2 sky130_asc_cap_mim_m3_1_4/Cout VDD sky130_asc_cap_mim_m3_1_9/Cin
+ VSS VDD sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_res_xhigh_po_2p85_1_30 sky130_asc_res_xhigh_po_2p85_1_30/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_20 sky130_asc_res_xhigh_po_2p85_1_20/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pnp_05v5_W3p40L3p40_7_0 sky130_asc_res_xhigh_po_2p85_1_12/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_7
Xsky130_asc_res_xhigh_po_2p85_1_10 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_2_0/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_21 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_13/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_2_0 sky130_asc_res_xhigh_po_2p85_2_0/Rin VSS VDD VSS
+ sky130_asc_res_xhigh_po_2p85_2
Xsky130_asc_res_xhigh_po_2p85_1_11 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_20/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_22 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_11/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_2_1 sky130_asc_res_xhigh_po_2p85_2_1/Rin VSS VDD VSS
+ sky130_asc_res_xhigh_po_2p85_2
Xsky130_asc_res_xhigh_po_2p85_1_12 sky130_asc_res_xhigh_po_2p85_1_12/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rout
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_23 sky130_asc_res_xhigh_po_2p85_1_23/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_13 sky130_asc_res_xhigh_po_2p85_1_13/Rin sky130_asc_nfet_01v8_lvt_9_1/GATE
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_24 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_28/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_12_0 sky130_asc_cap_mim_m3_1_4/Cout VDD sky130_asc_nfet_01v8_lvt_1_1/GATE
+ VSS VDD sky130_asc_pfet_01v8_lvt_12
Xsky130_asc_res_xhigh_po_2p85_1_14 sky130_asc_nfet_01v8_lvt_9_1/GATE sky130_asc_res_xhigh_po_2p85_1_12/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_25 sky130_asc_res_xhigh_po_2p85_1_25/Rin sky130_asc_res_xhigh_po_2p85_1_29/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_12_1 VDD VDD sky130_asc_cap_mim_m3_1_9/Cin VSS VDD sky130_asc_pfet_01v8_lvt_12
Xsky130_asc_res_xhigh_po_2p85_1_15 sky130_asc_res_xhigh_po_2p85_1_9/Rout sky130_asc_res_xhigh_po_2p85_1_16/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_26 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_res_xhigh_po_2p85_1_25/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_16 sky130_asc_res_xhigh_po_2p85_1_16/Rin sky130_asc_res_xhigh_po_2p85_1_17/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_27 sky130_asc_res_xhigh_po_2p85_1_27/Rin sky130_asc_res_xhigh_po_2p85_2_1/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_17 sky130_asc_res_xhigh_po_2p85_1_17/Rin sky130_asc_res_xhigh_po_2p85_1_18/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_28 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_10/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_nfet_01v8_lvt_9_0 porst VSS sky130_asc_cap_mim_m3_1_4/Cout VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_pfet_01v8_lvt_6_0 sky130_asc_pfet_01v8_lvt_6_1/GATE VDD sky130_asc_pfet_01v8_lvt_6_1/GATE
+ VSS VDD sky130_asc_pfet_01v8_lvt_6
Xsky130_asc_res_xhigh_po_2p85_1_18 sky130_asc_res_xhigh_po_2p85_1_18/Rin sky130_asc_res_xhigh_po_2p85_1_30/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_29 sky130_asc_res_xhigh_po_2p85_1_29/Rin sky130_asc_res_xhigh_po_2p85_1_27/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_nfet_01v8_lvt_9_1 sky130_asc_nfet_01v8_lvt_9_1/GATE sky130_asc_nfet_01v8_lvt_1_0/DRAIN
+ sky130_asc_pfet_01v8_lvt_6_1/GATE VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_pfet_01v8_lvt_6_1 sky130_asc_pfet_01v8_lvt_6_1/GATE VDD sky130_asc_cap_mim_m3_1_4/Cout
+ VSS VDD sky130_asc_pfet_01v8_lvt_6
Xsky130_asc_res_xhigh_po_2p85_1_19 sky130_asc_res_xhigh_po_2p85_1_19/Rin sky130_asc_res_xhigh_po_2p85_1_26/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pnp_05v5_W3p40L3p40_1_0 sky130_asc_cap_mim_m3_1_9/Cin VSS VSS VDD VSS
+ sky130_asc_pnp_05v5_W3p40L3p40_1
Xsky130_asc_nfet_01v8_lvt_9_2 sky130_asc_cap_mim_m3_1_9/Cin sky130_asc_nfet_01v8_lvt_1_0/DRAIN
+ sky130_asc_cap_mim_m3_1_4/Cout VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_cap_mim_m3_1_0 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_cap_mim_m3_1_1 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_0 sky130_asc_res_xhigh_po_2p85_1_12/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_2 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_1 sky130_asc_res_xhigh_po_2p85_1_12/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_3 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_2 sky130_asc_res_xhigh_po_2p85_1_12/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_4 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_3 sky130_asc_res_xhigh_po_2p85_1_12/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_5 sky130_asc_cap_mim_m3_1_9/Cin VSS VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_0 sky130_asc_res_xhigh_po_2p85_1_0/Rin sky130_asc_res_xhigh_po_2p85_1_8/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_6 sky130_asc_cap_mim_m3_1_9/Cin VSS VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_nfet_01v8_lvt_1_0 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS sky130_asc_nfet_01v8_lvt_1_0/DRAIN
+ VDD VSS sky130_asc_nfet_01v8_lvt_1
Xsky130_asc_res_xhigh_po_2p85_1_1 sky130_asc_res_xhigh_po_2p85_1_1/Rin sky130_asc_res_xhigh_po_2p85_1_5/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_7 sky130_asc_cap_mim_m3_1_9/Cin VSS VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_nfet_01v8_lvt_1_1 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS sky130_asc_nfet_01v8_lvt_1_1/GATE
+ VDD VSS sky130_asc_nfet_01v8_lvt_1
Xsky130_asc_res_xhigh_po_2p85_1_2 sky130_asc_res_xhigh_po_2p85_1_2/Rin sky130_asc_res_xhigh_po_2p85_1_4/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_8 sky130_asc_cap_mim_m3_1_9/Cin VSS VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_3 sky130_asc_res_xhigh_po_2p85_1_3/Rin VSS VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_9 sky130_asc_cap_mim_m3_1_9/Cin VSS VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_4 sky130_asc_res_xhigh_po_2p85_1_4/Rin sky130_asc_res_xhigh_po_2p85_1_0/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_5 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_6/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_6 sky130_asc_res_xhigh_po_2p85_1_6/Rin sky130_asc_res_xhigh_po_2p85_1_3/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
.ends

.subckt bgr_top porst vbg VDD VSS
Xsky130_asc_res_xhigh_po_2p85_1_7 sky130_asc_res_xhigh_po_2p85_1_7/Rin sky130_asc_res_xhigh_po_2p85_1_7/Rout
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_8 sky130_asc_res_xhigh_po_2p85_1_8/Rin sky130_asc_res_xhigh_po_2p85_1_7/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_9 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rout
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_60_0 sky130_asc_cap_mim_m3_1_9/Cout VDD sky130_asc_cap_mim_m3_1_4/Cin
+ VSS VDD sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_pfet_01v8_lvt_60_1 sky130_asc_cap_mim_m3_1_9/Cout VDD sky130_asc_nfet_01v8_lvt_9_1/GATE
+ VSS VDD sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_pfet_01v8_lvt_60_2 sky130_asc_cap_mim_m3_1_9/Cout VDD vbg VSS VDD sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_res_xhigh_po_2p85_1_30 sky130_asc_res_xhigh_po_2p85_1_9/Rout sky130_asc_res_xhigh_po_2p85_1_25/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_20 sky130_asc_res_xhigh_po_2p85_1_20/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pnp_05v5_W3p40L3p40_7_0 sky130_asc_res_xhigh_po_2p85_1_0/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_7
Xsky130_asc_res_xhigh_po_2p85_1_10 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_13/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_21 sky130_asc_res_xhigh_po_2p85_1_21/Rin sky130_asc_res_xhigh_po_2p85_1_20/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_2_0 sky130_asc_res_xhigh_po_2p85_2_0/Rin VSS VDD VSS
+ sky130_asc_res_xhigh_po_2p85_2
Xsky130_asc_res_xhigh_po_2p85_1_11 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_22 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_2_1 sky130_asc_res_xhigh_po_2p85_2_1/Rin VSS VDD VSS
+ sky130_asc_res_xhigh_po_2p85_2
Xsky130_asc_res_xhigh_po_2p85_1_12 sky130_asc_res_xhigh_po_2p85_1_7/Rout sky130_asc_res_xhigh_po_2p85_1_15/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_23 sky130_asc_res_xhigh_po_2p85_1_23/Rin sky130_asc_res_xhigh_po_2p85_2_1/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_13 sky130_asc_res_xhigh_po_2p85_1_13/Rin sky130_asc_res_xhigh_po_2p85_1_14/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_24 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_12_0 sky130_asc_cap_mim_m3_1_9/Cout VDD sky130_asc_nfet_01v8_lvt_1_1/GATE
+ VSS VDD sky130_asc_pfet_01v8_lvt_12
Xsky130_asc_res_xhigh_po_2p85_1_14 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_2_0/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_25 sky130_asc_res_xhigh_po_2p85_1_25/Rin sky130_asc_res_xhigh_po_2p85_1_4/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_12_1 VDD VDD sky130_asc_cap_mim_m3_1_4/Cin VSS VDD sky130_asc_pfet_01v8_lvt_12
Xsky130_asc_res_xhigh_po_2p85_1_15 sky130_asc_res_xhigh_po_2p85_1_15/Rin sky130_asc_res_xhigh_po_2p85_1_10/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_26 sky130_asc_res_xhigh_po_2p85_1_5/Rout VSS VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_16 sky130_asc_res_xhigh_po_2p85_1_16/Rin sky130_asc_res_xhigh_po_2p85_1_22/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_27 sky130_asc_res_xhigh_po_2p85_1_6/Rout sky130_asc_res_xhigh_po_2p85_1_28/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_17 sky130_asc_nfet_01v8_lvt_9_1/GATE sky130_asc_res_xhigh_po_2p85_1_0/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_28 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_18/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_nfet_01v8_lvt_9_0 sky130_asc_cap_mim_m3_1_4/Cin sky130_asc_nfet_01v8_lvt_1_1/DRAIN
+ sky130_asc_cap_mim_m3_1_9/Cout VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_pfet_01v8_lvt_6_0 sky130_asc_pfet_01v8_lvt_6_1/GATE VDD sky130_asc_cap_mim_m3_1_9/Cout
+ VSS VDD sky130_asc_pfet_01v8_lvt_6
Xsky130_asc_res_xhigh_po_2p85_1_18 sky130_asc_res_xhigh_po_2p85_1_18/Rin sky130_asc_res_xhigh_po_2p85_1_16/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_29 vbg sky130_asc_res_xhigh_po_2p85_1_11/Rin VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_nfet_01v8_lvt_9_1 sky130_asc_nfet_01v8_lvt_9_1/GATE sky130_asc_nfet_01v8_lvt_1_1/DRAIN
+ sky130_asc_pfet_01v8_lvt_6_1/GATE VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_res_xhigh_po_2p85_1_19 sky130_asc_res_xhigh_po_2p85_1_19/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_6_1 sky130_asc_pfet_01v8_lvt_6_1/GATE VDD sky130_asc_pfet_01v8_lvt_6_1/GATE
+ VSS VDD sky130_asc_pfet_01v8_lvt_6
Xsky130_asc_pnp_05v5_W3p40L3p40_1_0 sky130_asc_cap_mim_m3_1_4/Cin VSS VSS VDD VSS
+ sky130_asc_pnp_05v5_W3p40L3p40_1
Xsky130_asc_nfet_01v8_lvt_9_2 porst VSS sky130_asc_cap_mim_m3_1_9/Cout VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_cap_mim_m3_1_0 sky130_asc_cap_mim_m3_1_4/Cin VSS VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_cap_mim_m3_1_1 sky130_asc_cap_mim_m3_1_4/Cin VSS VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_0 sky130_asc_res_xhigh_po_2p85_1_0/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_2 sky130_asc_cap_mim_m3_1_4/Cin VSS VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_1 sky130_asc_res_xhigh_po_2p85_1_0/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_3 sky130_asc_cap_mim_m3_1_4/Cin VSS VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_2 sky130_asc_res_xhigh_po_2p85_1_0/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_4 sky130_asc_cap_mim_m3_1_4/Cin VSS VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_3 sky130_asc_res_xhigh_po_2p85_1_0/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_5 VDD sky130_asc_cap_mim_m3_1_9/Cout VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_0 sky130_asc_res_xhigh_po_2p85_1_0/Rin sky130_asc_res_xhigh_po_2p85_1_0/Rout
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_6 VDD sky130_asc_cap_mim_m3_1_9/Cout VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_nfet_01v8_lvt_1_0 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS sky130_asc_nfet_01v8_lvt_1_1/GATE
+ VDD VSS sky130_asc_nfet_01v8_lvt_1
Xsky130_asc_res_xhigh_po_2p85_1_1 sky130_asc_cap_mim_m3_1_4/Cin sky130_asc_res_xhigh_po_2p85_1_2/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_7 VDD sky130_asc_cap_mim_m3_1_9/Cout VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_nfet_01v8_lvt_1_1 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS sky130_asc_nfet_01v8_lvt_1_1/DRAIN
+ VDD VSS sky130_asc_nfet_01v8_lvt_1
Xsky130_asc_res_xhigh_po_2p85_1_2 sky130_asc_res_xhigh_po_2p85_1_2/Rin sky130_asc_res_xhigh_po_2p85_1_3/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_8 VDD sky130_asc_cap_mim_m3_1_9/Cout VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_3 sky130_asc_res_xhigh_po_2p85_1_3/Rin sky130_asc_res_xhigh_po_2p85_1_8/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_9 VDD sky130_asc_cap_mim_m3_1_9/Cout VDD VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_4 sky130_asc_res_xhigh_po_2p85_1_4/Rin sky130_asc_res_xhigh_po_2p85_1_5/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_5 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_5/Rout
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_6 sky130_asc_nfet_01v8_lvt_9_1/GATE sky130_asc_res_xhigh_po_2p85_1_6/Rout
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1
.ends

.subckt pmos_flat VGND SOURCE DRAIN GATE VPWR
X0 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X2 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X3 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X4 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X5 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X6 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X7 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X8 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X9 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X10 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X11 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X12 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X13 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X14 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X15 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X16 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X17 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X18 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X19 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[4] io_analog[5] io_analog[6] io_analog[7]
+ io_analog[8] io_analog[9] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xpuf_top_0 la_data_out[0] io_in[20] io_in[18] io_out[25] io_in[21] io_in[26] io_in[23]
+ io_in[17] io_in[22] vccd2 io_out[24] la_data_out[1] vssd2 io_in[19] puf_top
Xnmos_flat_0 vccd1 vssd2 gpio_analog[2] vssd2 vssd2 nmos_flat
Xsky130_fd_pr__res_generic_m4_LS59QM_0 vssd2 vssa1 sky130_fd_pr__res_generic_m4_LS59QM
Xnmos_flat_1 vccd1 vssd2 gpio_analog[1] vssd2 vssd2 nmos_flat
Xnmos_flat_3 vccd1 vssd2 gpio_analog[4] vssd2 vssd2 nmos_flat
Xnmos_flat_2 vccd1 vssd2 gpio_analog[3] vssd2 vssd2 nmos_flat
Xnmos_flat_4 vccd1 vssd2 gpio_analog[6] vssd2 vssd2 nmos_flat
Xnmos_flat_5 vccd1 vssd2 gpio_analog[5] vssd2 vssd2 nmos_flat
Xbandgaptop_flat_io_0 gpio_analog[6] vccd1 vssd2 gpio_analog[5] bandgaptop_flat_io
Xbgr_gen7_0 gpio_analog[2] gpio_analog[1] vssd2 vccd1 bgr_gen7
Xbgr_top_0 gpio_analog[4] gpio_analog[3] vccd1 vssd2 bgr_top
Xpmos_flat_0 vssd2 vccd1 gpio_analog[4] vccd1 vccd1 pmos_flat
Xpmos_flat_1 vssd2 vccd1 gpio_analog[3] vccd1 vccd1 pmos_flat
Xpmos_flat_2 vssd2 vccd1 gpio_analog[2] vccd1 vccd1 pmos_flat
Xpmos_flat_3 vssd2 vccd1 gpio_analog[1] vccd1 vccd1 pmos_flat
Xpmos_flat_4 vssd2 vccd1 gpio_analog[6] vccd1 vccd1 pmos_flat
Xpmos_flat_5 vssd2 vccd1 gpio_analog[5] vccd1 vccd1 pmos_flat
.ends

