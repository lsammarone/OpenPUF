//-----------------------------------------------------------------------------
// BR32 - Bistable Ring PUF 32-bit 
//-----------------------------------------------------------------------------
// dump-vcd: False
// verilator-xinit: zeros
module BR32 
(
  input wire RESET,
  input wire [31:0] C,
  output wire OUT
);
  supply1 VDD;
  supply0 VSS;
  // empty module
  // see lib file
  
endmodule
