magic
tech sky130A
magscale 1 2
timestamp 1483428465
<< checkpaint >>
rect -1569 -1402 1569 1402
<< metal4 >>
rect -309 118 309 142
rect -309 -118 -278 118
rect -42 -118 42 118
rect 278 -118 309 118
rect -309 -142 309 -118
<< via4 >>
rect -278 -118 -42 118
rect 42 -118 278 118
<< metal5 >>
rect -309 118 309 142
rect -309 -118 -278 118
rect -42 -118 42 118
rect 278 -118 309 118
rect -309 -142 309 -118
<< end >>
