magic
tech sky130A
magscale 1 2
timestamp 1655322987
<< metal4 >>
rect -1000 438 1000 571
rect -1000 -438 -918 438
rect 918 -438 1000 438
rect -1000 -571 1000 -438
<< via4 >>
rect -918 -438 918 438
<< metal5 >>
rect -1000 438 1000 571
rect -1000 -438 -918 438
rect 918 -438 1000 438
rect -1000 -571 1000 -438
<< end >>
