magic
tech sky130A
magscale 1 2
timestamp 1654736712
<< nwell >>
rect 10784 7195 10824 7516
rect 11708 7195 11748 7516
<< locali >>
rect 10990 7299 11034 7300
rect 10990 7265 10995 7299
rect 11029 7265 11034 7299
rect 10990 7264 11034 7265
rect 10072 7188 10124 7190
rect 10072 7154 10081 7188
rect 10115 7154 10124 7188
rect 10620 7189 10662 7190
rect 10620 7155 10624 7189
rect 10658 7155 10662 7189
rect 10620 7154 10662 7155
rect 10992 7187 11034 7188
rect 10072 7152 10124 7154
rect 10992 7153 10996 7187
rect 11030 7153 11034 7187
rect 11768 7160 11769 7194
rect 11803 7160 11804 7194
rect 10992 7152 11034 7153
<< viali >>
rect 10995 7265 11029 7299
rect 10081 7154 10115 7188
rect 10624 7155 10658 7189
rect 10996 7153 11030 7187
rect 11769 7160 11803 7194
<< metal1 >>
rect 10632 7430 10942 7526
rect 11576 7432 11866 7528
rect 10426 7299 11812 7306
rect 10426 7265 10995 7299
rect 11029 7265 11812 7299
rect 10426 7258 11812 7265
rect 10426 7198 10474 7258
rect 11764 7200 11812 7258
rect 10044 7188 10474 7198
rect 10044 7154 10081 7188
rect 10115 7154 10474 7188
rect 10044 7150 10474 7154
rect 10604 7189 11048 7196
rect 10604 7155 10624 7189
rect 10658 7187 11048 7189
rect 10658 7155 10996 7187
rect 10604 7153 10996 7155
rect 11030 7153 11048 7187
rect 11756 7194 11816 7200
rect 11756 7160 11769 7194
rect 11803 7160 11816 7194
rect 11756 7154 11816 7160
rect 10060 7146 10136 7150
rect 10604 7146 11048 7153
rect 10632 6886 10942 6982
rect 11542 6886 11832 6982
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0
timestamp 1654736712
transform 1 0 10496 0 1 6934
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0
timestamp 1654736712
transform 1 0 10852 0 1 6934
box -38 -48 866 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0
timestamp 1654736712
transform 1 0 11762 0 1 6934
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1654736712
transform 1 0 9030 0 1 6934
box -38 -48 1510 592
<< end >>
