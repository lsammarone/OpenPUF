magic
tech sky130A
timestamp 1654736712
<< metal4 >>
rect -155 459 155 500
rect -155 -459 -139 459
rect 139 -459 155 459
rect -155 -500 155 -459
<< via4 >>
rect -139 -459 139 459
<< metal5 >>
rect -155 459 155 500
rect -155 -459 -139 459
rect 139 -459 155 459
rect -155 -500 155 -459
<< end >>
