magic
tech sky130A
magscale 1 2
timestamp 1483428465
<< checkpaint >>
rect -1260 -3558 62809 11458
<< nwell >>
rect 31643 4383 32021 5502
rect 31376 4354 32021 4383
rect 31376 4062 31912 4354
rect 15656 3686 16038 4007
rect 45798 3846 46180 4167
<< nsubdiff >>
rect 45923 4019 46057 4038
rect 45923 3985 45995 4019
rect 46029 3985 46057 4019
rect 45923 3968 46057 3985
rect 15781 3859 15915 3878
rect 15781 3825 15853 3859
rect 15887 3825 15915 3859
rect 15781 3808 15915 3825
<< nsubdiffcont >>
rect 45995 3985 46029 4019
rect 15853 3825 15887 3859
<< locali >>
rect 30618 4060 30974 4066
rect 30618 4026 30665 4060
rect 30699 4026 30753 4060
rect 30787 4026 30974 4060
rect 30618 4016 30974 4026
rect 45720 4019 46263 4039
rect 45720 3985 45995 4019
rect 46029 3985 46263 4019
rect 45720 3967 46263 3985
rect 44589 3945 44623 3951
rect 44421 3938 44455 3944
rect 44925 3947 44959 3953
rect 44589 3906 44623 3911
rect 44757 3935 44791 3941
rect 44421 3899 44455 3904
rect 44925 3908 44959 3913
rect 45091 3945 45125 3951
rect 45091 3906 45125 3911
rect 45257 3947 45291 3953
rect 45257 3908 45291 3913
rect 45425 3947 45459 3953
rect 45425 3908 45459 3913
rect 45599 3945 45633 3951
rect 45599 3906 45633 3911
rect 46355 3939 46389 3945
rect 44757 3896 44791 3901
rect 46355 3900 46389 3905
rect 46517 3943 46551 3949
rect 46517 3904 46551 3909
rect 46687 3947 46721 3953
rect 46687 3908 46721 3913
rect 46851 3943 46885 3949
rect 46851 3904 46885 3909
rect 47021 3943 47055 3949
rect 47021 3904 47055 3909
rect 47189 3939 47223 3945
rect 47189 3900 47223 3905
rect 47357 3943 47391 3949
rect 47357 3904 47391 3909
rect 47531 3939 47565 3945
rect 47531 3900 47565 3905
rect 15578 3859 16121 3879
rect 15578 3825 15853 3859
rect 15887 3825 16121 3859
rect 15578 3807 16121 3825
rect 14447 3785 14481 3791
rect 14279 3778 14313 3784
rect 14783 3787 14817 3793
rect 14447 3746 14481 3751
rect 14615 3775 14649 3781
rect 14279 3739 14313 3744
rect 14783 3748 14817 3753
rect 14949 3785 14983 3791
rect 14949 3746 14983 3751
rect 15115 3787 15149 3793
rect 15115 3748 15149 3753
rect 15283 3787 15317 3793
rect 15283 3748 15317 3753
rect 15457 3785 15491 3791
rect 15457 3746 15491 3751
rect 16213 3779 16247 3785
rect 14615 3736 14649 3741
rect 16213 3740 16247 3745
rect 16375 3783 16409 3789
rect 16375 3744 16409 3749
rect 16545 3787 16579 3793
rect 16545 3748 16579 3753
rect 16709 3783 16743 3789
rect 16709 3744 16743 3749
rect 16879 3783 16913 3789
rect 16879 3744 16913 3749
rect 17047 3779 17081 3785
rect 17047 3740 17081 3745
rect 17215 3783 17249 3789
rect 17215 3744 17249 3749
rect 17389 3779 17423 3785
rect 17389 3740 17423 3745
<< viali >>
rect 30665 4026 30699 4060
rect 30753 4026 30787 4060
rect 31330 4058 31364 4092
rect 31601 4022 31635 4056
rect 31689 4022 31723 4056
rect 31777 4022 31811 4056
rect 31865 4022 31899 4056
rect 31953 4022 31987 4056
rect 32041 4022 32075 4056
rect 32129 4022 32163 4056
rect 32217 4022 32251 4056
rect 31330 3978 31364 4012
rect 31955 3920 31989 3954
rect 32121 3916 32155 3950
rect 32289 3922 32323 3956
rect 32456 3920 32490 3954
rect 32626 3921 32660 3955
rect 32790 3922 32824 3956
rect 44421 3904 44455 3938
rect 44589 3911 44623 3945
rect 44757 3901 44791 3935
rect 44925 3913 44959 3947
rect 45091 3911 45125 3945
rect 45257 3913 45291 3947
rect 45425 3913 45459 3947
rect 45599 3911 45633 3945
rect 46355 3905 46389 3939
rect 46517 3909 46551 3943
rect 46687 3913 46721 3947
rect 46851 3909 46885 3943
rect 47021 3909 47055 3943
rect 47189 3905 47223 3939
rect 47357 3909 47391 3943
rect 47531 3905 47565 3939
rect 44621 3808 44655 3842
rect 44721 3808 44755 3842
rect 44821 3808 44855 3842
rect 44921 3808 44955 3842
rect 45021 3808 45055 3842
rect 45121 3808 45155 3842
rect 45221 3808 45255 3842
rect 45321 3808 45355 3842
rect 46281 3808 46315 3842
rect 46381 3808 46415 3842
rect 46481 3808 46515 3842
rect 46581 3808 46615 3842
rect 46681 3808 46715 3842
rect 46781 3808 46815 3842
rect 46881 3808 46915 3842
rect 46981 3808 47015 3842
rect 14279 3744 14313 3778
rect 14447 3751 14481 3785
rect 14615 3741 14649 3775
rect 14783 3753 14817 3787
rect 14949 3751 14983 3785
rect 15115 3753 15149 3787
rect 15283 3753 15317 3787
rect 15457 3751 15491 3785
rect 16213 3745 16247 3779
rect 16375 3749 16409 3783
rect 16545 3753 16579 3787
rect 16709 3749 16743 3783
rect 16879 3749 16913 3783
rect 17047 3745 17081 3779
rect 17215 3749 17249 3783
rect 17389 3745 17423 3779
rect 14479 3648 14513 3682
rect 14579 3648 14613 3682
rect 14679 3648 14713 3682
rect 14779 3648 14813 3682
rect 14879 3648 14913 3682
rect 14979 3648 15013 3682
rect 15079 3648 15113 3682
rect 15179 3648 15213 3682
rect 16139 3648 16173 3682
rect 16239 3648 16273 3682
rect 16339 3648 16373 3682
rect 16439 3648 16473 3682
rect 16539 3648 16573 3682
rect 16639 3648 16673 3682
rect 16739 3648 16773 3682
rect 16839 3648 16873 3682
<< metal1 >>
rect 15330 4977 15585 5333
rect 31266 5000 31600 5324
rect 15330 4925 15350 4977
rect 15402 4925 15428 4977
rect 15480 4925 15521 4977
rect 15573 4925 15585 4977
rect 15330 4895 15585 4925
rect 31266 4948 31309 5000
rect 31361 4948 31422 5000
rect 31474 4948 31523 5000
rect 31575 4948 31600 5000
rect 31266 4904 31600 4948
rect 45470 4977 45697 5345
rect 45470 4925 45501 4977
rect 45553 4925 45584 4977
rect 45636 4925 45697 4977
rect 45470 4891 45697 4925
rect 7986 4760 8522 4844
rect 23020 4769 23628 4827
rect 38124 4777 38748 4835
rect 53130 4783 53863 4841
rect 31394 4380 31502 4393
rect 31394 4328 31424 4380
rect 31476 4328 31502 4380
rect 31394 4297 31502 4328
rect 32934 4297 32969 4393
rect 0 4161 18000 4227
rect 17934 4075 18000 4161
rect 45639 4153 46306 4162
rect 31315 4092 31394 4120
rect 45649 4104 46306 4153
rect 17934 4060 30881 4075
rect 17934 4026 30665 4060
rect 30699 4026 30753 4060
rect 30787 4026 30881 4060
rect 17934 4009 30881 4026
rect 31315 4058 31330 4092
rect 31364 4064 31394 4092
rect 31364 4058 32313 4064
rect 31315 4056 32313 4058
rect 31315 4022 31601 4056
rect 31635 4022 31689 4056
rect 31723 4022 31777 4056
rect 31811 4022 31865 4056
rect 31899 4022 31953 4056
rect 31987 4022 32041 4056
rect 32075 4022 32129 4056
rect 32163 4022 32217 4056
rect 32251 4022 32313 4056
rect 31315 4016 32313 4022
rect 31315 4012 31397 4016
rect 15549 3948 16198 3998
rect 31315 3978 31330 4012
rect 31364 3978 31397 4012
rect 31315 3960 31397 3978
rect 31886 3971 32831 3984
rect 15497 3940 16198 3948
rect 31886 3954 32102 3971
rect 31886 3920 31955 3954
rect 31989 3920 32102 3954
rect 32154 3950 32262 3971
rect 32314 3956 32395 3971
rect 31886 3919 32102 3920
rect 32155 3919 32262 3950
rect 32323 3922 32395 3956
rect 32314 3919 32395 3922
rect 32447 3954 32508 3971
rect 32447 3920 32456 3954
rect 32490 3920 32508 3954
rect 32447 3919 32508 3920
rect 32560 3956 32831 3971
rect 32560 3955 32790 3956
rect 32560 3921 32626 3955
rect 32660 3922 32790 3955
rect 32824 3922 32831 3956
rect 32660 3921 32831 3922
rect 32560 3919 32831 3921
rect 31886 3916 32121 3919
rect 32155 3916 32831 3919
rect 31886 3901 32831 3916
rect 38288 3947 53723 3963
rect 38288 3945 44925 3947
rect 38288 3944 44589 3945
rect 38288 3943 38470 3944
rect 38288 3891 38367 3943
rect 38419 3892 38470 3943
rect 38522 3938 44589 3944
rect 38522 3904 44421 3938
rect 44455 3911 44589 3938
rect 44623 3935 44925 3945
rect 44623 3911 44757 3935
rect 44455 3904 44757 3911
rect 38522 3901 44757 3904
rect 44791 3913 44925 3935
rect 44959 3945 45257 3947
rect 44959 3913 45091 3945
rect 44791 3911 45091 3913
rect 45125 3913 45257 3945
rect 45291 3913 45425 3947
rect 45459 3945 46687 3947
rect 45459 3913 45599 3945
rect 45125 3911 45599 3913
rect 45633 3943 46687 3945
rect 45633 3939 46517 3943
rect 45633 3911 46355 3939
rect 44791 3905 46355 3911
rect 46389 3909 46517 3939
rect 46551 3913 46687 3943
rect 46721 3944 53723 3947
rect 46721 3943 53571 3944
rect 46721 3913 46851 3943
rect 46551 3909 46851 3913
rect 46885 3909 47021 3943
rect 47055 3939 47357 3943
rect 47055 3909 47189 3939
rect 46389 3905 47189 3909
rect 47223 3909 47357 3939
rect 47391 3939 53571 3943
rect 47391 3909 47531 3939
rect 47223 3905 47531 3909
rect 47565 3905 53480 3939
rect 44791 3901 53480 3905
rect 38522 3892 53480 3901
rect 38419 3891 53480 3892
rect 38288 3887 53480 3891
rect 53532 3892 53571 3939
rect 53623 3892 53723 3944
rect 53532 3887 53723 3892
rect 38288 3882 53723 3887
rect 31394 3830 31497 3849
rect 31394 3827 31484 3830
rect 8131 3788 23497 3803
rect 8131 3736 8172 3788
rect 8224 3736 8268 3788
rect 8320 3787 23497 3788
rect 8320 3785 14783 3787
rect 8320 3778 14447 3785
rect 8320 3744 14279 3778
rect 14313 3751 14447 3778
rect 14481 3775 14783 3785
rect 14481 3751 14615 3775
rect 14313 3744 14615 3751
rect 8320 3741 14615 3744
rect 14649 3753 14783 3775
rect 14817 3785 15115 3787
rect 14817 3753 14949 3785
rect 14649 3751 14949 3753
rect 14983 3753 15115 3785
rect 15149 3753 15283 3787
rect 15317 3785 16545 3787
rect 15317 3753 15457 3785
rect 14983 3751 15457 3753
rect 15491 3783 16545 3785
rect 15491 3779 16375 3783
rect 15491 3751 16213 3779
rect 14649 3745 16213 3751
rect 16247 3749 16375 3779
rect 16409 3753 16545 3783
rect 16579 3786 23497 3787
rect 16579 3783 23382 3786
rect 16579 3753 16709 3783
rect 16409 3749 16709 3753
rect 16743 3749 16879 3783
rect 16913 3779 17215 3783
rect 16913 3749 17047 3779
rect 16247 3745 17047 3749
rect 17081 3749 17215 3779
rect 17249 3779 23382 3783
rect 17249 3749 17389 3779
rect 17081 3745 17389 3749
rect 17423 3745 23283 3779
rect 14649 3741 23283 3745
rect 8320 3736 23283 3741
rect 8131 3727 23283 3736
rect 23335 3734 23382 3779
rect 23434 3734 23497 3786
rect 31425 3778 31484 3827
rect 31425 3775 31497 3778
rect 31394 3753 31497 3775
rect 32934 3753 32969 3849
rect 44589 3842 47192 3848
rect 44589 3808 44621 3842
rect 44655 3808 44721 3842
rect 44755 3808 44821 3842
rect 44855 3808 44921 3842
rect 44955 3808 45021 3842
rect 45055 3808 45121 3842
rect 45155 3808 45221 3842
rect 45255 3808 45321 3842
rect 45355 3808 46281 3842
rect 46315 3808 46381 3842
rect 46415 3808 46481 3842
rect 46515 3808 46581 3842
rect 46615 3808 46681 3842
rect 46715 3808 46781 3842
rect 46815 3808 46881 3842
rect 46915 3808 46981 3842
rect 47015 3808 47192 3842
rect 44589 3803 47192 3808
rect 44589 3800 46035 3803
rect 45885 3799 46035 3800
rect 23335 3727 23497 3734
rect 8131 3722 23497 3727
rect 45885 3747 45930 3799
rect 45982 3751 46035 3799
rect 46087 3800 47192 3803
rect 46087 3751 46113 3800
rect 45982 3747 46113 3751
rect 45885 3708 46113 3747
rect 14447 3682 17050 3688
rect 14447 3648 14479 3682
rect 14513 3648 14579 3682
rect 14613 3648 14679 3682
rect 14713 3648 14779 3682
rect 14813 3648 14879 3682
rect 14913 3648 14979 3682
rect 15013 3648 15079 3682
rect 15113 3648 15179 3682
rect 15213 3648 16139 3682
rect 16173 3648 16239 3682
rect 16273 3648 16339 3682
rect 16373 3648 16439 3682
rect 16473 3648 16539 3682
rect 16573 3648 16639 3682
rect 16673 3648 16739 3682
rect 16773 3648 16839 3682
rect 16873 3648 17050 3682
rect 14447 3643 17050 3648
rect 14447 3640 15893 3643
rect 15743 3639 15893 3640
rect 15743 3587 15788 3639
rect 15840 3591 15893 3639
rect 15945 3640 17050 3643
rect 15945 3591 15971 3640
rect 15840 3587 15971 3591
rect 15743 3548 15971 3587
rect 45639 3556 46391 3614
rect 14109 3378 14160 3474
rect 15497 3402 16178 3460
rect 20628 3405 46139 3449
rect 20628 3403 46027 3405
rect 14109 3377 14159 3378
rect 20628 3351 32091 3403
rect 32143 3351 32235 3403
rect 32287 3351 32379 3403
rect 32431 3402 46027 3403
rect 32431 3351 45938 3402
rect 20628 3350 45938 3351
rect 45990 3353 46027 3402
rect 46079 3353 46139 3405
rect 45990 3350 46139 3353
rect 20628 3326 46139 3350
rect 20628 3319 45938 3326
rect 20628 3267 32090 3319
rect 32142 3267 32234 3319
rect 32286 3267 32378 3319
rect 32430 3274 45938 3319
rect 45990 3274 46031 3326
rect 46083 3274 46139 3326
rect 32430 3267 46139 3274
rect 15755 3243 46139 3267
rect 15755 3222 20834 3243
rect 15755 3170 15792 3222
rect 15844 3217 20834 3222
rect 15844 3170 15886 3217
rect 15755 3165 15886 3170
rect 15938 3165 20834 3217
rect 15755 3144 20834 3165
rect 15755 3142 15886 3144
rect 7922 3068 8585 3126
rect 15755 3090 15792 3142
rect 15844 3092 15886 3142
rect 15938 3092 20834 3144
rect 15844 3090 20834 3092
rect 15755 3061 20834 3090
rect 23020 3080 23648 3138
rect 38032 3080 38795 3138
rect 53222 3071 53873 3129
rect 61289 1010 61511 1088
<< via1 >>
rect 8171 4991 8223 5043
rect 8252 4990 8304 5042
rect 23287 4988 23339 5040
rect 23382 4988 23434 5040
rect 15350 4925 15402 4977
rect 15428 4925 15480 4977
rect 15521 4925 15573 4977
rect 31309 4948 31361 5000
rect 31422 4948 31474 5000
rect 31523 4948 31575 5000
rect 38364 4990 38416 5042
rect 38466 4990 38518 5042
rect 45501 4925 45553 4977
rect 45584 4925 45636 4977
rect 53482 4963 53534 5015
rect 53577 4963 53629 5015
rect 7179 4769 7231 4821
rect 7286 4771 7338 4823
rect 7388 4771 7440 4823
rect 7488 4772 7540 4824
rect 22209 4775 22261 4827
rect 22312 4775 22364 4827
rect 22395 4775 22447 4827
rect 22496 4775 22548 4827
rect 22583 4775 22635 4827
rect 37341 4771 37393 4823
rect 37429 4771 37481 4823
rect 37514 4776 37566 4828
rect 54257 4768 54309 4820
rect 54351 4768 54403 4820
rect 54428 4768 54480 4820
rect 54508 4767 54560 4819
rect 54582 4768 54634 4820
rect 31321 4325 31373 4377
rect 31424 4328 31476 4380
rect 31525 4328 31577 4380
rect 45507 4100 45559 4152
rect 45597 4101 45649 4153
rect 15374 3948 15426 4000
rect 15497 3948 15549 4000
rect 32102 3950 32154 3971
rect 32262 3956 32314 3971
rect 32102 3919 32121 3950
rect 32121 3919 32154 3950
rect 32262 3922 32289 3956
rect 32289 3922 32314 3956
rect 32262 3919 32314 3922
rect 32395 3919 32447 3971
rect 32508 3919 32560 3971
rect 38367 3891 38419 3943
rect 38470 3892 38522 3944
rect 53480 3887 53532 3939
rect 53571 3892 53623 3944
rect 8172 3736 8224 3788
rect 8268 3736 8320 3788
rect 23283 3727 23335 3779
rect 23382 3734 23434 3786
rect 31277 3773 31329 3825
rect 31373 3775 31425 3827
rect 31484 3778 31536 3830
rect 31576 3775 31628 3827
rect 45930 3747 45982 3799
rect 46035 3751 46087 3803
rect 15788 3587 15840 3639
rect 15893 3591 15945 3643
rect 46942 3560 46994 3612
rect 47034 3561 47086 3613
rect 47124 3560 47176 3612
rect 47212 3559 47264 3611
rect 14587 3399 14639 3451
rect 14671 3399 14723 3451
rect 14764 3400 14816 3452
rect 32091 3351 32143 3403
rect 32235 3351 32287 3403
rect 32379 3351 32431 3403
rect 45938 3350 45990 3402
rect 46027 3353 46079 3405
rect 32090 3267 32142 3319
rect 32234 3267 32286 3319
rect 32378 3267 32430 3319
rect 45938 3274 45990 3326
rect 46031 3274 46083 3326
rect 15792 3170 15844 3222
rect 15886 3165 15938 3217
rect 7173 3071 7225 3123
rect 7271 3071 7323 3123
rect 7366 3071 7418 3123
rect 7471 3071 7523 3123
rect 15792 3090 15844 3142
rect 15886 3092 15938 3144
rect 22223 3076 22275 3128
rect 22323 3076 22375 3128
rect 22422 3076 22474 3128
rect 22525 3076 22577 3128
rect 37331 3070 37383 3122
rect 37419 3070 37471 3122
rect 37517 3066 37569 3118
rect 54253 3067 54305 3119
rect 54341 3067 54393 3119
rect 54424 3067 54476 3119
rect 54511 3067 54563 3119
rect 8172 2853 8224 2905
rect 8252 2851 8304 2903
rect 23288 2868 23340 2920
rect 23371 2868 23423 2920
rect 38366 2858 38418 2910
rect 38457 2858 38509 2910
rect 53483 2843 53535 2895
rect 53566 2843 53618 2895
<< metal2 >>
rect 2297 6878 2341 8034
rect 4185 6878 4229 8034
rect 6073 6878 6117 8034
rect 7961 6878 8005 8034
rect 9849 6878 9893 8034
rect 11737 6878 11781 8034
rect 13625 6878 13669 8034
rect 15513 6878 15557 8034
rect 17401 6878 17445 8034
rect 19289 6878 19333 8034
rect 21177 6878 21221 8034
rect 23065 6878 23109 8034
rect 24953 6878 24997 8034
rect 26841 6878 26885 8034
rect 28729 6878 28773 8034
rect 30617 6878 30661 8034
rect 32505 6878 32549 8034
rect 34393 6878 34437 8034
rect 36281 6878 36325 8034
rect 38169 6878 38213 8034
rect 40057 6878 40101 8034
rect 41945 6878 41989 8034
rect 43833 6878 43877 8034
rect 45721 6878 45765 8034
rect 47609 6878 47653 8034
rect 49497 6878 49541 8034
rect 51385 6878 51429 8034
rect 53273 6878 53317 8034
rect 55161 6878 55205 8034
rect 57049 6878 57093 8034
rect 58937 6878 58981 8034
rect 60825 6878 60869 8034
rect 61398 6196 61512 6243
rect 271 6160 513 6196
rect 60845 6160 61512 6196
rect 271 6106 387 6160
rect 278 1740 368 6106
rect 8147 5043 8336 5073
rect 8147 4991 8171 5043
rect 8223 5042 8336 5043
rect 8223 4991 8252 5042
rect 8147 4990 8252 4991
rect 8304 4990 8336 5042
rect 7115 4824 7599 4949
rect 7115 4823 7488 4824
rect 7115 4821 7286 4823
rect 7115 4769 7179 4821
rect 7231 4771 7286 4821
rect 7338 4771 7388 4823
rect 7440 4772 7488 4823
rect 7540 4772 7599 4824
rect 7440 4771 7599 4772
rect 7231 4769 7599 4771
rect 7115 3602 7599 4769
rect 7115 3546 7182 3602
rect 7238 3546 7296 3602
rect 7352 3546 7410 3602
rect 7466 3546 7599 3602
rect 7115 3487 7599 3546
rect 7115 3431 7182 3487
rect 7238 3431 7296 3487
rect 7352 3431 7410 3487
rect 7466 3431 7599 3487
rect 7115 3372 7599 3431
rect 7115 3316 7182 3372
rect 7238 3316 7296 3372
rect 7352 3316 7410 3372
rect 7466 3316 7599 3372
rect 7115 3123 7599 3316
rect 7115 3071 7173 3123
rect 7225 3071 7271 3123
rect 7323 3071 7366 3123
rect 7418 3071 7471 3123
rect 7523 3071 7599 3123
rect 7115 2959 7599 3071
rect 8147 3788 8336 4990
rect 15330 4977 15590 5048
rect 15330 4925 15350 4977
rect 15402 4925 15428 4977
rect 15480 4925 15521 4977
rect 15573 4925 15590 4977
rect 23258 5040 23447 5063
rect 23258 4988 23287 5040
rect 23339 4988 23382 5040
rect 23434 4988 23447 5040
rect 15330 4000 15590 4925
rect 15330 3948 15374 4000
rect 15426 3948 15497 4000
rect 15549 3948 15590 4000
rect 15330 3904 15590 3948
rect 22171 4827 22638 4927
rect 22171 4775 22209 4827
rect 22261 4775 22312 4827
rect 22364 4775 22395 4827
rect 22447 4775 22496 4827
rect 22548 4775 22583 4827
rect 22635 4775 22638 4827
rect 8147 3736 8172 3788
rect 8224 3736 8268 3788
rect 8320 3736 8336 3788
rect 8147 2905 8336 3736
rect 15755 3643 15961 3688
rect 15755 3639 15893 3643
rect 15755 3587 15788 3639
rect 15840 3591 15893 3639
rect 15945 3591 15961 3643
rect 15840 3587 15961 3591
rect 8147 2853 8172 2905
rect 8224 2903 8336 2905
rect 8224 2853 8252 2903
rect 8147 2851 8252 2853
rect 8304 2851 8336 2903
rect 14536 3452 14889 3498
rect 14536 3451 14764 3452
rect 14536 3399 14587 3451
rect 14639 3399 14671 3451
rect 14723 3400 14764 3451
rect 14816 3400 14889 3452
rect 14723 3399 14889 3400
rect 14536 3041 14889 3399
rect 15755 3222 15961 3587
rect 15755 3170 15792 3222
rect 15844 3217 15961 3222
rect 15844 3170 15886 3217
rect 15755 3165 15886 3170
rect 15938 3165 15961 3217
rect 15755 3144 15961 3165
rect 15755 3142 15886 3144
rect 15755 3090 15792 3142
rect 15844 3092 15886 3142
rect 15938 3092 15961 3144
rect 15844 3090 15961 3092
rect 15755 3061 15961 3090
rect 22171 3512 22638 4775
rect 22171 3456 22221 3512
rect 22277 3456 22325 3512
rect 22381 3456 22429 3512
rect 22485 3456 22533 3512
rect 22589 3456 22638 3512
rect 22171 3396 22638 3456
rect 22171 3340 22221 3396
rect 22277 3340 22325 3396
rect 22381 3340 22429 3396
rect 22485 3340 22533 3396
rect 22589 3340 22638 3396
rect 22171 3280 22638 3340
rect 22171 3224 22221 3280
rect 22277 3224 22325 3280
rect 22381 3224 22429 3280
rect 22485 3224 22533 3280
rect 22589 3224 22638 3280
rect 22171 3128 22638 3224
rect 22171 3076 22223 3128
rect 22275 3076 22323 3128
rect 22375 3076 22422 3128
rect 22474 3076 22525 3128
rect 22577 3076 22638 3128
rect 14536 2985 14576 3041
rect 14632 2985 14684 3041
rect 14740 2985 14792 3041
rect 14848 2985 14889 3041
rect 14536 2947 14889 2985
rect 22171 2976 22638 3076
rect 23258 3786 23447 4988
rect 31263 5000 31598 5043
rect 31263 4948 31309 5000
rect 31361 4948 31422 5000
rect 31474 4948 31523 5000
rect 31575 4948 31598 5000
rect 31263 4380 31598 4948
rect 38349 5042 38536 5061
rect 38349 4990 38364 5042
rect 38416 4990 38466 5042
rect 38518 4990 38536 5042
rect 31263 4377 31424 4380
rect 31263 4325 31321 4377
rect 31373 4328 31424 4377
rect 31476 4328 31525 4380
rect 31577 4328 31598 4380
rect 31373 4325 31598 4328
rect 31263 4293 31598 4325
rect 37287 4828 37587 4925
rect 37287 4823 37514 4828
rect 37287 4771 37341 4823
rect 37393 4771 37429 4823
rect 37481 4776 37514 4823
rect 37566 4776 37587 4828
rect 37481 4771 37587 4776
rect 32034 3971 32573 3994
rect 32034 3919 32102 3971
rect 32154 3919 32262 3971
rect 32314 3919 32395 3971
rect 32447 3919 32508 3971
rect 32560 3919 32573 3971
rect 23258 3779 23382 3786
rect 23258 3727 23283 3779
rect 23335 3734 23382 3779
rect 23434 3734 23447 3786
rect 23335 3727 23447 3734
rect 14536 2891 14576 2947
rect 14632 2891 14684 2947
rect 14740 2891 14792 2947
rect 14848 2891 14889 2947
rect 14536 2865 14889 2891
rect 23258 2920 23447 3727
rect 31225 3830 31650 3848
rect 31225 3827 31484 3830
rect 31225 3825 31373 3827
rect 31225 3773 31277 3825
rect 31329 3775 31373 3825
rect 31425 3778 31484 3827
rect 31536 3827 31650 3830
rect 31536 3778 31576 3827
rect 31425 3775 31576 3778
rect 31628 3775 31650 3827
rect 31329 3773 31650 3775
rect 31225 3161 31650 3773
rect 32034 3403 32573 3919
rect 32034 3351 32091 3403
rect 32143 3351 32235 3403
rect 32287 3351 32379 3403
rect 32431 3351 32573 3403
rect 32034 3319 32573 3351
rect 32034 3267 32090 3319
rect 32142 3267 32234 3319
rect 32286 3267 32378 3319
rect 32430 3267 32573 3319
rect 32034 3193 32573 3267
rect 37287 3861 37587 4771
rect 37287 3805 37308 3861
rect 37364 3805 37402 3861
rect 37458 3805 37496 3861
rect 37552 3805 37587 3861
rect 37287 3773 37587 3805
rect 37287 3717 37308 3773
rect 37364 3717 37402 3773
rect 37458 3717 37496 3773
rect 37552 3717 37587 3773
rect 37287 3685 37587 3717
rect 37287 3629 37308 3685
rect 37364 3629 37402 3685
rect 37458 3629 37496 3685
rect 37552 3629 37587 3685
rect 31225 3105 31271 3161
rect 31327 3105 31396 3161
rect 31452 3105 31521 3161
rect 31577 3105 31650 3161
rect 31225 3065 31650 3105
rect 31225 3009 31271 3065
rect 31327 3009 31396 3065
rect 31452 3009 31521 3065
rect 31577 3009 31650 3065
rect 31225 2977 31650 3009
rect 37287 3122 37587 3629
rect 37287 3070 37331 3122
rect 37383 3070 37419 3122
rect 37471 3118 37587 3122
rect 37471 3070 37517 3118
rect 37287 3066 37517 3070
rect 37569 3066 37587 3118
rect 37287 2973 37587 3066
rect 38349 3944 38536 4990
rect 45478 4977 45697 5030
rect 45478 4925 45501 4977
rect 45553 4925 45584 4977
rect 45636 4925 45697 4977
rect 45478 4153 45697 4925
rect 45478 4152 45597 4153
rect 45478 4100 45507 4152
rect 45559 4101 45597 4152
rect 45649 4101 45697 4153
rect 45559 4100 45697 4101
rect 45478 4065 45697 4100
rect 53453 5015 53642 5038
rect 53453 4963 53482 5015
rect 53534 4963 53577 5015
rect 53629 4963 53642 5015
rect 38349 3943 38470 3944
rect 38349 3891 38367 3943
rect 38419 3892 38470 3943
rect 38522 3892 38536 3944
rect 38419 3891 38536 3892
rect 23258 2868 23288 2920
rect 23340 2868 23371 2920
rect 23423 2868 23447 2920
rect 23258 2855 23447 2868
rect 38349 2910 38536 3891
rect 53453 3944 53642 4963
rect 53453 3939 53571 3944
rect 53453 3887 53480 3939
rect 53532 3892 53571 3939
rect 53623 3892 53642 3944
rect 53532 3887 53642 3892
rect 45897 3803 46103 3848
rect 45897 3799 46035 3803
rect 45897 3747 45930 3799
rect 45982 3751 46035 3799
rect 46087 3751 46103 3803
rect 45982 3747 46103 3751
rect 45897 3405 46103 3747
rect 45897 3402 46027 3405
rect 45897 3350 45938 3402
rect 45990 3353 46027 3402
rect 46079 3353 46103 3405
rect 45990 3350 46103 3353
rect 45897 3326 46103 3350
rect 45897 3274 45938 3326
rect 45990 3274 46031 3326
rect 46083 3274 46103 3326
rect 45897 3231 46103 3274
rect 46905 3613 47319 3635
rect 46905 3612 47034 3613
rect 46905 3560 46942 3612
rect 46994 3561 47034 3612
rect 47086 3612 47319 3613
rect 47086 3561 47124 3612
rect 46994 3560 47124 3561
rect 47176 3611 47319 3612
rect 47176 3560 47212 3611
rect 46905 3559 47212 3560
rect 47264 3559 47319 3611
rect 38349 2858 38366 2910
rect 38418 2858 38457 2910
rect 38509 2858 38536 2910
rect 8147 2833 8336 2851
rect 38349 2850 38536 2858
rect 46905 3014 47319 3559
rect 46905 2958 46942 3014
rect 46998 2958 47035 3014
rect 47091 2958 47128 3014
rect 47184 2958 47221 3014
rect 47277 2958 47319 3014
rect 46905 2932 47319 2958
rect 46905 2876 46942 2932
rect 46998 2876 47035 2932
rect 47091 2876 47128 2932
rect 47184 2876 47221 2932
rect 47277 2876 47319 2932
rect 46905 2839 47319 2876
rect 53453 2895 53642 3887
rect 54218 4820 54639 4925
rect 54218 4768 54257 4820
rect 54309 4768 54351 4820
rect 54403 4768 54428 4820
rect 54480 4819 54582 4820
rect 54480 4768 54508 4819
rect 54218 4767 54508 4768
rect 54560 4768 54582 4819
rect 54634 4768 54639 4820
rect 54560 4767 54639 4768
rect 54218 3406 54639 4767
rect 54218 3350 54255 3406
rect 54311 3350 54359 3406
rect 54415 3350 54463 3406
rect 54519 3350 54567 3406
rect 54623 3350 54639 3406
rect 54218 3316 54639 3350
rect 54218 3260 54255 3316
rect 54311 3260 54359 3316
rect 54415 3260 54463 3316
rect 54519 3260 54567 3316
rect 54623 3260 54639 3316
rect 54218 3119 54639 3260
rect 54218 3067 54253 3119
rect 54305 3067 54341 3119
rect 54393 3067 54424 3119
rect 54476 3067 54511 3119
rect 54563 3067 54639 3119
rect 54218 2975 54639 3067
rect 53453 2843 53483 2895
rect 53535 2843 53566 2895
rect 53618 2843 53642 2895
rect 53453 2830 53642 2843
rect 61398 1818 61512 6160
rect 61355 1740 61549 1818
rect 273 1704 958 1740
rect 61283 1704 61549 1740
rect 278 1621 368 1704
rect 927 124 971 1022
rect 2815 124 2859 1022
rect 4703 124 4747 1022
rect 6591 124 6635 1022
rect 8479 124 8523 1022
rect 10367 124 10411 1022
rect 12255 124 12299 1022
rect 14143 124 14187 1022
rect 16031 124 16075 1022
rect 17919 124 17963 1022
rect 19807 124 19851 1022
rect 21695 124 21739 1022
rect 23583 124 23627 1022
rect 25471 124 25515 1022
rect 27359 24 27403 1022
rect 29247 124 29291 1022
rect 31135 124 31179 1022
rect 33023 124 33067 1022
rect 34911 124 34955 1022
rect 36799 124 36843 1022
rect 38687 124 38731 1022
rect 40575 0 40619 1022
rect 42463 124 42507 1022
rect 44351 124 44395 1022
rect 46239 124 46283 1022
rect 48127 124 48171 1022
rect 50015 124 50059 1022
rect 51903 124 51947 1022
rect 53791 124 53835 1022
rect 55679 124 55723 1022
rect 57567 902 57611 1022
rect 57567 124 57613 902
rect 59455 124 59499 1022
rect 57569 4 57613 124
<< via2 >>
rect 7182 3546 7238 3602
rect 7296 3546 7352 3602
rect 7410 3546 7466 3602
rect 7182 3431 7238 3487
rect 7296 3431 7352 3487
rect 7410 3431 7466 3487
rect 7182 3316 7238 3372
rect 7296 3316 7352 3372
rect 7410 3316 7466 3372
rect 22221 3456 22277 3512
rect 22325 3456 22381 3512
rect 22429 3456 22485 3512
rect 22533 3456 22589 3512
rect 22221 3340 22277 3396
rect 22325 3340 22381 3396
rect 22429 3340 22485 3396
rect 22533 3340 22589 3396
rect 22221 3224 22277 3280
rect 22325 3224 22381 3280
rect 22429 3224 22485 3280
rect 22533 3224 22589 3280
rect 14576 2985 14632 3041
rect 14684 2985 14740 3041
rect 14792 2985 14848 3041
rect 14576 2891 14632 2947
rect 14684 2891 14740 2947
rect 14792 2891 14848 2947
rect 37308 3805 37364 3861
rect 37402 3805 37458 3861
rect 37496 3805 37552 3861
rect 37308 3717 37364 3773
rect 37402 3717 37458 3773
rect 37496 3717 37552 3773
rect 37308 3629 37364 3685
rect 37402 3629 37458 3685
rect 37496 3629 37552 3685
rect 31271 3105 31327 3161
rect 31396 3105 31452 3161
rect 31521 3105 31577 3161
rect 31271 3009 31327 3065
rect 31396 3009 31452 3065
rect 31521 3009 31577 3065
rect 46942 2958 46998 3014
rect 47035 2958 47091 3014
rect 47128 2958 47184 3014
rect 47221 2958 47277 3014
rect 46942 2876 46998 2932
rect 47035 2876 47091 2932
rect 47128 2876 47184 2932
rect 47221 2876 47277 2932
rect 54255 3350 54311 3406
rect 54359 3350 54415 3406
rect 54463 3350 54519 3406
rect 54567 3350 54623 3406
rect 54255 3260 54311 3316
rect 54359 3260 54415 3316
rect 54463 3260 54519 3316
rect 54567 3260 54623 3316
<< metal3 >>
rect 3425 7602 3531 7619
rect 3425 7538 3446 7602
rect 3510 7538 3531 7602
rect 3425 7522 3531 7538
rect 3425 7458 3446 7522
rect 3510 7458 3531 7522
rect 3425 7441 3531 7458
rect 3634 7601 3740 7618
rect 3634 7537 3655 7601
rect 3719 7537 3740 7601
rect 3634 7521 3740 7537
rect 3634 7457 3655 7521
rect 3719 7457 3740 7521
rect 3634 7440 3740 7457
rect 3800 7601 3906 7618
rect 3800 7537 3821 7601
rect 3885 7537 3906 7601
rect 3800 7521 3906 7537
rect 3800 7457 3821 7521
rect 3885 7457 3906 7521
rect 3800 7440 3906 7457
rect 3980 7603 4086 7620
rect 3980 7539 4001 7603
rect 4065 7539 4086 7603
rect 3980 7523 4086 7539
rect 3980 7459 4001 7523
rect 4065 7459 4086 7523
rect 3980 7442 4086 7459
rect 20054 7619 20160 7636
rect 20054 7555 20075 7619
rect 20139 7555 20160 7619
rect 20054 7539 20160 7555
rect 20054 7475 20075 7539
rect 20139 7475 20160 7539
rect 20054 7458 20160 7475
rect 20270 7619 20376 7636
rect 20270 7555 20291 7619
rect 20355 7555 20376 7619
rect 20270 7539 20376 7555
rect 20270 7475 20291 7539
rect 20355 7475 20376 7539
rect 20270 7458 20376 7475
rect 20486 7619 20592 7636
rect 20486 7555 20507 7619
rect 20571 7555 20592 7619
rect 20486 7539 20592 7555
rect 20486 7475 20507 7539
rect 20571 7475 20592 7539
rect 20486 7458 20592 7475
rect 28546 7618 28652 7635
rect 28546 7554 28567 7618
rect 28631 7554 28652 7618
rect 28546 7538 28652 7554
rect 28546 7474 28567 7538
rect 28631 7474 28652 7538
rect 28546 7457 28652 7474
rect 28762 7618 28868 7635
rect 28762 7554 28783 7618
rect 28847 7554 28868 7618
rect 28762 7538 28868 7554
rect 28762 7474 28783 7538
rect 28847 7474 28868 7538
rect 28762 7457 28868 7474
rect 28978 7618 29084 7635
rect 28978 7554 28999 7618
rect 29063 7554 29084 7618
rect 28978 7538 29084 7554
rect 28978 7474 28999 7538
rect 29063 7474 29084 7538
rect 28978 7457 29084 7474
rect 42074 7624 42180 7641
rect 42074 7560 42095 7624
rect 42159 7560 42180 7624
rect 42074 7544 42180 7560
rect 42074 7480 42095 7544
rect 42159 7480 42180 7544
rect 42074 7463 42180 7480
rect 42290 7624 42396 7641
rect 42290 7560 42311 7624
rect 42375 7560 42396 7624
rect 42290 7544 42396 7560
rect 42290 7480 42311 7544
rect 42375 7480 42396 7544
rect 42290 7463 42396 7480
rect 42506 7624 42612 7641
rect 42506 7560 42527 7624
rect 42591 7560 42612 7624
rect 42506 7544 42612 7560
rect 42506 7480 42527 7544
rect 42591 7480 42612 7544
rect 42506 7463 42612 7480
rect 58559 7617 58665 7634
rect 58559 7553 58580 7617
rect 58644 7553 58665 7617
rect 58559 7537 58665 7553
rect 58559 7473 58580 7537
rect 58644 7473 58665 7537
rect 58559 7456 58665 7473
rect 58775 7617 58881 7634
rect 58775 7553 58796 7617
rect 58860 7553 58881 7617
rect 58775 7537 58881 7553
rect 58775 7473 58796 7537
rect 58860 7473 58881 7537
rect 58775 7456 58881 7473
rect 58991 7617 59097 7634
rect 58991 7553 59012 7617
rect 59076 7553 59097 7617
rect 58991 7537 59097 7553
rect 58991 7473 59012 7537
rect 59076 7473 59097 7537
rect 58991 7456 59097 7473
rect 18519 5505 18625 5522
rect 2191 5484 2297 5501
rect 2191 5420 2212 5484
rect 2276 5420 2297 5484
rect 2191 5404 2297 5420
rect 2191 5340 2212 5404
rect 2276 5340 2297 5404
rect 2191 5323 2297 5340
rect 2363 5485 2469 5502
rect 2363 5421 2384 5485
rect 2448 5421 2469 5485
rect 2363 5405 2469 5421
rect 2363 5341 2384 5405
rect 2448 5341 2469 5405
rect 2363 5324 2469 5341
rect 2537 5484 2643 5501
rect 2537 5420 2558 5484
rect 2622 5420 2643 5484
rect 2537 5404 2643 5420
rect 2537 5340 2558 5404
rect 2622 5340 2643 5404
rect 18519 5441 18540 5505
rect 18604 5441 18625 5505
rect 18519 5425 18625 5441
rect 18519 5361 18540 5425
rect 18604 5361 18625 5425
rect 18519 5344 18625 5361
rect 18735 5505 18841 5522
rect 18735 5441 18756 5505
rect 18820 5441 18841 5505
rect 18735 5425 18841 5441
rect 18735 5361 18756 5425
rect 18820 5361 18841 5425
rect 18735 5344 18841 5361
rect 18951 5505 19057 5522
rect 18951 5441 18972 5505
rect 19036 5441 19057 5505
rect 18951 5425 19057 5441
rect 18951 5361 18972 5425
rect 19036 5361 19057 5425
rect 18951 5344 19057 5361
rect 27027 5497 27133 5514
rect 27027 5433 27048 5497
rect 27112 5433 27133 5497
rect 27027 5417 27133 5433
rect 27027 5353 27048 5417
rect 27112 5353 27133 5417
rect 2537 5323 2643 5340
rect 27027 5336 27133 5353
rect 27243 5497 27349 5514
rect 27243 5433 27264 5497
rect 27328 5433 27349 5497
rect 27243 5417 27349 5433
rect 27243 5353 27264 5417
rect 27328 5353 27349 5417
rect 27243 5336 27349 5353
rect 27459 5497 27565 5514
rect 27459 5433 27480 5497
rect 27544 5433 27565 5497
rect 27459 5417 27565 5433
rect 27459 5353 27480 5417
rect 27544 5353 27565 5417
rect 27459 5336 27565 5353
rect 40499 5492 40605 5509
rect 40499 5428 40520 5492
rect 40584 5428 40605 5492
rect 40499 5412 40605 5428
rect 40499 5348 40520 5412
rect 40584 5348 40605 5412
rect 40499 5331 40605 5348
rect 40715 5492 40821 5509
rect 40715 5428 40736 5492
rect 40800 5428 40821 5492
rect 40715 5412 40821 5428
rect 40715 5348 40736 5412
rect 40800 5348 40821 5412
rect 40715 5331 40821 5348
rect 40931 5492 41037 5509
rect 40931 5428 40952 5492
rect 41016 5428 41037 5492
rect 40931 5412 41037 5428
rect 40931 5348 40952 5412
rect 41016 5348 41037 5412
rect 40931 5331 41037 5348
rect 57050 5484 57156 5501
rect 57050 5420 57071 5484
rect 57135 5420 57156 5484
rect 57050 5404 57156 5420
rect 57050 5340 57071 5404
rect 57135 5340 57156 5404
rect 57050 5323 57156 5340
rect 57266 5484 57372 5501
rect 57266 5420 57287 5484
rect 57351 5420 57372 5484
rect 57266 5404 57372 5420
rect 57266 5340 57287 5404
rect 57351 5340 57372 5404
rect 57266 5323 57372 5340
rect 57482 5484 57588 5501
rect 57482 5420 57503 5484
rect 57567 5420 57588 5484
rect 57482 5404 57588 5420
rect 57482 5340 57503 5404
rect 57567 5340 57588 5404
rect 57482 5323 57588 5340
rect 37285 3861 37589 3875
rect 37285 3805 37308 3861
rect 37364 3805 37402 3861
rect 37458 3805 37496 3861
rect 37552 3805 37589 3861
rect 37285 3773 37589 3805
rect 37285 3717 37308 3773
rect 37364 3738 37402 3773
rect 37396 3717 37402 3738
rect 37458 3739 37496 3773
rect 37458 3717 37486 3739
rect 37552 3717 37589 3773
rect 37285 3685 37332 3717
rect 37396 3685 37486 3717
rect 37550 3685 37589 3717
rect 7181 3628 7523 3661
rect 37285 3629 37308 3685
rect 37396 3674 37402 3685
rect 37364 3629 37402 3674
rect 37458 3675 37486 3685
rect 37458 3629 37496 3675
rect 37552 3629 37589 3685
rect 7113 3602 7602 3628
rect 37285 3609 37589 3629
rect 7113 3546 7182 3602
rect 7238 3546 7296 3602
rect 7352 3546 7410 3602
rect 7466 3546 7602 3602
rect 7113 3487 7602 3546
rect 7113 3431 7182 3487
rect 7238 3445 7296 3487
rect 7352 3451 7410 3487
rect 7254 3431 7296 3445
rect 7405 3431 7410 3451
rect 7466 3451 7602 3487
rect 7466 3431 7486 3451
rect 7113 3381 7190 3431
rect 7254 3387 7341 3431
rect 7405 3387 7486 3431
rect 7550 3387 7602 3451
rect 7254 3381 7602 3387
rect 7113 3372 7602 3381
rect 7113 3316 7182 3372
rect 7238 3316 7296 3372
rect 7352 3316 7410 3372
rect 7466 3316 7602 3372
rect 7113 3261 7602 3316
rect 22171 3512 22638 3566
rect 22171 3456 22221 3512
rect 22277 3459 22325 3512
rect 22297 3456 22325 3459
rect 22381 3459 22429 3512
rect 22381 3456 22400 3459
rect 22485 3456 22533 3512
rect 22589 3456 22638 3512
rect 22171 3396 22233 3456
rect 22297 3396 22400 3456
rect 22464 3396 22638 3456
rect 22171 3340 22221 3396
rect 22297 3395 22325 3396
rect 22277 3340 22325 3395
rect 22381 3395 22400 3396
rect 22381 3340 22429 3395
rect 22485 3340 22533 3396
rect 22589 3340 22638 3396
rect 22171 3298 22638 3340
rect 22171 3280 22233 3298
rect 22297 3280 22400 3298
rect 22464 3280 22638 3298
rect 22171 3224 22221 3280
rect 22297 3234 22325 3280
rect 22277 3224 22325 3234
rect 22381 3234 22400 3280
rect 22381 3224 22429 3234
rect 22485 3224 22533 3280
rect 22589 3224 22638 3280
rect 54218 3406 54640 3434
rect 54218 3350 54255 3406
rect 54336 3350 54359 3406
rect 54457 3350 54463 3406
rect 54519 3350 54531 3406
rect 54623 3350 54640 3406
rect 54218 3342 54272 3350
rect 54336 3342 54393 3350
rect 54457 3342 54531 3350
rect 54595 3342 54640 3350
rect 54218 3326 54640 3342
rect 54218 3316 54272 3326
rect 54336 3316 54393 3326
rect 54457 3316 54531 3326
rect 54595 3316 54640 3326
rect 54218 3260 54255 3316
rect 54336 3262 54359 3316
rect 54457 3262 54463 3316
rect 54311 3260 54359 3262
rect 54415 3260 54463 3262
rect 54519 3262 54531 3316
rect 54519 3260 54567 3262
rect 54623 3260 54640 3316
rect 54218 3226 54640 3260
rect 22171 3180 22638 3224
rect 31223 3161 31648 3199
rect 31223 3105 31271 3161
rect 31327 3105 31396 3161
rect 31452 3105 31521 3161
rect 31577 3105 31648 3161
rect 31223 3098 31648 3105
rect 31223 3065 31280 3098
rect 31344 3065 31399 3098
rect 14536 3041 14889 3064
rect 14536 2990 14576 3041
rect 14632 2990 14684 3041
rect 14740 2990 14792 3041
rect 14536 2926 14566 2990
rect 14632 2985 14669 2990
rect 14740 2985 14772 2990
rect 14848 2985 14889 3041
rect 14630 2947 14669 2985
rect 14733 2947 14772 2985
rect 14836 2947 14889 2985
rect 31223 3009 31271 3065
rect 31344 3034 31396 3065
rect 31463 3034 31518 3098
rect 31582 3034 31648 3098
rect 31327 3009 31396 3034
rect 31452 3009 31521 3034
rect 31577 3009 31648 3034
rect 31223 2972 31648 3009
rect 46905 3031 47320 3081
rect 46905 3030 47093 3031
rect 46905 3014 46953 3030
rect 47017 3014 47093 3030
rect 47157 3014 47221 3031
rect 14632 2926 14669 2947
rect 14740 2926 14772 2947
rect 14536 2891 14576 2926
rect 14632 2891 14684 2926
rect 14740 2891 14792 2926
rect 14848 2891 14889 2947
rect 14536 2865 14889 2891
rect 46905 2958 46942 3014
rect 47017 2966 47035 3014
rect 46998 2958 47035 2966
rect 47091 2967 47093 3014
rect 47091 2958 47128 2967
rect 47184 2958 47221 3014
rect 47285 2967 47320 3031
rect 47277 2958 47320 2967
rect 46905 2951 47320 2958
rect 46905 2950 47093 2951
rect 46905 2932 46953 2950
rect 47017 2932 47093 2950
rect 47157 2932 47221 2951
rect 46905 2876 46942 2932
rect 47017 2886 47035 2932
rect 46998 2876 47035 2886
rect 47091 2887 47093 2932
rect 47091 2876 47128 2887
rect 47184 2876 47221 2932
rect 47285 2887 47320 2951
rect 47277 2876 47320 2887
rect 46905 2840 47320 2876
rect 2193 2536 2299 2553
rect 2193 2472 2214 2536
rect 2278 2472 2299 2536
rect 2193 2456 2299 2472
rect 2193 2392 2214 2456
rect 2278 2392 2299 2456
rect 2193 2375 2299 2392
rect 2398 2538 2504 2555
rect 2398 2474 2419 2538
rect 2483 2474 2504 2538
rect 2398 2458 2504 2474
rect 2398 2394 2419 2458
rect 2483 2394 2504 2458
rect 2398 2377 2504 2394
rect 2597 2538 2703 2555
rect 2597 2474 2618 2538
rect 2682 2474 2703 2538
rect 2597 2458 2703 2474
rect 2597 2394 2618 2458
rect 2682 2394 2703 2458
rect 2597 2377 2703 2394
rect 18510 2554 18616 2571
rect 18510 2490 18531 2554
rect 18595 2490 18616 2554
rect 18510 2474 18616 2490
rect 18510 2410 18531 2474
rect 18595 2410 18616 2474
rect 18510 2393 18616 2410
rect 18726 2554 18832 2571
rect 18726 2490 18747 2554
rect 18811 2490 18832 2554
rect 18726 2474 18832 2490
rect 18726 2410 18747 2474
rect 18811 2410 18832 2474
rect 18726 2393 18832 2410
rect 18942 2554 19048 2571
rect 18942 2490 18963 2554
rect 19027 2490 19048 2554
rect 18942 2474 19048 2490
rect 18942 2410 18963 2474
rect 19027 2410 19048 2474
rect 18942 2393 19048 2410
rect 27032 2549 27138 2566
rect 27032 2485 27053 2549
rect 27117 2485 27138 2549
rect 27032 2469 27138 2485
rect 27032 2405 27053 2469
rect 27117 2405 27138 2469
rect 27032 2388 27138 2405
rect 27248 2549 27354 2566
rect 27248 2485 27269 2549
rect 27333 2485 27354 2549
rect 27248 2469 27354 2485
rect 27248 2405 27269 2469
rect 27333 2405 27354 2469
rect 27248 2388 27354 2405
rect 27464 2549 27570 2566
rect 27464 2485 27485 2549
rect 27549 2485 27570 2549
rect 27464 2469 27570 2485
rect 27464 2405 27485 2469
rect 27549 2405 27570 2469
rect 27464 2388 27570 2405
rect 40535 2551 40641 2568
rect 40535 2487 40556 2551
rect 40620 2487 40641 2551
rect 40535 2471 40641 2487
rect 40535 2407 40556 2471
rect 40620 2407 40641 2471
rect 40535 2390 40641 2407
rect 40751 2551 40857 2568
rect 40751 2487 40772 2551
rect 40836 2487 40857 2551
rect 40751 2471 40857 2487
rect 40751 2407 40772 2471
rect 40836 2407 40857 2471
rect 40751 2390 40857 2407
rect 40967 2551 41073 2568
rect 40967 2487 40988 2551
rect 41052 2487 41073 2551
rect 40967 2471 41073 2487
rect 40967 2407 40988 2471
rect 41052 2407 41073 2471
rect 40967 2390 41073 2407
rect 57030 2562 57136 2579
rect 57030 2498 57051 2562
rect 57115 2498 57136 2562
rect 57030 2482 57136 2498
rect 57030 2418 57051 2482
rect 57115 2418 57136 2482
rect 57030 2401 57136 2418
rect 57246 2562 57352 2579
rect 57246 2498 57267 2562
rect 57331 2498 57352 2562
rect 57246 2482 57352 2498
rect 57246 2418 57267 2482
rect 57331 2418 57352 2482
rect 57246 2401 57352 2418
rect 57462 2562 57568 2579
rect 57462 2498 57483 2562
rect 57547 2498 57568 2562
rect 57462 2482 57568 2498
rect 57462 2418 57483 2482
rect 57547 2418 57568 2482
rect 57462 2401 57568 2418
rect 3439 425 3545 442
rect 3439 361 3460 425
rect 3524 361 3545 425
rect 3439 345 3545 361
rect 3439 281 3460 345
rect 3524 281 3545 345
rect 3439 264 3545 281
rect 3660 425 3766 442
rect 3660 361 3681 425
rect 3745 361 3766 425
rect 3660 345 3766 361
rect 3660 281 3681 345
rect 3745 281 3766 345
rect 3660 264 3766 281
rect 3869 425 3975 442
rect 3869 361 3890 425
rect 3954 361 3975 425
rect 3869 345 3975 361
rect 3869 281 3890 345
rect 3954 281 3975 345
rect 3869 264 3975 281
rect 4043 425 4149 442
rect 4043 361 4064 425
rect 4128 361 4149 425
rect 14686 436 14763 439
rect 4043 345 4149 361
rect 4043 281 4064 345
rect 4128 281 4149 345
rect 7167 373 7253 387
rect 7167 309 7178 373
rect 7242 309 7253 373
rect 7167 296 7253 309
rect 7315 373 7401 387
rect 7315 309 7326 373
rect 7390 309 7401 373
rect 7315 296 7401 309
rect 7463 373 7549 387
rect 7463 309 7474 373
rect 7538 309 7549 373
rect 14686 372 14692 436
rect 14756 372 14763 436
rect 14686 370 14763 372
rect 20072 424 20178 441
rect 20072 360 20093 424
rect 20157 360 20178 424
rect 20072 344 20178 360
rect 7463 296 7549 309
rect 14709 317 14786 320
rect 4043 264 4149 281
rect 14709 253 14715 317
rect 14779 253 14786 317
rect 20072 280 20093 344
rect 20157 280 20178 344
rect 20072 263 20178 280
rect 20288 424 20394 441
rect 20288 360 20309 424
rect 20373 360 20394 424
rect 20288 344 20394 360
rect 20288 280 20309 344
rect 20373 280 20394 344
rect 20288 263 20394 280
rect 20504 424 20610 441
rect 20504 360 20525 424
rect 20589 360 20610 424
rect 28501 429 28607 446
rect 20504 344 20610 360
rect 20504 280 20525 344
rect 20589 280 20610 344
rect 22224 377 22320 399
rect 22224 313 22240 377
rect 22304 313 22320 377
rect 22224 291 22320 313
rect 22357 377 22453 399
rect 22357 313 22373 377
rect 22437 313 22453 377
rect 22357 291 22453 313
rect 22490 377 22586 399
rect 22490 313 22506 377
rect 22570 313 22586 377
rect 22490 291 22586 313
rect 28501 365 28522 429
rect 28586 365 28607 429
rect 28501 349 28607 365
rect 20504 263 20610 280
rect 28501 285 28522 349
rect 28586 285 28607 349
rect 28501 268 28607 285
rect 28717 429 28823 446
rect 28717 365 28738 429
rect 28802 365 28823 429
rect 28717 349 28823 365
rect 28717 285 28738 349
rect 28802 285 28823 349
rect 28717 268 28823 285
rect 28933 429 29039 446
rect 28933 365 28954 429
rect 29018 365 29039 429
rect 42019 419 42125 436
rect 28933 349 29039 365
rect 28933 285 28954 349
rect 29018 285 29039 349
rect 28933 268 29039 285
rect 31290 366 31377 390
rect 31290 302 31301 366
rect 31365 302 31377 366
rect 31290 278 31377 302
rect 31413 366 31500 390
rect 31413 302 31424 366
rect 31488 302 31500 366
rect 31413 278 31500 302
rect 31545 366 31632 390
rect 31545 302 31556 366
rect 31620 302 31632 366
rect 31545 278 31632 302
rect 37319 363 37406 387
rect 37319 299 37330 363
rect 37394 299 37406 363
rect 37319 275 37406 299
rect 37488 363 37575 387
rect 37488 299 37499 363
rect 37563 299 37575 363
rect 37488 275 37575 299
rect 42019 355 42040 419
rect 42104 355 42125 419
rect 42019 339 42125 355
rect 42019 275 42040 339
rect 42104 275 42125 339
rect 42019 258 42125 275
rect 42235 419 42341 436
rect 42235 355 42256 419
rect 42320 355 42341 419
rect 42235 339 42341 355
rect 42235 275 42256 339
rect 42320 275 42341 339
rect 42235 258 42341 275
rect 42451 419 42557 436
rect 54268 423 54352 430
rect 42451 355 42472 419
rect 42536 355 42557 419
rect 42451 339 42557 355
rect 42451 275 42472 339
rect 42536 275 42557 339
rect 42451 258 42557 275
rect 46945 413 47029 420
rect 46945 349 46955 413
rect 47019 349 47029 413
rect 46945 333 47029 349
rect 46945 269 46955 333
rect 47019 269 47029 333
rect 46945 262 47029 269
rect 47058 413 47142 420
rect 47058 349 47068 413
rect 47132 349 47142 413
rect 47058 333 47142 349
rect 47058 269 47068 333
rect 47132 269 47142 333
rect 47058 262 47142 269
rect 47173 413 47257 420
rect 47173 349 47183 413
rect 47247 349 47257 413
rect 47173 333 47257 349
rect 47173 269 47183 333
rect 47247 269 47257 333
rect 54268 359 54278 423
rect 54342 359 54352 423
rect 54268 343 54352 359
rect 54268 279 54278 343
rect 54342 279 54352 343
rect 54268 272 54352 279
rect 54387 423 54471 430
rect 54387 359 54397 423
rect 54461 359 54471 423
rect 54387 343 54471 359
rect 54387 279 54397 343
rect 54461 279 54471 343
rect 54387 272 54471 279
rect 54516 423 54600 430
rect 54516 359 54526 423
rect 54590 359 54600 423
rect 54516 343 54600 359
rect 54516 279 54526 343
rect 54590 279 54600 343
rect 54516 272 54600 279
rect 58531 414 58637 431
rect 58531 350 58552 414
rect 58616 350 58637 414
rect 58531 334 58637 350
rect 47173 262 47257 269
rect 58531 270 58552 334
rect 58616 270 58637 334
rect 58531 253 58637 270
rect 58747 414 58853 431
rect 58747 350 58768 414
rect 58832 350 58853 414
rect 58747 334 58853 350
rect 58747 270 58768 334
rect 58832 270 58853 334
rect 58747 253 58853 270
rect 58963 414 59069 431
rect 58963 350 58984 414
rect 59048 350 59069 414
rect 58963 334 59069 350
rect 58963 270 58984 334
rect 59048 270 59069 334
rect 58963 253 59069 270
rect 14709 251 14786 253
<< via3 >>
rect 3446 7538 3510 7602
rect 3446 7458 3510 7522
rect 3655 7537 3719 7601
rect 3655 7457 3719 7521
rect 3821 7537 3885 7601
rect 3821 7457 3885 7521
rect 4001 7539 4065 7603
rect 4001 7459 4065 7523
rect 20075 7555 20139 7619
rect 20075 7475 20139 7539
rect 20291 7555 20355 7619
rect 20291 7475 20355 7539
rect 20507 7555 20571 7619
rect 20507 7475 20571 7539
rect 28567 7554 28631 7618
rect 28567 7474 28631 7538
rect 28783 7554 28847 7618
rect 28783 7474 28847 7538
rect 28999 7554 29063 7618
rect 28999 7474 29063 7538
rect 42095 7560 42159 7624
rect 42095 7480 42159 7544
rect 42311 7560 42375 7624
rect 42311 7480 42375 7544
rect 42527 7560 42591 7624
rect 42527 7480 42591 7544
rect 58580 7553 58644 7617
rect 58580 7473 58644 7537
rect 58796 7553 58860 7617
rect 58796 7473 58860 7537
rect 59012 7553 59076 7617
rect 59012 7473 59076 7537
rect 2212 5420 2276 5484
rect 2212 5340 2276 5404
rect 2384 5421 2448 5485
rect 2384 5341 2448 5405
rect 2558 5420 2622 5484
rect 2558 5340 2622 5404
rect 18540 5441 18604 5505
rect 18540 5361 18604 5425
rect 18756 5441 18820 5505
rect 18756 5361 18820 5425
rect 18972 5441 19036 5505
rect 18972 5361 19036 5425
rect 27048 5433 27112 5497
rect 27048 5353 27112 5417
rect 27264 5433 27328 5497
rect 27264 5353 27328 5417
rect 27480 5433 27544 5497
rect 27480 5353 27544 5417
rect 40520 5428 40584 5492
rect 40520 5348 40584 5412
rect 40736 5428 40800 5492
rect 40736 5348 40800 5412
rect 40952 5428 41016 5492
rect 40952 5348 41016 5412
rect 57071 5420 57135 5484
rect 57071 5340 57135 5404
rect 57287 5420 57351 5484
rect 57287 5340 57351 5404
rect 57503 5420 57567 5484
rect 57503 5340 57567 5404
rect 37332 3717 37364 3738
rect 37364 3717 37396 3738
rect 37486 3717 37496 3739
rect 37496 3717 37550 3739
rect 37332 3685 37396 3717
rect 37486 3685 37550 3717
rect 37332 3674 37364 3685
rect 37364 3674 37396 3685
rect 37486 3675 37496 3685
rect 37496 3675 37550 3685
rect 7190 3431 7238 3445
rect 7238 3431 7254 3445
rect 7341 3431 7352 3451
rect 7352 3431 7405 3451
rect 7190 3381 7254 3431
rect 7341 3387 7405 3431
rect 7486 3387 7550 3451
rect 22233 3456 22277 3459
rect 22277 3456 22297 3459
rect 22400 3456 22429 3459
rect 22429 3456 22464 3459
rect 22233 3396 22297 3456
rect 22400 3396 22464 3456
rect 22233 3395 22277 3396
rect 22277 3395 22297 3396
rect 22400 3395 22429 3396
rect 22429 3395 22464 3396
rect 22233 3280 22297 3298
rect 22400 3280 22464 3298
rect 22233 3234 22277 3280
rect 22277 3234 22297 3280
rect 22400 3234 22429 3280
rect 22429 3234 22464 3280
rect 54272 3350 54311 3406
rect 54311 3350 54336 3406
rect 54393 3350 54415 3406
rect 54415 3350 54457 3406
rect 54531 3350 54567 3406
rect 54567 3350 54595 3406
rect 54272 3342 54336 3350
rect 54393 3342 54457 3350
rect 54531 3342 54595 3350
rect 54272 3316 54336 3326
rect 54393 3316 54457 3326
rect 54531 3316 54595 3326
rect 54272 3262 54311 3316
rect 54311 3262 54336 3316
rect 54393 3262 54415 3316
rect 54415 3262 54457 3316
rect 54531 3262 54567 3316
rect 54567 3262 54595 3316
rect 31280 3065 31344 3098
rect 31399 3065 31463 3098
rect 14566 2985 14576 2990
rect 14576 2985 14630 2990
rect 14669 2985 14684 2990
rect 14684 2985 14733 2990
rect 14772 2985 14792 2990
rect 14792 2985 14836 2990
rect 14566 2947 14630 2985
rect 14669 2947 14733 2985
rect 14772 2947 14836 2985
rect 31280 3034 31327 3065
rect 31327 3034 31344 3065
rect 31399 3034 31452 3065
rect 31452 3034 31463 3065
rect 31518 3065 31582 3098
rect 31518 3034 31521 3065
rect 31521 3034 31577 3065
rect 31577 3034 31582 3065
rect 46953 3014 47017 3030
rect 47093 3014 47157 3031
rect 47221 3014 47285 3031
rect 14566 2926 14576 2947
rect 14576 2926 14630 2947
rect 14669 2926 14684 2947
rect 14684 2926 14733 2947
rect 14772 2926 14792 2947
rect 14792 2926 14836 2947
rect 46953 2966 46998 3014
rect 46998 2966 47017 3014
rect 47093 2967 47128 3014
rect 47128 2967 47157 3014
rect 47221 2967 47277 3014
rect 47277 2967 47285 3014
rect 46953 2932 47017 2950
rect 47093 2932 47157 2951
rect 47221 2932 47285 2951
rect 46953 2886 46998 2932
rect 46998 2886 47017 2932
rect 47093 2887 47128 2932
rect 47128 2887 47157 2932
rect 47221 2887 47277 2932
rect 47277 2887 47285 2932
rect 2214 2472 2278 2536
rect 2214 2392 2278 2456
rect 2419 2474 2483 2538
rect 2419 2394 2483 2458
rect 2618 2474 2682 2538
rect 2618 2394 2682 2458
rect 18531 2490 18595 2554
rect 18531 2410 18595 2474
rect 18747 2490 18811 2554
rect 18747 2410 18811 2474
rect 18963 2490 19027 2554
rect 18963 2410 19027 2474
rect 27053 2485 27117 2549
rect 27053 2405 27117 2469
rect 27269 2485 27333 2549
rect 27269 2405 27333 2469
rect 27485 2485 27549 2549
rect 27485 2405 27549 2469
rect 40556 2487 40620 2551
rect 40556 2407 40620 2471
rect 40772 2487 40836 2551
rect 40772 2407 40836 2471
rect 40988 2487 41052 2551
rect 40988 2407 41052 2471
rect 57051 2498 57115 2562
rect 57051 2418 57115 2482
rect 57267 2498 57331 2562
rect 57267 2418 57331 2482
rect 57483 2498 57547 2562
rect 57483 2418 57547 2482
rect 3460 361 3524 425
rect 3460 281 3524 345
rect 3681 361 3745 425
rect 3681 281 3745 345
rect 3890 361 3954 425
rect 3890 281 3954 345
rect 4064 361 4128 425
rect 4064 281 4128 345
rect 7178 309 7242 373
rect 7326 309 7390 373
rect 7474 309 7538 373
rect 14692 372 14756 436
rect 20093 360 20157 424
rect 14715 253 14779 317
rect 20093 280 20157 344
rect 20309 360 20373 424
rect 20309 280 20373 344
rect 20525 360 20589 424
rect 20525 280 20589 344
rect 22240 313 22304 377
rect 22373 313 22437 377
rect 22506 313 22570 377
rect 28522 365 28586 429
rect 28522 285 28586 349
rect 28738 365 28802 429
rect 28738 285 28802 349
rect 28954 365 29018 429
rect 28954 285 29018 349
rect 31301 302 31365 366
rect 31424 302 31488 366
rect 31556 302 31620 366
rect 37330 299 37394 363
rect 37499 299 37563 363
rect 42040 355 42104 419
rect 42040 275 42104 339
rect 42256 355 42320 419
rect 42256 275 42320 339
rect 42472 355 42536 419
rect 42472 275 42536 339
rect 46955 349 47019 413
rect 46955 269 47019 333
rect 47068 349 47132 413
rect 47068 269 47132 333
rect 47183 349 47247 413
rect 47183 269 47247 333
rect 54278 359 54342 423
rect 54278 279 54342 343
rect 54397 359 54461 423
rect 54397 279 54461 343
rect 54526 359 54590 423
rect 54526 279 54590 343
rect 58552 350 58616 414
rect 58552 270 58616 334
rect 58768 350 58832 414
rect 58768 270 58832 334
rect 58984 350 59048 414
rect 58984 270 59048 334
<< metal4 >>
rect 2047 5485 2853 7801
rect 2047 5484 2384 5485
rect 2047 5420 2212 5484
rect 2276 5421 2384 5484
rect 2448 5484 2853 5485
rect 2448 5421 2558 5484
rect 2276 5420 2558 5421
rect 2622 5420 2853 5484
rect 2047 5405 2853 5420
rect 2047 5404 2384 5405
rect 2047 5340 2212 5404
rect 2276 5341 2384 5404
rect 2448 5404 2853 5405
rect 2448 5341 2558 5404
rect 2276 5340 2558 5341
rect 2622 5340 2853 5404
rect 2047 2538 2853 5340
rect 2047 2536 2419 2538
rect 2047 2472 2214 2536
rect 2278 2474 2419 2536
rect 2483 2474 2618 2538
rect 2682 2474 2853 2538
rect 2278 2472 2853 2474
rect 2047 2458 2853 2472
rect 2047 2456 2419 2458
rect 2047 2392 2214 2456
rect 2278 2394 2419 2456
rect 2483 2394 2618 2458
rect 2682 2394 2853 2458
rect 2278 2392 2853 2394
rect 2047 95 2853 2392
rect 3390 7603 4196 7802
rect 3390 7602 4001 7603
rect 3390 7538 3446 7602
rect 3510 7601 4001 7602
rect 3510 7538 3655 7601
rect 3390 7537 3655 7538
rect 3719 7537 3821 7601
rect 3885 7539 4001 7601
rect 4065 7539 4196 7603
rect 3885 7537 4196 7539
rect 3390 7523 4196 7537
rect 3390 7522 4001 7523
rect 3390 7458 3446 7522
rect 3510 7521 4001 7522
rect 3510 7458 3655 7521
rect 3390 7457 3655 7458
rect 3719 7457 3821 7521
rect 3885 7459 4001 7521
rect 4065 7459 4196 7523
rect 3885 7457 4196 7459
rect 3390 425 4196 7457
rect 18390 5505 19196 7802
rect 18390 5441 18540 5505
rect 18604 5441 18756 5505
rect 18820 5441 18972 5505
rect 19036 5441 19196 5505
rect 18390 5425 19196 5441
rect 18390 5361 18540 5425
rect 18604 5361 18756 5425
rect 18820 5361 18972 5425
rect 19036 5361 19196 5425
rect 3390 361 3460 425
rect 3524 361 3681 425
rect 3745 361 3890 425
rect 3954 361 4064 425
rect 4128 361 4196 425
rect 3390 345 4196 361
rect 3390 281 3460 345
rect 3524 281 3681 345
rect 3745 281 3890 345
rect 3954 281 4064 345
rect 4128 281 4196 345
rect 3390 96 4196 281
rect 7121 3451 7590 3580
rect 7121 3445 7341 3451
rect 7121 3381 7190 3445
rect 7254 3387 7341 3445
rect 7405 3387 7486 3451
rect 7550 3387 7590 3451
rect 7254 3381 7590 3387
rect 7121 373 7590 3381
rect 14536 2990 14890 3065
rect 14536 2926 14566 2990
rect 14630 2926 14669 2990
rect 14733 2926 14772 2990
rect 14836 2926 14890 2990
rect 14536 2864 14890 2926
rect 7121 309 7178 373
rect 7242 309 7326 373
rect 7390 309 7474 373
rect 7538 309 7590 373
rect 7121 197 7590 309
rect 14612 436 14813 2864
rect 14612 372 14692 436
rect 14756 372 14813 436
rect 14612 317 14813 372
rect 14612 253 14715 317
rect 14779 253 14813 317
rect 14612 172 14813 253
rect 18390 2554 19196 5361
rect 18390 2490 18531 2554
rect 18595 2490 18747 2554
rect 18811 2490 18963 2554
rect 19027 2490 19196 2554
rect 18390 2474 19196 2490
rect 18390 2410 18531 2474
rect 18595 2410 18747 2474
rect 18811 2410 18963 2474
rect 19027 2410 19196 2474
rect 18390 96 19196 2410
rect 19890 7619 20696 7802
rect 19890 7555 20075 7619
rect 20139 7555 20291 7619
rect 20355 7555 20507 7619
rect 20571 7555 20696 7619
rect 19890 7539 20696 7555
rect 19890 7475 20075 7539
rect 20139 7475 20291 7539
rect 20355 7475 20507 7539
rect 20571 7475 20696 7539
rect 19890 424 20696 7475
rect 26890 5497 27696 7802
rect 26890 5433 27048 5497
rect 27112 5433 27264 5497
rect 27328 5433 27480 5497
rect 27544 5433 27696 5497
rect 26890 5417 27696 5433
rect 26890 5353 27048 5417
rect 27112 5353 27264 5417
rect 27328 5353 27480 5417
rect 27544 5353 27696 5417
rect 19890 360 20093 424
rect 20157 360 20309 424
rect 20373 360 20525 424
rect 20589 360 20696 424
rect 19890 344 20696 360
rect 19890 280 20093 344
rect 20157 280 20309 344
rect 20373 280 20525 344
rect 20589 280 20696 344
rect 19890 96 20696 280
rect 22171 3459 22638 3594
rect 22171 3395 22233 3459
rect 22297 3395 22400 3459
rect 22464 3395 22638 3459
rect 22171 3298 22638 3395
rect 22171 3234 22233 3298
rect 22297 3234 22400 3298
rect 22464 3234 22638 3298
rect 22171 377 22638 3234
rect 22171 313 22240 377
rect 22304 313 22373 377
rect 22437 313 22506 377
rect 22570 313 22638 377
rect 22171 222 22638 313
rect 26890 2549 27696 5353
rect 26890 2485 27053 2549
rect 27117 2485 27269 2549
rect 27333 2485 27485 2549
rect 27549 2485 27696 2549
rect 26890 2469 27696 2485
rect 26890 2405 27053 2469
rect 27117 2405 27269 2469
rect 27333 2405 27485 2469
rect 27549 2405 27696 2469
rect 26890 96 27696 2405
rect 28390 7618 29196 7802
rect 28390 7554 28567 7618
rect 28631 7554 28783 7618
rect 28847 7554 28999 7618
rect 29063 7554 29196 7618
rect 28390 7538 29196 7554
rect 28390 7474 28567 7538
rect 28631 7474 28783 7538
rect 28847 7474 28999 7538
rect 29063 7474 29196 7538
rect 28390 429 29196 7474
rect 40390 5492 41196 7802
rect 40390 5428 40520 5492
rect 40584 5428 40736 5492
rect 40800 5428 40952 5492
rect 41016 5428 41196 5492
rect 40390 5412 41196 5428
rect 40390 5348 40520 5412
rect 40584 5348 40736 5412
rect 40800 5348 40952 5412
rect 41016 5348 41196 5412
rect 37285 3739 37590 3920
rect 37285 3738 37486 3739
rect 37285 3674 37332 3738
rect 37396 3675 37486 3738
rect 37550 3675 37590 3739
rect 37396 3674 37590 3675
rect 28390 365 28522 429
rect 28586 365 28738 429
rect 28802 365 28954 429
rect 29018 365 29196 429
rect 28390 349 29196 365
rect 28390 285 28522 349
rect 28586 285 28738 349
rect 28802 285 28954 349
rect 29018 285 29196 349
rect 28390 96 29196 285
rect 31223 3098 31648 3201
rect 31223 3034 31280 3098
rect 31344 3034 31399 3098
rect 31463 3034 31518 3098
rect 31582 3034 31648 3098
rect 31223 366 31648 3034
rect 31223 302 31301 366
rect 31365 302 31424 366
rect 31488 302 31556 366
rect 31620 302 31648 366
rect 31223 236 31648 302
rect 37285 363 37590 3674
rect 37285 299 37330 363
rect 37394 299 37499 363
rect 37563 299 37590 363
rect 37285 227 37590 299
rect 40390 2551 41196 5348
rect 40390 2487 40556 2551
rect 40620 2487 40772 2551
rect 40836 2487 40988 2551
rect 41052 2487 41196 2551
rect 40390 2471 41196 2487
rect 40390 2407 40556 2471
rect 40620 2407 40772 2471
rect 40836 2407 40988 2471
rect 41052 2407 41196 2471
rect 40390 96 41196 2407
rect 41890 7624 42696 7802
rect 41890 7560 42095 7624
rect 42159 7560 42311 7624
rect 42375 7560 42527 7624
rect 42591 7560 42696 7624
rect 41890 7544 42696 7560
rect 41890 7480 42095 7544
rect 42159 7480 42311 7544
rect 42375 7480 42527 7544
rect 42591 7480 42696 7544
rect 41890 419 42696 7480
rect 56890 5484 57696 7802
rect 56890 5420 57071 5484
rect 57135 5420 57287 5484
rect 57351 5420 57503 5484
rect 57567 5420 57696 5484
rect 56890 5404 57696 5420
rect 56890 5340 57071 5404
rect 57135 5340 57287 5404
rect 57351 5340 57503 5404
rect 57567 5340 57696 5404
rect 54218 3406 54643 3436
rect 54218 3342 54272 3406
rect 54336 3342 54393 3406
rect 54457 3342 54531 3406
rect 54595 3342 54643 3406
rect 54218 3326 54643 3342
rect 54218 3262 54272 3326
rect 54336 3262 54393 3326
rect 54457 3262 54531 3326
rect 54595 3262 54643 3326
rect 41890 355 42040 419
rect 42104 355 42256 419
rect 42320 355 42472 419
rect 42536 355 42696 419
rect 41890 339 42696 355
rect 41890 275 42040 339
rect 42104 275 42256 339
rect 42320 275 42472 339
rect 42536 275 42696 339
rect 41890 96 42696 275
rect 46905 3031 47319 3127
rect 46905 3030 47093 3031
rect 46905 2966 46953 3030
rect 47017 2967 47093 3030
rect 47157 2967 47221 3031
rect 47285 2967 47319 3031
rect 47017 2966 47319 2967
rect 46905 2951 47319 2966
rect 46905 2950 47093 2951
rect 46905 2886 46953 2950
rect 47017 2887 47093 2950
rect 47157 2887 47221 2951
rect 47285 2887 47319 2951
rect 47017 2886 47319 2887
rect 46905 413 47319 2886
rect 46905 349 46955 413
rect 47019 349 47068 413
rect 47132 349 47183 413
rect 47247 349 47319 413
rect 46905 333 47319 349
rect 46905 269 46955 333
rect 47019 269 47068 333
rect 47132 269 47183 333
rect 47247 269 47319 333
rect 46905 174 47319 269
rect 54218 423 54643 3262
rect 54218 359 54278 423
rect 54342 359 54397 423
rect 54461 359 54526 423
rect 54590 359 54643 423
rect 54218 343 54643 359
rect 54218 279 54278 343
rect 54342 279 54397 343
rect 54461 279 54526 343
rect 54590 279 54643 343
rect 54218 186 54643 279
rect 56890 2562 57696 5340
rect 56890 2498 57051 2562
rect 57115 2498 57267 2562
rect 57331 2498 57483 2562
rect 57547 2498 57696 2562
rect 56890 2482 57696 2498
rect 56890 2418 57051 2482
rect 57115 2418 57267 2482
rect 57331 2418 57483 2482
rect 57547 2418 57696 2482
rect 56890 96 57696 2418
rect 58390 7617 59196 7802
rect 58390 7553 58580 7617
rect 58644 7553 58796 7617
rect 58860 7553 59012 7617
rect 59076 7553 59196 7617
rect 58390 7537 59196 7553
rect 58390 7473 58580 7537
rect 58644 7473 58796 7537
rect 58860 7473 59012 7537
rect 59076 7473 59196 7537
rect 58390 414 59196 7473
rect 58390 350 58552 414
rect 58616 350 58768 414
rect 58832 350 58984 414
rect 59048 350 59196 414
rect 58390 334 59196 350
rect 58390 270 58552 334
rect 58616 270 58768 334
rect 58832 270 58984 334
rect 59048 270 59196 334
rect 58390 96 59196 270
use brbufhalf  brbufhalf_0
timestamp 1483428465
transform -1 0 27135 0 -1 10198
box -3552 2527 26658 5446
use brbufhalf  brbufhalf_1
timestamp 1483428465
transform -1 0 57337 0 -1 10198
box -3552 2527 26658 5446
use brbufhalf  brbufhalf_2
timestamp 1483428465
transform 1 0 34661 0 1 -2298
box -3552 2527 26658 5446
use brbufhalf  brbufhalf_3
timestamp 1483428465
transform 1 0 4459 0 1 -2298
box -3552 2527 26658 5446
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0
timestamp 1483428465
transform 1 0 30934 0 1 3801
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0
timestamp 1483428465
transform 1 0 44288 0 1 3585
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1483428465
transform 1 0 46218 0 1 3585
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_2
timestamp 1483428465
transform 1 0 31482 0 1 3801
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_3
timestamp 1483428465
transform 1 0 14146 0 1 3425
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_4
timestamp 1483428465
transform 1 0 16076 0 1 3425
box -38 -48 1510 592
<< labels >>
flabel metal1 s 61289 1010 61511 1088 1 FreeSans 2000 0 0 0 OUT
port 1 nsew
flabel metal1 s 0 4161 254 4227 1 FreeSans 2000 0 0 0 RESET
port 2 nsew
flabel metal4 s 2047 95 2853 7801 1 FreeSans 2000 0 0 0 VDD
port 3 nsew
flabel metal4 s 18390 96 19196 7802 1 FreeSans 2000 0 0 0 VDD
port 3 nsew
flabel metal4 s 26890 96 27696 7802 1 FreeSans 2000 0 0 0 VDD
port 3 nsew
flabel metal4 s 40390 96 41196 7802 1 FreeSans 2000 0 0 0 VDD
port 3 nsew
flabel metal4 s 56890 96 57696 7802 1 FreeSans 2000 0 0 0 VDD
port 3 nsew
flabel metal4 s 3390 96 4196 7802 1 FreeSans 2000 0 0 0 VSS
port 4 nsew
flabel metal4 s 19890 96 20696 7802 1 FreeSans 2000 0 0 0 VSS
port 4 nsew
flabel metal4 s 28390 96 29196 7802 1 FreeSans 2000 0 0 0 VSS
port 4 nsew
flabel metal4 s 41890 96 42696 7802 1 FreeSans 2000 0 0 0 VSS
port 4 nsew
flabel metal4 s 58390 96 59196 7802 1 FreeSans 2000 0 0 0 VSS
port 4 nsew
flabel metal2 s 59455 124 59499 1022 1 FreeSans 2000 0 0 0 C[63]
port 5 nsew
flabel metal2 s 55679 124 55723 1022 1 FreeSans 2000 0 0 0 C[61]
port 6 nsew
flabel metal2 s 53791 124 53835 1022 1 FreeSans 2000 0 0 0 C[60]
port 7 nsew
flabel metal2 s 51903 124 51947 1022 1 FreeSans 2000 0 0 0 C[59]
port 8 nsew
flabel metal2 s 50015 124 50059 1022 1 FreeSans 2000 0 0 0 C[58]
port 9 nsew
flabel metal2 s 48127 124 48171 1022 1 FreeSans 2000 0 0 0 C[57]
port 10 nsew
flabel metal2 s 46239 124 46283 1022 1 FreeSans 2000 0 0 0 C[56]
port 11 nsew
flabel metal2 s 44351 124 44395 1022 1 FreeSans 2000 0 0 0 C[55]
port 12 nsew
flabel metal2 s 42463 124 42507 1022 1 FreeSans 2000 0 0 0 C[54]
port 13 nsew
flabel metal2 s 38687 124 38731 1022 1 FreeSans 2000 0 0 0 C[52]
port 14 nsew
flabel metal2 s 36799 124 36843 1022 1 FreeSans 2000 0 0 0 C[51]
port 15 nsew
flabel metal2 s 34911 124 34955 1022 1 FreeSans 2000 0 0 0 C[50]
port 16 nsew
flabel metal2 s 33023 124 33067 1022 1 FreeSans 2000 0 0 0 C[49]
port 17 nsew
flabel metal2 s 31135 124 31179 1022 1 FreeSans 2000 0 0 0 C[48]
port 18 nsew
flabel metal2 s 29247 124 29291 1022 1 FreeSans 2000 0 0 0 C[47]
port 19 nsew
flabel metal2 s 25471 124 25515 1022 1 FreeSans 2000 0 0 0 C[45]
port 20 nsew
flabel metal2 s 23583 124 23627 1022 1 FreeSans 2000 0 0 0 C[44]
port 21 nsew
flabel metal2 s 21695 124 21739 1022 1 FreeSans 2000 0 0 0 C[43]
port 22 nsew
flabel metal2 s 19807 124 19851 1022 1 FreeSans 2000 0 0 0 C[42]
port 23 nsew
flabel metal2 s 17919 124 17963 1022 1 FreeSans 2000 0 0 0 C[41]
port 24 nsew
flabel metal2 s 16031 124 16075 1022 1 FreeSans 2000 0 0 0 C[40]
port 25 nsew
flabel metal2 s 14143 124 14187 1022 1 FreeSans 2000 0 0 0 C[39]
port 26 nsew
flabel metal2 s 12255 124 12299 1022 1 FreeSans 2000 0 0 0 C[38]
port 27 nsew
flabel metal2 s 10367 124 10411 1022 1 FreeSans 2000 0 0 0 C[37]
port 28 nsew
flabel metal2 s 8479 124 8523 1022 1 FreeSans 2000 0 0 0 C[36]
port 29 nsew
flabel metal2 s 6591 124 6635 1022 1 FreeSans 2000 0 0 0 C[35]
port 30 nsew
flabel metal2 s 4703 124 4747 1022 1 FreeSans 2000 0 0 0 C[34]
port 31 nsew
flabel metal2 s 2815 124 2859 1022 1 FreeSans 2000 0 0 0 C[33]
port 32 nsew
flabel metal2 s 927 124 971 1022 1 FreeSans 2000 0 0 0 C[32]
port 33 nsew
flabel metal2 s 2297 6878 2341 8034 1 FreeSans 2000 0 0 0 C[31]
port 34 nsew
flabel metal2 s 4185 6878 4229 8034 1 FreeSans 2000 0 0 0 C[30]
port 35 nsew
flabel metal2 s 6073 6878 6117 8034 1 FreeSans 2000 0 0 0 C[29]
port 36 nsew
flabel metal2 s 7961 6878 8005 8034 1 FreeSans 2000 0 0 0 C[28]
port 37 nsew
flabel metal2 s 9849 6878 9893 8034 1 FreeSans 2000 0 0 0 C[27]
port 38 nsew
flabel metal2 s 11737 6878 11781 8034 1 FreeSans 2000 0 0 0 C[26]
port 39 nsew
flabel metal2 s 13625 6878 13669 8034 1 FreeSans 2000 0 0 0 C[25]
port 40 nsew
flabel metal2 s 15513 6878 15557 8034 1 FreeSans 2000 0 0 0 C[24]
port 41 nsew
flabel metal2 s 17401 6878 17445 8034 1 FreeSans 2000 0 0 0 C[23]
port 42 nsew
flabel metal2 s 19289 6878 19333 8034 1 FreeSans 2000 0 0 0 C[22]
port 43 nsew
flabel metal2 s 21177 6878 21221 8034 1 FreeSans 2000 0 0 0 C[21]
port 44 nsew
flabel metal2 s 23065 6878 23109 8034 1 FreeSans 2000 0 0 0 C[20]
port 45 nsew
flabel metal2 s 24953 6878 24997 8034 1 FreeSans 2000 0 0 0 C[19]
port 46 nsew
flabel metal2 s 26841 6878 26885 8034 1 FreeSans 2000 0 0 0 C[18]
port 47 nsew
flabel metal2 s 28729 6878 28773 8034 1 FreeSans 2000 0 0 0 C[17]
port 48 nsew
flabel metal2 s 30617 6878 30661 8034 1 FreeSans 2000 0 0 0 C[16]
port 49 nsew
flabel metal2 s 32505 6878 32549 8034 1 FreeSans 2000 0 0 0 C[15]
port 50 nsew
flabel metal2 s 34393 6878 34437 8034 1 FreeSans 2000 0 0 0 C[14]
port 51 nsew
flabel metal2 s 36281 6878 36325 8034 1 FreeSans 2000 0 0 0 C[13]
port 52 nsew
flabel metal2 s 38169 6878 38213 8034 1 FreeSans 2000 0 0 0 C[12]
port 53 nsew
flabel metal2 s 40057 6878 40101 8034 1 FreeSans 2000 0 0 0 C[11]
port 54 nsew
flabel metal2 s 41945 6878 41989 8034 1 FreeSans 2000 0 0 0 C[10]
port 55 nsew
flabel metal2 s 43833 6878 43877 8034 1 FreeSans 2000 0 0 0 C[9]
port 56 nsew
flabel metal2 s 45721 6878 45765 8034 1 FreeSans 2000 0 0 0 C[8]
port 57 nsew
flabel metal2 s 47609 6878 47653 8034 1 FreeSans 2000 0 0 0 C[7]
port 58 nsew
flabel metal2 s 49497 6878 49541 8034 1 FreeSans 2000 0 0 0 C[6]
port 59 nsew
flabel metal2 s 51385 6878 51429 8034 1 FreeSans 2000 0 0 0 C[5]
port 60 nsew
flabel metal2 s 53273 6878 53317 8034 1 FreeSans 2000 0 0 0 C[4]
port 61 nsew
flabel metal2 s 55161 6878 55205 8034 1 FreeSans 2000 0 0 0 C[3]
port 62 nsew
flabel metal2 s 57049 6878 57093 8034 1 FreeSans 2000 0 0 0 C[2]
port 63 nsew
flabel metal2 s 58937 6878 58981 8034 1 FreeSans 2000 0 0 0 C[1]
port 64 nsew
flabel metal2 s 60825 6878 60869 8034 1 FreeSans 2000 0 0 0 C[0]
port 65 nsew
flabel metal2 s 27359 24 27403 922 1 FreeSans 2000 0 0 0 C[46]
port 66 nsew
flabel metal2 s 40575 0 40619 898 1 FreeSans 2000 0 0 0 C[53]
port 67 nsew
flabel metal2 s 57569 4 57613 902 1 FreeSans 2000 0 0 0 C[62]
port 68 nsew
<< end >>
