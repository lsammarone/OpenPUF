magic
tech sky130A
timestamp 1654736712
<< metal3 >>
rect -500 16 500 24
rect -500 -16 -496 16
rect -464 -16 -456 16
rect -424 -16 -416 16
rect -384 -16 -376 16
rect -344 -16 -336 16
rect -304 -16 -296 16
rect -264 -16 -256 16
rect -224 -16 -216 16
rect -184 -16 -176 16
rect -144 -16 -136 16
rect -104 -16 -96 16
rect -64 -16 -56 16
rect -24 -16 -16 16
rect 16 -16 24 16
rect 56 -16 64 16
rect 96 -16 104 16
rect 136 -16 144 16
rect 176 -16 184 16
rect 216 -16 224 16
rect 256 -16 264 16
rect 296 -16 304 16
rect 336 -16 344 16
rect 376 -16 384 16
rect 416 -16 424 16
rect 456 -16 464 16
rect 496 -16 500 16
rect -500 -24 500 -16
<< via3 >>
rect -496 -16 -464 16
rect -456 -16 -424 16
rect -416 -16 -384 16
rect -376 -16 -344 16
rect -336 -16 -304 16
rect -296 -16 -264 16
rect -256 -16 -224 16
rect -216 -16 -184 16
rect -176 -16 -144 16
rect -136 -16 -104 16
rect -96 -16 -64 16
rect -56 -16 -24 16
rect -16 -16 16 16
rect 24 -16 56 16
rect 64 -16 96 16
rect 104 -16 136 16
rect 144 -16 176 16
rect 184 -16 216 16
rect 224 -16 256 16
rect 264 -16 296 16
rect 304 -16 336 16
rect 344 -16 376 16
rect 384 -16 416 16
rect 424 -16 456 16
rect 464 -16 496 16
<< metal4 >>
rect -500 16 500 24
rect -500 -16 -496 16
rect -464 -16 -456 16
rect -424 -16 -416 16
rect -384 -16 -376 16
rect -344 -16 -336 16
rect -304 -16 -296 16
rect -264 -16 -256 16
rect -224 -16 -216 16
rect -184 -16 -176 16
rect -144 -16 -136 16
rect -104 -16 -96 16
rect -64 -16 -56 16
rect -24 -16 -16 16
rect 16 -16 24 16
rect 56 -16 64 16
rect 96 -16 104 16
rect 136 -16 144 16
rect 176 -16 184 16
rect 216 -16 224 16
rect 256 -16 264 16
rect 296 -16 304 16
rect 336 -16 344 16
rect 376 -16 384 16
rect 416 -16 424 16
rect 456 -16 464 16
rect 496 -16 500 16
rect -500 -24 500 -16
<< end >>
