magic
tech sky130A
timestamp 1654736712
<< metal4 >>
rect -500 139 500 155
rect -500 -139 -459 139
rect 459 -139 500 139
rect -500 -155 500 -139
<< via4 >>
rect -459 -139 459 139
<< metal5 >>
rect -500 139 500 155
rect -500 -139 -459 139
rect 459 -139 500 139
rect -500 -155 500 -139
<< end >>
