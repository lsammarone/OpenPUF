magic
tech sky130A
magscale 1 2
timestamp 1656729169
<< nwell >>
rect -38 261 130 582
<< pwell >>
rect 3 38 89 195
<< psubdiff >>
rect 29 145 63 169
rect 29 64 63 111
<< nsubdiff >>
rect 29 456 63 480
rect 29 363 63 422
rect 29 305 63 329
<< psubdiffcont >>
rect 29 111 63 145
<< nsubdiffcont >>
rect 29 422 63 456
rect 29 329 63 363
<< locali >>
rect 0 527 29 561
rect 63 527 92 561
rect 17 456 75 527
rect 17 422 29 456
rect 63 422 75 456
rect 17 363 75 422
rect 17 329 29 363
rect 63 329 75 363
rect 17 294 75 329
rect 17 145 75 162
rect 17 111 29 145
rect 63 111 75 145
rect 17 17 75 111
rect 0 -17 29 17
rect 63 -17 92 17
<< viali >>
rect 29 527 63 561
rect 29 -17 63 17
<< metal1 >>
rect 0 561 92 592
rect 0 527 29 561
rect 63 527 92 561
rect 0 496 92 527
rect 0 17 92 48
rect 0 -17 29 17
rect 63 -17 92 17
rect 0 -48 92 -17
<< labels >>
flabel metal1 s 22 524 75 553 0 FreeSans 200 0 0 0 VPWR
port 1 nsew
flabel metal1 s 21 -18 72 20 0 FreeSans 200 0 0 0 VGND
port 2 nsew
rlabel comment s 0 0 0 0 4 tapvpwrvgnd_1
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 1 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
port 2 nsew
rlabel comment s 0 0 0 0 4 tapvpwrvgnd_1
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 1 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
port 2 nsew
rlabel comment s 0 0 0 0 4 tapvpwrvgnd_1
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 1 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
port 2 nsew
rlabel comment s 0 0 0 0 4 tapvpwrvgnd_1
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 1 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
port 2 nsew
rlabel comment s 0 0 0 0 4 tapvpwrvgnd_1
<< properties >>
string FIXED_BBOX 0 0 92 544
string GDS_END 9277134
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/merge/design_merged.gds
string GDS_START 9269050
<< end >>
