magic
tech sky130A
magscale 1 2
timestamp 1656729169
<< error_p >>
rect -38 261 314 582
rect 29 47 81 177
rect 111 47 165 177
rect 195 47 247 177
<< nwell >>
rect -38 261 314 582
<< pwell >>
rect 3 21 273 203
rect 29 -17 63 21
<< scnmos >>
rect 81 47 111 177
rect 165 47 195 177
<< scpmoshvt >>
rect 81 297 111 497
rect 165 297 195 497
<< ndiff >>
rect 29 165 81 177
rect 29 131 37 165
rect 71 131 81 165
rect 29 93 81 131
rect 29 59 37 93
rect 71 59 81 93
rect 29 47 81 59
rect 111 165 165 177
rect 111 131 121 165
rect 155 131 165 165
rect 111 93 165 131
rect 111 59 121 93
rect 155 59 165 93
rect 111 47 165 59
rect 195 165 247 177
rect 195 131 205 165
rect 239 131 247 165
rect 195 93 247 131
rect 195 59 205 93
rect 239 59 247 93
rect 195 47 247 59
<< pdiff >>
rect 29 485 81 497
rect 29 451 37 485
rect 71 451 81 485
rect 29 417 81 451
rect 29 383 37 417
rect 71 383 81 417
rect 29 349 81 383
rect 29 315 37 349
rect 71 315 81 349
rect 29 297 81 315
rect 111 485 165 497
rect 111 451 121 485
rect 155 451 165 485
rect 111 417 165 451
rect 111 383 121 417
rect 155 383 165 417
rect 111 349 165 383
rect 111 315 121 349
rect 155 315 165 349
rect 111 297 165 315
rect 195 485 247 497
rect 195 451 205 485
rect 239 451 247 485
rect 195 417 247 451
rect 195 383 205 417
rect 239 383 247 417
rect 195 349 247 383
rect 195 315 205 349
rect 239 315 247 349
rect 195 297 247 315
<< ndiffc >>
rect 37 131 71 165
rect 37 59 71 93
rect 121 131 155 165
rect 121 59 155 93
rect 205 131 239 165
rect 205 59 239 93
<< pdiffc >>
rect 37 451 71 485
rect 37 383 71 417
rect 37 315 71 349
rect 121 451 155 485
rect 121 383 155 417
rect 121 315 155 349
rect 205 451 239 485
rect 205 383 239 417
rect 205 315 239 349
<< poly >>
rect 81 497 111 523
rect 165 497 195 523
rect 81 265 111 297
rect 165 265 195 297
rect 21 249 195 265
rect 21 215 37 249
rect 71 215 195 249
rect 21 199 195 215
rect 81 177 111 199
rect 165 177 195 199
rect 81 21 111 47
rect 165 21 195 47
<< polycont >>
rect 37 215 71 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 25 485 71 527
rect 25 451 37 485
rect 25 417 71 451
rect 25 383 37 417
rect 25 349 71 383
rect 25 315 37 349
rect 25 299 71 315
rect 105 485 171 493
rect 105 451 121 485
rect 155 451 171 485
rect 105 417 171 451
rect 105 383 121 417
rect 155 383 171 417
rect 105 349 171 383
rect 105 315 121 349
rect 155 315 171 349
rect 105 297 171 315
rect 205 485 247 527
rect 239 451 247 485
rect 205 417 247 451
rect 239 383 247 417
rect 205 349 247 383
rect 239 315 247 349
rect 205 299 247 315
rect 21 249 87 265
rect 21 215 37 249
rect 71 215 87 249
rect 25 165 71 181
rect 121 177 171 297
rect 25 131 37 165
rect 25 93 71 131
rect 25 59 37 93
rect 25 17 71 59
rect 105 165 171 177
rect 105 131 121 165
rect 155 131 171 165
rect 105 93 171 131
rect 105 59 121 93
rect 155 59 171 93
rect 105 51 171 59
rect 205 165 247 181
rect 239 131 247 165
rect 205 93 247 131
rect 239 59 247 93
rect 205 17 247 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
<< metal1 >>
rect 0 561 276 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 496 276 527
rect 0 17 276 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 0 -48 276 -17
<< labels >>
flabel locali s 29 221 63 255 0 FreeSans 531 0 0 0 A
port 1 nsew
flabel locali s 121 153 155 187 0 FreeSans 531 0 0 0 Y
port 2 nsew
flabel locali s 121 289 155 323 0 FreeSans 531 0 0 0 Y
port 2 nsew
flabel locali s 121 221 155 255 0 FreeSans 531 0 0 0 Y
port 2 nsew
flabel nwell s 29 527 63 561 0 FreeSans 312 0 0 0 VPB
port 3 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 312 0 0 0 VNB
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 312 0 0 0 VPWR
port 5 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 312 0 0 0 VGND
port 6 nsew
flabel locali s 46 238 46 238 0 FreeSans 531 0 0 0 A
port 1 nsew
flabel locali s 138 170 138 170 0 FreeSans 531 0 0 0 Y
port 2 nsew
flabel locali s 138 306 138 306 0 FreeSans 531 0 0 0 Y
port 2 nsew
flabel locali s 138 238 138 238 0 FreeSans 531 0 0 0 Y
port 2 nsew
flabel nwell s 46 544 46 544 0 FreeSans 312 0 0 0 VPB
port 3 nsew
flabel pwell s 46 0 46 0 0 FreeSans 312 0 0 0 VNB
port 4 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 312 0 0 0 VPWR
port 5 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 312 0 0 0 VGND
port 6 nsew
flabel locali s 46 238 46 238 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel locali s 138 170 138 170 0 FreeSans 340 0 0 0 Y
port 2 nsew
flabel locali s 138 306 138 306 0 FreeSans 340 0 0 0 Y
port 2 nsew
flabel locali s 138 238 138 238 0 FreeSans 340 0 0 0 Y
port 2 nsew
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 3 nsew
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
port 6 nsew
rlabel comment s 0 0 0 0 4 inv_2
<< properties >>
string FIXED_BBOX 0 0 276 544
string GDS_END 9932344
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/merge/design_merged.gds
string GDS_START 9920420
string path 0.000 0.000 6.900 0.000 
<< end >>
