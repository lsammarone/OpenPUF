magic
tech sky130A
timestamp 1655322987
<< metal2 >>
rect -90 34 90 45
rect -90 -34 -74 34
rect 74 -34 90 34
rect -90 -45 90 -34
<< via2 >>
rect -74 -34 74 34
<< metal3 >>
rect -90 34 90 45
rect -90 -34 -74 34
rect 74 -34 90 34
rect -90 -45 90 -34
<< end >>
