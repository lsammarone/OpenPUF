magic
tech sky130A
magscale 1 2
timestamp 1656729169
<< error_p >>
rect -33 32 33 33
rect -38 -32 -32 32
rect -33 -33 33 -32
<< metal3 >>
rect -38 -32 -32 32
rect 32 -32 38 32
<< via3 >>
rect -32 -32 32 32
<< metal4 >>
rect -33 32 33 33
rect -33 -32 -32 32
rect 32 -32 33 32
rect -33 -33 33 -32
<< end >>
