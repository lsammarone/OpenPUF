magic
tech sky130A
magscale 1 2
timestamp 1655322987
<< metal4 >>
rect -180 918 180 969
rect -180 682 -118 918
rect 118 682 180 918
rect -180 598 180 682
rect -180 362 -118 598
rect 118 362 180 598
rect -180 278 180 362
rect -180 42 -118 278
rect 118 42 180 278
rect -180 -42 180 42
rect -180 -278 -118 -42
rect 118 -278 180 -42
rect -180 -362 180 -278
rect -180 -598 -118 -362
rect 118 -598 180 -362
rect -180 -682 180 -598
rect -180 -918 -118 -682
rect 118 -918 180 -682
rect -180 -969 180 -918
<< via4 >>
rect -118 682 118 918
rect -118 362 118 598
rect -118 42 118 278
rect -118 -278 118 -42
rect -118 -598 118 -362
rect -118 -918 118 -682
<< metal5 >>
rect -180 918 180 969
rect -180 682 -118 918
rect 118 682 180 918
rect -180 598 180 682
rect -180 362 -118 598
rect 118 362 180 598
rect -180 278 180 362
rect -180 42 -118 278
rect 118 42 180 278
rect -180 -42 180 42
rect -180 -278 -118 -42
rect 118 -278 180 -42
rect -180 -362 180 -278
rect -180 -598 -118 -362
rect 118 -598 180 -362
rect -180 -682 180 -598
rect -180 -918 -118 -682
rect 118 -918 180 -682
rect -180 -969 180 -918
<< end >>
