magic
tech sky130A
magscale 1 2
timestamp 1656729169
<< locali >>
rect 122 1897 7290 1910
rect 122 1863 305 1897
rect 339 1863 705 1897
rect 739 1863 1105 1897
rect 1139 1863 1505 1897
rect 1539 1863 1905 1897
rect 1939 1863 2305 1897
rect 2339 1863 2705 1897
rect 2739 1863 3105 1897
rect 3139 1863 3505 1897
rect 3539 1863 3905 1897
rect 3939 1863 4305 1897
rect 4339 1863 4705 1897
rect 4739 1863 5105 1897
rect 5139 1863 5505 1897
rect 5539 1863 5905 1897
rect 5939 1863 6305 1897
rect 6339 1863 6705 1897
rect 6739 1863 7105 1897
rect 7139 1863 7290 1897
rect 122 1850 7290 1863
rect 122 17 7290 30
rect 122 -17 305 17
rect 339 -17 705 17
rect 739 -17 1105 17
rect 1139 -17 1505 17
rect 1539 -17 1905 17
rect 1939 -17 2305 17
rect 2339 -17 2705 17
rect 2739 -17 3105 17
rect 3139 -17 3505 17
rect 3539 -17 3905 17
rect 3939 -17 4305 17
rect 4339 -17 4705 17
rect 4739 -17 5105 17
rect 5139 -17 5505 17
rect 5539 -17 5905 17
rect 5939 -17 6305 17
rect 6339 -17 6705 17
rect 6739 -17 7105 17
rect 7139 -17 7290 17
rect 122 -30 7290 -17
<< viali >>
rect 305 1863 339 1897
rect 705 1863 739 1897
rect 1105 1863 1139 1897
rect 1505 1863 1539 1897
rect 1905 1863 1939 1897
rect 2305 1863 2339 1897
rect 2705 1863 2739 1897
rect 3105 1863 3139 1897
rect 3505 1863 3539 1897
rect 3905 1863 3939 1897
rect 4305 1863 4339 1897
rect 4705 1863 4739 1897
rect 5105 1863 5139 1897
rect 5505 1863 5539 1897
rect 5905 1863 5939 1897
rect 6305 1863 6339 1897
rect 6705 1863 6739 1897
rect 7105 1863 7139 1897
rect 305 -17 339 17
rect 705 -17 739 17
rect 1105 -17 1139 17
rect 1505 -17 1539 17
rect 1905 -17 1939 17
rect 2305 -17 2339 17
rect 2705 -17 2739 17
rect 3105 -17 3139 17
rect 3505 -17 3539 17
rect 3905 -17 3939 17
rect 4305 -17 4339 17
rect 4705 -17 4739 17
rect 5105 -17 5139 17
rect 5505 -17 5539 17
rect 5905 -17 5939 17
rect 6305 -17 6339 17
rect 6705 -17 6739 17
rect 7105 -17 7139 17
<< metal1 >>
rect 122 1897 7290 1940
rect 122 1863 305 1897
rect 339 1863 705 1897
rect 739 1863 1105 1897
rect 1139 1863 1505 1897
rect 1539 1863 1905 1897
rect 1939 1863 2305 1897
rect 2339 1863 2705 1897
rect 2739 1863 3105 1897
rect 3139 1863 3505 1897
rect 3539 1863 3905 1897
rect 3939 1863 4305 1897
rect 4339 1863 4705 1897
rect 4739 1863 5105 1897
rect 5139 1863 5505 1897
rect 5539 1863 5905 1897
rect 5939 1863 6305 1897
rect 6339 1863 6705 1897
rect 6739 1863 7105 1897
rect 7139 1863 7290 1897
rect 122 1820 7290 1863
rect 122 17 7290 60
rect 122 -17 305 17
rect 339 -17 705 17
rect 739 -17 1105 17
rect 1139 -17 1505 17
rect 1539 -17 1905 17
rect 1939 -17 2305 17
rect 2339 -17 2705 17
rect 2739 -17 3105 17
rect 3139 -17 3505 17
rect 3539 -17 3905 17
rect 3939 -17 4305 17
rect 4339 -17 4705 17
rect 4739 -17 5105 17
rect 5139 -17 5505 17
rect 5539 -17 5905 17
rect 5939 -17 6305 17
rect 6339 -17 6705 17
rect 6739 -17 7105 17
rect 7139 -17 7290 17
rect 122 -60 7290 -17
<< metal2 >>
rect 120 1638 320 1650
rect 120 1582 152 1638
rect 208 1582 232 1638
rect 288 1582 320 1638
rect 120 1570 320 1582
rect 142 218 302 240
rect 142 162 194 218
rect 250 162 302 218
rect 142 140 302 162
<< via2 >>
rect 152 1582 208 1638
rect 232 1582 288 1638
rect 194 162 250 218
<< metal3 >>
rect 120 1638 7292 1650
rect 120 1582 152 1638
rect 208 1582 232 1638
rect 288 1622 7292 1638
rect 288 1582 736 1622
rect 120 1558 736 1582
rect 800 1558 1455 1622
rect 1519 1558 2174 1622
rect 2238 1558 2893 1622
rect 2957 1558 3612 1622
rect 3676 1558 4331 1622
rect 4395 1558 5050 1622
rect 5114 1558 5769 1622
rect 5833 1558 6488 1622
rect 6552 1558 7207 1622
rect 7271 1558 7292 1622
rect 120 1542 7292 1558
rect 120 1478 736 1542
rect 800 1478 1455 1542
rect 1519 1478 2174 1542
rect 2238 1478 2893 1542
rect 2957 1478 3612 1542
rect 3676 1478 4331 1542
rect 4395 1478 5050 1542
rect 5114 1478 5769 1542
rect 5833 1478 6488 1542
rect 6552 1478 7207 1542
rect 7271 1478 7292 1542
rect 120 1462 7292 1478
rect 120 1398 736 1462
rect 800 1398 1455 1462
rect 1519 1398 2174 1462
rect 2238 1398 2893 1462
rect 2957 1398 3612 1462
rect 3676 1398 4331 1462
rect 4395 1398 5050 1462
rect 5114 1398 5769 1462
rect 5833 1398 6488 1462
rect 6552 1398 7207 1462
rect 7271 1398 7292 1462
rect 120 1382 7292 1398
rect 120 1318 736 1382
rect 800 1318 1455 1382
rect 1519 1318 2174 1382
rect 2238 1318 2893 1382
rect 2957 1318 3612 1382
rect 3676 1318 4331 1382
rect 4395 1318 5050 1382
rect 5114 1318 5769 1382
rect 5833 1318 6488 1382
rect 6552 1318 7207 1382
rect 7271 1318 7292 1382
rect 120 1302 7292 1318
rect 120 1238 736 1302
rect 800 1238 1455 1302
rect 1519 1238 2174 1302
rect 2238 1238 2893 1302
rect 2957 1238 3612 1302
rect 3676 1238 4331 1302
rect 4395 1238 5050 1302
rect 5114 1238 5769 1302
rect 5833 1238 6488 1302
rect 6552 1238 7207 1302
rect 7271 1238 7292 1302
rect 120 1222 7292 1238
rect 120 1158 736 1222
rect 800 1158 1455 1222
rect 1519 1158 2174 1222
rect 2238 1158 2893 1222
rect 2957 1158 3612 1222
rect 3676 1158 4331 1222
rect 4395 1158 5050 1222
rect 5114 1158 5769 1222
rect 5833 1158 6488 1222
rect 6552 1158 7207 1222
rect 7271 1158 7292 1222
rect 120 1142 7292 1158
rect 120 1078 736 1142
rect 800 1078 1455 1142
rect 1519 1078 2174 1142
rect 2238 1078 2893 1142
rect 2957 1078 3612 1142
rect 3676 1078 4331 1142
rect 4395 1078 5050 1142
rect 5114 1078 5769 1142
rect 5833 1078 6488 1142
rect 6552 1078 7207 1142
rect 7271 1078 7292 1142
rect 120 922 7292 1078
rect 120 858 736 922
rect 800 858 1455 922
rect 1519 858 2174 922
rect 2238 858 2893 922
rect 2957 858 3612 922
rect 3676 858 4331 922
rect 4395 858 5050 922
rect 5114 858 5769 922
rect 5833 858 6488 922
rect 6552 858 7207 922
rect 7271 858 7292 922
rect 120 842 7292 858
rect 120 778 736 842
rect 800 778 1455 842
rect 1519 778 2174 842
rect 2238 778 2893 842
rect 2957 778 3612 842
rect 3676 778 4331 842
rect 4395 778 5050 842
rect 5114 778 5769 842
rect 5833 778 6488 842
rect 6552 778 7207 842
rect 7271 778 7292 842
rect 120 762 7292 778
rect 120 698 736 762
rect 800 698 1455 762
rect 1519 698 2174 762
rect 2238 698 2893 762
rect 2957 698 3612 762
rect 3676 698 4331 762
rect 4395 698 5050 762
rect 5114 698 5769 762
rect 5833 698 6488 762
rect 6552 698 7207 762
rect 7271 698 7292 762
rect 120 682 7292 698
rect 120 618 736 682
rect 800 618 1455 682
rect 1519 618 2174 682
rect 2238 618 2893 682
rect 2957 618 3612 682
rect 3676 618 4331 682
rect 4395 618 5050 682
rect 5114 618 5769 682
rect 5833 618 6488 682
rect 6552 618 7207 682
rect 7271 618 7292 682
rect 120 602 7292 618
rect 120 538 736 602
rect 800 538 1455 602
rect 1519 538 2174 602
rect 2238 538 2893 602
rect 2957 538 3612 602
rect 3676 538 4331 602
rect 4395 538 5050 602
rect 5114 538 5769 602
rect 5833 538 6488 602
rect 6552 538 7207 602
rect 7271 538 7292 602
rect 120 522 7292 538
rect 120 458 736 522
rect 800 458 1455 522
rect 1519 458 2174 522
rect 2238 458 2893 522
rect 2957 458 3612 522
rect 3676 458 4331 522
rect 4395 458 5050 522
rect 5114 458 5769 522
rect 5833 458 6488 522
rect 6552 458 7207 522
rect 7271 458 7292 522
rect 120 442 7292 458
rect 120 378 736 442
rect 800 378 1455 442
rect 1519 378 2174 442
rect 2238 378 2893 442
rect 2957 378 3612 442
rect 3676 378 4331 442
rect 4395 378 5050 442
rect 5114 378 5769 442
rect 5833 378 6488 442
rect 6552 378 7207 442
rect 7271 378 7292 442
rect 120 350 7292 378
rect 122 222 322 250
rect 122 158 150 222
rect 214 218 230 222
rect 214 158 230 162
rect 294 158 322 222
rect 122 130 322 158
<< via3 >>
rect 736 1558 800 1622
rect 1455 1558 1519 1622
rect 2174 1558 2238 1622
rect 2893 1558 2957 1622
rect 3612 1558 3676 1622
rect 4331 1558 4395 1622
rect 5050 1558 5114 1622
rect 5769 1558 5833 1622
rect 6488 1558 6552 1622
rect 7207 1558 7271 1622
rect 736 1478 800 1542
rect 1455 1478 1519 1542
rect 2174 1478 2238 1542
rect 2893 1478 2957 1542
rect 3612 1478 3676 1542
rect 4331 1478 4395 1542
rect 5050 1478 5114 1542
rect 5769 1478 5833 1542
rect 6488 1478 6552 1542
rect 7207 1478 7271 1542
rect 736 1398 800 1462
rect 1455 1398 1519 1462
rect 2174 1398 2238 1462
rect 2893 1398 2957 1462
rect 3612 1398 3676 1462
rect 4331 1398 4395 1462
rect 5050 1398 5114 1462
rect 5769 1398 5833 1462
rect 6488 1398 6552 1462
rect 7207 1398 7271 1462
rect 736 1318 800 1382
rect 1455 1318 1519 1382
rect 2174 1318 2238 1382
rect 2893 1318 2957 1382
rect 3612 1318 3676 1382
rect 4331 1318 4395 1382
rect 5050 1318 5114 1382
rect 5769 1318 5833 1382
rect 6488 1318 6552 1382
rect 7207 1318 7271 1382
rect 736 1238 800 1302
rect 1455 1238 1519 1302
rect 2174 1238 2238 1302
rect 2893 1238 2957 1302
rect 3612 1238 3676 1302
rect 4331 1238 4395 1302
rect 5050 1238 5114 1302
rect 5769 1238 5833 1302
rect 6488 1238 6552 1302
rect 7207 1238 7271 1302
rect 736 1158 800 1222
rect 1455 1158 1519 1222
rect 2174 1158 2238 1222
rect 2893 1158 2957 1222
rect 3612 1158 3676 1222
rect 4331 1158 4395 1222
rect 5050 1158 5114 1222
rect 5769 1158 5833 1222
rect 6488 1158 6552 1222
rect 7207 1158 7271 1222
rect 736 1078 800 1142
rect 1455 1078 1519 1142
rect 2174 1078 2238 1142
rect 2893 1078 2957 1142
rect 3612 1078 3676 1142
rect 4331 1078 4395 1142
rect 5050 1078 5114 1142
rect 5769 1078 5833 1142
rect 6488 1078 6552 1142
rect 7207 1078 7271 1142
rect 736 858 800 922
rect 1455 858 1519 922
rect 2174 858 2238 922
rect 2893 858 2957 922
rect 3612 858 3676 922
rect 4331 858 4395 922
rect 5050 858 5114 922
rect 5769 858 5833 922
rect 6488 858 6552 922
rect 7207 858 7271 922
rect 736 778 800 842
rect 1455 778 1519 842
rect 2174 778 2238 842
rect 2893 778 2957 842
rect 3612 778 3676 842
rect 4331 778 4395 842
rect 5050 778 5114 842
rect 5769 778 5833 842
rect 6488 778 6552 842
rect 7207 778 7271 842
rect 736 698 800 762
rect 1455 698 1519 762
rect 2174 698 2238 762
rect 2893 698 2957 762
rect 3612 698 3676 762
rect 4331 698 4395 762
rect 5050 698 5114 762
rect 5769 698 5833 762
rect 6488 698 6552 762
rect 7207 698 7271 762
rect 736 618 800 682
rect 1455 618 1519 682
rect 2174 618 2238 682
rect 2893 618 2957 682
rect 3612 618 3676 682
rect 4331 618 4395 682
rect 5050 618 5114 682
rect 5769 618 5833 682
rect 6488 618 6552 682
rect 7207 618 7271 682
rect 736 538 800 602
rect 1455 538 1519 602
rect 2174 538 2238 602
rect 2893 538 2957 602
rect 3612 538 3676 602
rect 4331 538 4395 602
rect 5050 538 5114 602
rect 5769 538 5833 602
rect 6488 538 6552 602
rect 7207 538 7271 602
rect 736 458 800 522
rect 1455 458 1519 522
rect 2174 458 2238 522
rect 2893 458 2957 522
rect 3612 458 3676 522
rect 4331 458 4395 522
rect 5050 458 5114 522
rect 5769 458 5833 522
rect 6488 458 6552 522
rect 7207 458 7271 522
rect 736 378 800 442
rect 1455 378 1519 442
rect 2174 378 2238 442
rect 2893 378 2957 442
rect 3612 378 3676 442
rect 4331 378 4395 442
rect 5050 378 5114 442
rect 5769 378 5833 442
rect 6488 378 6552 442
rect 7207 378 7271 442
rect 150 218 214 222
rect 230 218 294 222
rect 150 162 194 218
rect 194 162 214 218
rect 230 162 250 218
rect 250 162 294 218
rect 150 158 214 162
rect 230 158 294 162
<< mimcap >>
rect 221 1502 621 1550
rect 221 1198 269 1502
rect 573 1198 621 1502
rect 221 1150 621 1198
rect 940 1502 1340 1550
rect 940 1198 988 1502
rect 1292 1198 1340 1502
rect 940 1150 1340 1198
rect 1659 1502 2059 1550
rect 1659 1198 1707 1502
rect 2011 1198 2059 1502
rect 1659 1150 2059 1198
rect 2378 1502 2778 1550
rect 2378 1198 2426 1502
rect 2730 1198 2778 1502
rect 2378 1150 2778 1198
rect 3097 1502 3497 1550
rect 3097 1198 3145 1502
rect 3449 1198 3497 1502
rect 3097 1150 3497 1198
rect 3816 1502 4216 1550
rect 3816 1198 3864 1502
rect 4168 1198 4216 1502
rect 3816 1150 4216 1198
rect 4535 1502 4935 1550
rect 4535 1198 4583 1502
rect 4887 1198 4935 1502
rect 4535 1150 4935 1198
rect 5254 1502 5654 1550
rect 5254 1198 5302 1502
rect 5606 1198 5654 1502
rect 5254 1150 5654 1198
rect 5973 1502 6373 1550
rect 5973 1198 6021 1502
rect 6325 1198 6373 1502
rect 5973 1150 6373 1198
rect 6692 1502 7092 1550
rect 6692 1198 6740 1502
rect 7044 1198 7092 1502
rect 6692 1150 7092 1198
rect 221 802 621 850
rect 221 498 269 802
rect 573 498 621 802
rect 221 450 621 498
rect 940 802 1340 850
rect 940 498 988 802
rect 1292 498 1340 802
rect 940 450 1340 498
rect 1659 802 2059 850
rect 1659 498 1707 802
rect 2011 498 2059 802
rect 1659 450 2059 498
rect 2378 802 2778 850
rect 2378 498 2426 802
rect 2730 498 2778 802
rect 2378 450 2778 498
rect 3097 802 3497 850
rect 3097 498 3145 802
rect 3449 498 3497 802
rect 3097 450 3497 498
rect 3816 802 4216 850
rect 3816 498 3864 802
rect 4168 498 4216 802
rect 3816 450 4216 498
rect 4535 802 4935 850
rect 4535 498 4583 802
rect 4887 498 4935 802
rect 4535 450 4935 498
rect 5254 802 5654 850
rect 5254 498 5302 802
rect 5606 498 5654 802
rect 5254 450 5654 498
rect 5973 802 6373 850
rect 5973 498 6021 802
rect 6325 498 6373 802
rect 5973 450 6373 498
rect 6692 802 7092 850
rect 6692 498 6740 802
rect 7044 498 7092 802
rect 6692 450 7092 498
<< mimcapcontact >>
rect 269 1198 573 1502
rect 988 1198 1292 1502
rect 1707 1198 2011 1502
rect 2426 1198 2730 1502
rect 3145 1198 3449 1502
rect 3864 1198 4168 1502
rect 4583 1198 4887 1502
rect 5302 1198 5606 1502
rect 6021 1198 6325 1502
rect 6740 1198 7044 1502
rect 269 498 573 802
rect 988 498 1292 802
rect 1707 498 2011 802
rect 2426 498 2730 802
rect 3145 498 3449 802
rect 3864 498 4168 802
rect 4583 498 4887 802
rect 5302 498 5606 802
rect 6021 498 6325 802
rect 6740 498 7044 802
<< metal4 >>
rect 720 1622 816 1638
rect 720 1558 736 1622
rect 800 1558 816 1622
rect 720 1542 816 1558
rect 260 1511 580 1530
rect 260 1502 582 1511
rect 260 1198 269 1502
rect 573 1198 582 1502
rect 260 1189 582 1198
rect 720 1478 736 1542
rect 800 1478 816 1542
rect 1439 1622 1535 1638
rect 1439 1558 1455 1622
rect 1519 1558 1535 1622
rect 1439 1542 1535 1558
rect 980 1511 1300 1530
rect 720 1462 816 1478
rect 720 1398 736 1462
rect 800 1398 816 1462
rect 720 1382 816 1398
rect 720 1318 736 1382
rect 800 1318 816 1382
rect 720 1302 816 1318
rect 720 1238 736 1302
rect 800 1238 816 1302
rect 720 1222 816 1238
rect 260 811 580 1189
rect 720 1158 736 1222
rect 800 1158 816 1222
rect 979 1502 1301 1511
rect 979 1198 988 1502
rect 1292 1198 1301 1502
rect 979 1189 1301 1198
rect 1439 1478 1455 1542
rect 1519 1478 1535 1542
rect 2158 1622 2254 1638
rect 2158 1558 2174 1622
rect 2238 1558 2254 1622
rect 2158 1542 2254 1558
rect 1700 1511 2020 1530
rect 1439 1462 1535 1478
rect 1439 1398 1455 1462
rect 1519 1398 1535 1462
rect 1439 1382 1535 1398
rect 1439 1318 1455 1382
rect 1519 1318 1535 1382
rect 1439 1302 1535 1318
rect 1439 1238 1455 1302
rect 1519 1238 1535 1302
rect 1439 1222 1535 1238
rect 720 1142 816 1158
rect 720 1078 736 1142
rect 800 1078 816 1142
rect 720 1062 816 1078
rect 720 922 816 938
rect 720 858 736 922
rect 800 858 816 922
rect 720 842 816 858
rect 260 802 582 811
rect 260 498 269 802
rect 573 498 582 802
rect 260 489 582 498
rect 720 778 736 842
rect 800 778 816 842
rect 980 811 1300 1189
rect 1439 1158 1455 1222
rect 1519 1158 1535 1222
rect 1698 1502 2020 1511
rect 1698 1198 1707 1502
rect 2011 1198 2020 1502
rect 1698 1189 2020 1198
rect 1439 1142 1535 1158
rect 1439 1078 1455 1142
rect 1519 1078 1535 1142
rect 1439 1062 1535 1078
rect 1439 922 1535 938
rect 1439 858 1455 922
rect 1519 858 1535 922
rect 1439 842 1535 858
rect 720 762 816 778
rect 720 698 736 762
rect 800 698 816 762
rect 720 682 816 698
rect 720 618 736 682
rect 800 618 816 682
rect 720 602 816 618
rect 720 538 736 602
rect 800 538 816 602
rect 720 522 816 538
rect 260 250 580 489
rect 720 458 736 522
rect 800 458 816 522
rect 979 802 1301 811
rect 979 498 988 802
rect 1292 498 1301 802
rect 979 489 1301 498
rect 1439 778 1455 842
rect 1519 778 1535 842
rect 1700 811 2020 1189
rect 2158 1478 2174 1542
rect 2238 1478 2254 1542
rect 2877 1622 2973 1638
rect 2877 1558 2893 1622
rect 2957 1558 2973 1622
rect 2877 1542 2973 1558
rect 2420 1511 2740 1530
rect 2158 1462 2254 1478
rect 2158 1398 2174 1462
rect 2238 1398 2254 1462
rect 2158 1382 2254 1398
rect 2158 1318 2174 1382
rect 2238 1318 2254 1382
rect 2158 1302 2254 1318
rect 2158 1238 2174 1302
rect 2238 1238 2254 1302
rect 2158 1222 2254 1238
rect 2158 1158 2174 1222
rect 2238 1158 2254 1222
rect 2417 1502 2740 1511
rect 2417 1198 2426 1502
rect 2730 1198 2740 1502
rect 2417 1189 2740 1198
rect 2158 1142 2254 1158
rect 2158 1078 2174 1142
rect 2238 1078 2254 1142
rect 2158 1062 2254 1078
rect 1439 762 1535 778
rect 1439 698 1455 762
rect 1519 698 1535 762
rect 1439 682 1535 698
rect 1439 618 1455 682
rect 1519 618 1535 682
rect 1439 602 1535 618
rect 1439 538 1455 602
rect 1519 538 1535 602
rect 1439 522 1535 538
rect 720 442 816 458
rect 720 378 736 442
rect 800 378 816 442
rect 720 362 816 378
rect 980 250 1300 489
rect 1439 458 1455 522
rect 1519 458 1535 522
rect 1698 802 2020 811
rect 1698 498 1707 802
rect 2011 498 2020 802
rect 1698 489 2020 498
rect 1439 442 1535 458
rect 1439 378 1455 442
rect 1519 378 1535 442
rect 1439 362 1535 378
rect 1700 250 2020 489
rect 2158 922 2254 938
rect 2158 858 2174 922
rect 2238 858 2254 922
rect 2158 842 2254 858
rect 2158 778 2174 842
rect 2238 778 2254 842
rect 2420 811 2740 1189
rect 2877 1478 2893 1542
rect 2957 1478 2973 1542
rect 3596 1622 3692 1638
rect 3596 1558 3612 1622
rect 3676 1558 3692 1622
rect 3596 1542 3692 1558
rect 3140 1511 3460 1530
rect 2877 1462 2973 1478
rect 2877 1398 2893 1462
rect 2957 1398 2973 1462
rect 2877 1382 2973 1398
rect 2877 1318 2893 1382
rect 2957 1318 2973 1382
rect 2877 1302 2973 1318
rect 2877 1238 2893 1302
rect 2957 1238 2973 1302
rect 2877 1222 2973 1238
rect 2877 1158 2893 1222
rect 2957 1158 2973 1222
rect 3136 1502 3460 1511
rect 3136 1198 3145 1502
rect 3449 1198 3460 1502
rect 3136 1189 3460 1198
rect 2877 1142 2973 1158
rect 2877 1078 2893 1142
rect 2957 1078 2973 1142
rect 2877 1062 2973 1078
rect 2158 762 2254 778
rect 2158 698 2174 762
rect 2238 698 2254 762
rect 2158 682 2254 698
rect 2158 618 2174 682
rect 2238 618 2254 682
rect 2158 602 2254 618
rect 2158 538 2174 602
rect 2238 538 2254 602
rect 2158 522 2254 538
rect 2158 458 2174 522
rect 2238 458 2254 522
rect 2417 802 2740 811
rect 2417 498 2426 802
rect 2730 498 2740 802
rect 2417 489 2740 498
rect 2158 442 2254 458
rect 2158 378 2174 442
rect 2238 378 2254 442
rect 2158 362 2254 378
rect 2420 250 2740 489
rect 2877 922 2973 938
rect 2877 858 2893 922
rect 2957 858 2973 922
rect 2877 842 2973 858
rect 2877 778 2893 842
rect 2957 778 2973 842
rect 3140 811 3460 1189
rect 3596 1478 3612 1542
rect 3676 1478 3692 1542
rect 4315 1622 4411 1638
rect 4315 1558 4331 1622
rect 4395 1558 4411 1622
rect 4315 1542 4411 1558
rect 3860 1511 4180 1530
rect 3596 1462 3692 1478
rect 3596 1398 3612 1462
rect 3676 1398 3692 1462
rect 3596 1382 3692 1398
rect 3596 1318 3612 1382
rect 3676 1318 3692 1382
rect 3596 1302 3692 1318
rect 3596 1238 3612 1302
rect 3676 1238 3692 1302
rect 3596 1222 3692 1238
rect 3596 1158 3612 1222
rect 3676 1158 3692 1222
rect 3855 1502 4180 1511
rect 3855 1198 3864 1502
rect 4168 1198 4180 1502
rect 3855 1189 4180 1198
rect 3596 1142 3692 1158
rect 3596 1078 3612 1142
rect 3676 1078 3692 1142
rect 3596 1062 3692 1078
rect 2877 762 2973 778
rect 2877 698 2893 762
rect 2957 698 2973 762
rect 2877 682 2973 698
rect 2877 618 2893 682
rect 2957 618 2973 682
rect 2877 602 2973 618
rect 2877 538 2893 602
rect 2957 538 2973 602
rect 2877 522 2973 538
rect 2877 458 2893 522
rect 2957 458 2973 522
rect 3136 802 3460 811
rect 3136 498 3145 802
rect 3449 498 3460 802
rect 3136 489 3460 498
rect 2877 442 2973 458
rect 2877 378 2893 442
rect 2957 378 2973 442
rect 2877 362 2973 378
rect 3140 250 3460 489
rect 3596 922 3692 938
rect 3596 858 3612 922
rect 3676 858 3692 922
rect 3596 842 3692 858
rect 3596 778 3612 842
rect 3676 778 3692 842
rect 3860 811 4180 1189
rect 4315 1478 4331 1542
rect 4395 1478 4411 1542
rect 5034 1622 5130 1638
rect 5034 1558 5050 1622
rect 5114 1558 5130 1622
rect 5034 1542 5130 1558
rect 4580 1511 4900 1530
rect 4315 1462 4411 1478
rect 4315 1398 4331 1462
rect 4395 1398 4411 1462
rect 4315 1382 4411 1398
rect 4315 1318 4331 1382
rect 4395 1318 4411 1382
rect 4315 1302 4411 1318
rect 4315 1238 4331 1302
rect 4395 1238 4411 1302
rect 4315 1222 4411 1238
rect 4315 1158 4331 1222
rect 4395 1158 4411 1222
rect 4574 1502 4900 1511
rect 4574 1198 4583 1502
rect 4887 1198 4900 1502
rect 4574 1189 4900 1198
rect 4315 1142 4411 1158
rect 4315 1078 4331 1142
rect 4395 1078 4411 1142
rect 4315 1062 4411 1078
rect 3596 762 3692 778
rect 3596 698 3612 762
rect 3676 698 3692 762
rect 3596 682 3692 698
rect 3596 618 3612 682
rect 3676 618 3692 682
rect 3596 602 3692 618
rect 3596 538 3612 602
rect 3676 538 3692 602
rect 3596 522 3692 538
rect 3596 458 3612 522
rect 3676 458 3692 522
rect 3855 802 4180 811
rect 3855 498 3864 802
rect 4168 498 4180 802
rect 3855 489 4180 498
rect 3596 442 3692 458
rect 3596 378 3612 442
rect 3676 378 3692 442
rect 3596 362 3692 378
rect 3860 250 4180 489
rect 4315 922 4411 938
rect 4315 858 4331 922
rect 4395 858 4411 922
rect 4315 842 4411 858
rect 4315 778 4331 842
rect 4395 778 4411 842
rect 4580 811 4900 1189
rect 5034 1478 5050 1542
rect 5114 1478 5130 1542
rect 5753 1622 5849 1638
rect 5753 1558 5769 1622
rect 5833 1558 5849 1622
rect 5753 1542 5849 1558
rect 5300 1511 5620 1530
rect 5034 1462 5130 1478
rect 5034 1398 5050 1462
rect 5114 1398 5130 1462
rect 5034 1382 5130 1398
rect 5034 1318 5050 1382
rect 5114 1318 5130 1382
rect 5034 1302 5130 1318
rect 5034 1238 5050 1302
rect 5114 1238 5130 1302
rect 5034 1222 5130 1238
rect 5034 1158 5050 1222
rect 5114 1158 5130 1222
rect 5293 1502 5620 1511
rect 5293 1198 5302 1502
rect 5606 1198 5620 1502
rect 5293 1189 5620 1198
rect 5034 1142 5130 1158
rect 5034 1078 5050 1142
rect 5114 1078 5130 1142
rect 5034 1062 5130 1078
rect 4315 762 4411 778
rect 4315 698 4331 762
rect 4395 698 4411 762
rect 4315 682 4411 698
rect 4315 618 4331 682
rect 4395 618 4411 682
rect 4315 602 4411 618
rect 4315 538 4331 602
rect 4395 538 4411 602
rect 4315 522 4411 538
rect 4315 458 4331 522
rect 4395 458 4411 522
rect 4574 802 4900 811
rect 4574 498 4583 802
rect 4887 498 4900 802
rect 4574 489 4900 498
rect 4315 442 4411 458
rect 4315 378 4331 442
rect 4395 378 4411 442
rect 4315 362 4411 378
rect 4580 250 4900 489
rect 5034 922 5130 938
rect 5034 858 5050 922
rect 5114 858 5130 922
rect 5034 842 5130 858
rect 5034 778 5050 842
rect 5114 778 5130 842
rect 5300 811 5620 1189
rect 5753 1478 5769 1542
rect 5833 1478 5849 1542
rect 6472 1622 6568 1638
rect 6472 1558 6488 1622
rect 6552 1558 6568 1622
rect 6472 1542 6568 1558
rect 6020 1511 6340 1530
rect 5753 1462 5849 1478
rect 5753 1398 5769 1462
rect 5833 1398 5849 1462
rect 5753 1382 5849 1398
rect 5753 1318 5769 1382
rect 5833 1318 5849 1382
rect 5753 1302 5849 1318
rect 5753 1238 5769 1302
rect 5833 1238 5849 1302
rect 5753 1222 5849 1238
rect 5753 1158 5769 1222
rect 5833 1158 5849 1222
rect 6012 1502 6340 1511
rect 6012 1198 6021 1502
rect 6325 1198 6340 1502
rect 6012 1189 6340 1198
rect 5753 1142 5849 1158
rect 5753 1078 5769 1142
rect 5833 1078 5849 1142
rect 5753 1062 5849 1078
rect 5034 762 5130 778
rect 5034 698 5050 762
rect 5114 698 5130 762
rect 5034 682 5130 698
rect 5034 618 5050 682
rect 5114 618 5130 682
rect 5034 602 5130 618
rect 5034 538 5050 602
rect 5114 538 5130 602
rect 5034 522 5130 538
rect 5034 458 5050 522
rect 5114 458 5130 522
rect 5293 802 5620 811
rect 5293 498 5302 802
rect 5606 498 5620 802
rect 5293 489 5620 498
rect 5034 442 5130 458
rect 5034 378 5050 442
rect 5114 378 5130 442
rect 5034 362 5130 378
rect 5300 250 5620 489
rect 5753 922 5849 938
rect 5753 858 5769 922
rect 5833 858 5849 922
rect 5753 842 5849 858
rect 5753 778 5769 842
rect 5833 778 5849 842
rect 6020 811 6340 1189
rect 6472 1478 6488 1542
rect 6552 1478 6568 1542
rect 7191 1622 7287 1638
rect 7191 1558 7207 1622
rect 7271 1558 7287 1622
rect 7191 1542 7287 1558
rect 6740 1511 7060 1530
rect 6472 1462 6568 1478
rect 6472 1398 6488 1462
rect 6552 1398 6568 1462
rect 6472 1382 6568 1398
rect 6472 1318 6488 1382
rect 6552 1318 6568 1382
rect 6472 1302 6568 1318
rect 6472 1238 6488 1302
rect 6552 1238 6568 1302
rect 6472 1222 6568 1238
rect 6472 1158 6488 1222
rect 6552 1158 6568 1222
rect 6731 1502 7060 1511
rect 6731 1198 6740 1502
rect 7044 1198 7060 1502
rect 6731 1189 7060 1198
rect 6472 1142 6568 1158
rect 6472 1078 6488 1142
rect 6552 1078 6568 1142
rect 6472 1062 6568 1078
rect 5753 762 5849 778
rect 5753 698 5769 762
rect 5833 698 5849 762
rect 5753 682 5849 698
rect 5753 618 5769 682
rect 5833 618 5849 682
rect 5753 602 5849 618
rect 5753 538 5769 602
rect 5833 538 5849 602
rect 5753 522 5849 538
rect 5753 458 5769 522
rect 5833 458 5849 522
rect 6012 802 6340 811
rect 6012 498 6021 802
rect 6325 498 6340 802
rect 6012 489 6340 498
rect 5753 442 5849 458
rect 5753 378 5769 442
rect 5833 378 5849 442
rect 5753 362 5849 378
rect 6020 250 6340 489
rect 6472 922 6568 938
rect 6472 858 6488 922
rect 6552 858 6568 922
rect 6472 842 6568 858
rect 6472 778 6488 842
rect 6552 778 6568 842
rect 6740 811 7060 1189
rect 7191 1478 7207 1542
rect 7271 1478 7287 1542
rect 7191 1462 7287 1478
rect 7191 1398 7207 1462
rect 7271 1398 7287 1462
rect 7191 1382 7287 1398
rect 7191 1318 7207 1382
rect 7271 1318 7287 1382
rect 7191 1302 7287 1318
rect 7191 1238 7207 1302
rect 7271 1238 7287 1302
rect 7191 1222 7287 1238
rect 7191 1158 7207 1222
rect 7271 1158 7287 1222
rect 7191 1142 7287 1158
rect 7191 1078 7207 1142
rect 7271 1078 7287 1142
rect 7191 1062 7287 1078
rect 6472 762 6568 778
rect 6472 698 6488 762
rect 6552 698 6568 762
rect 6472 682 6568 698
rect 6472 618 6488 682
rect 6552 618 6568 682
rect 6472 602 6568 618
rect 6472 538 6488 602
rect 6552 538 6568 602
rect 6472 522 6568 538
rect 6472 458 6488 522
rect 6552 458 6568 522
rect 6731 802 7060 811
rect 6731 498 6740 802
rect 7044 498 7060 802
rect 6731 489 7060 498
rect 6472 442 6568 458
rect 6472 378 6488 442
rect 6552 378 6568 442
rect 6472 362 6568 378
rect 6740 250 7060 489
rect 7191 922 7287 938
rect 7191 858 7207 922
rect 7271 858 7287 922
rect 7191 842 7287 858
rect 7191 778 7207 842
rect 7271 778 7287 842
rect 7191 762 7287 778
rect 7191 698 7207 762
rect 7271 698 7287 762
rect 7191 682 7287 698
rect 7191 618 7207 682
rect 7271 618 7287 682
rect 7191 602 7287 618
rect 7191 538 7207 602
rect 7271 538 7287 602
rect 7191 522 7287 538
rect 7191 458 7207 522
rect 7271 458 7287 522
rect 7191 442 7287 458
rect 7191 378 7207 442
rect 7271 378 7287 442
rect 7191 362 7287 378
rect 122 222 7290 250
rect 122 158 150 222
rect 214 158 230 222
rect 294 158 7290 222
rect 122 130 7290 158
<< labels >>
flabel metal2 s 120 1570 320 1650 1 FreeSans 1250 0 0 0 Cin
port 1 nsew
flabel metal4 s 142 140 302 240 1 FreeSans 1250 0 0 0 Cout
port 2 nsew
flabel metal1 s 122 1850 182 1910 1 FreeSans 1250 0 0 0 VPWR
port 3 nsew
flabel metal1 s 122 -30 182 30 1 FreeSans 1250 0 0 0 VGND
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 7411 1880
<< end >>
