magic
tech sky130A
magscale 1 2
timestamp 1483428465
<< checkpaint >>
rect -1260 -1260 62908 21444
<< nwell >>
rect 30591 9642 30703 9963
rect 30870 9642 30959 9963
<< viali >>
rect 27864 9722 27898 9756
rect 29381 9735 29415 9769
rect 29549 9735 29583 9769
rect 29717 9735 29751 9769
rect 29885 9735 29919 9769
rect 30053 9735 30087 9769
rect 30221 9735 30255 9769
rect 30389 9735 30423 9769
rect 31129 9734 31163 9768
rect 31297 9734 31331 9768
rect 31465 9734 31499 9768
rect 31633 9734 31667 9768
rect 31801 9734 31835 9768
rect 31969 9734 32003 9768
rect 32137 9734 32171 9768
rect 27678 9596 27712 9630
rect 28353 9602 28387 9636
rect 28435 9602 28469 9636
rect 28526 9602 28560 9636
rect 28620 9602 28654 9636
rect 28940 9595 28974 9629
rect 29141 9600 29175 9634
rect 29260 9600 29294 9634
rect 29379 9600 29413 9634
rect 29498 9600 29532 9634
rect 29617 9600 29651 9634
rect 29736 9600 29770 9634
rect 29855 9600 29889 9634
rect 31065 9602 31099 9636
rect 31184 9602 31218 9636
rect 31303 9602 31337 9636
rect 31422 9602 31456 9636
rect 31541 9602 31575 9636
rect 31660 9602 31694 9636
rect 31779 9602 31813 9636
<< metal1 >>
rect 427 13891 785 13911
rect 427 13890 727 13891
rect 427 13838 451 13890
rect 503 13839 727 13890
rect 779 13839 785 13891
rect 503 13838 785 13839
rect 427 13814 785 13838
rect 61150 13149 61394 13227
rect 0 12219 29210 12224
rect 0 12167 29120 12219
rect 29172 12167 29210 12219
rect 0 12163 29210 12167
rect 30969 12216 61648 12221
rect 30969 12164 31007 12216
rect 31059 12164 61648 12216
rect 30969 12160 61648 12164
rect 0 12077 27302 12082
rect 0 12025 27232 12077
rect 27284 12025 27302 12077
rect 0 12021 27302 12025
rect 32877 12074 61648 12079
rect 32877 12022 32895 12074
rect 32947 12022 61648 12074
rect 32877 12018 61648 12022
rect 0 11936 25444 11940
rect 0 11884 25345 11936
rect 25397 11884 25444 11936
rect 0 11879 25444 11884
rect 34735 11933 61648 11937
rect 34735 11881 34782 11933
rect 34834 11881 61648 11933
rect 34735 11876 61648 11881
rect 0 11795 23520 11798
rect 0 11743 23456 11795
rect 23508 11743 23520 11795
rect 0 11737 23520 11743
rect 36659 11792 61648 11795
rect 36659 11740 36671 11792
rect 36723 11740 61648 11792
rect 36659 11734 61648 11740
rect 0 11652 21644 11656
rect 0 11600 21568 11652
rect 21620 11600 21644 11652
rect 0 11595 21644 11600
rect 38535 11649 61648 11653
rect 38535 11597 38559 11649
rect 38611 11597 61648 11649
rect 38535 11592 61648 11597
rect 0 11509 19762 11514
rect 0 11457 19678 11509
rect 19730 11457 19762 11509
rect 0 11453 19762 11457
rect 40417 11506 61648 11511
rect 40417 11454 40449 11506
rect 40501 11454 61648 11506
rect 40417 11450 61648 11454
rect 0 11368 17854 11372
rect 0 11316 17792 11368
rect 17844 11316 17854 11368
rect 0 11311 17854 11316
rect 42325 11365 61648 11369
rect 42325 11313 42335 11365
rect 42387 11313 61648 11365
rect 42325 11308 61648 11313
rect 0 11225 15978 11230
rect 0 11173 15904 11225
rect 15956 11173 15978 11225
rect 0 11169 15978 11173
rect 44201 11222 61648 11227
rect 44201 11170 44223 11222
rect 44275 11170 61648 11222
rect 44201 11166 61648 11170
rect 0 11083 14108 11088
rect 0 11031 14023 11083
rect 14075 11031 14108 11083
rect 0 11027 14108 11031
rect 46071 11080 61648 11085
rect 46071 11028 46104 11080
rect 46156 11028 61648 11080
rect 46071 11024 61648 11028
rect 0 10940 12236 10946
rect 0 10888 12135 10940
rect 12187 10888 12236 10940
rect 0 10885 12236 10888
rect 47943 10937 61648 10943
rect 47943 10885 47992 10937
rect 48044 10885 61648 10937
rect 47943 10882 61648 10885
rect 0 10798 10350 10804
rect 0 10746 10247 10798
rect 10299 10746 10350 10798
rect 0 10743 10350 10746
rect 49829 10800 59808 10801
rect 61176 10800 61648 10801
rect 49829 10795 61648 10800
rect 49829 10743 49880 10795
rect 49932 10743 61648 10795
rect 49829 10740 61648 10743
rect 59711 10739 61648 10740
rect 0 10656 8439 10662
rect 0 10604 8360 10656
rect 8412 10604 8439 10656
rect 0 10601 8439 10604
rect 51740 10653 61648 10659
rect 51740 10601 51767 10653
rect 51819 10601 61648 10653
rect 51740 10598 61648 10601
rect 0 10515 6563 10520
rect 0 10463 6470 10515
rect 6522 10463 6563 10515
rect 0 10459 6563 10463
rect 53616 10512 61648 10517
rect 53616 10460 53657 10512
rect 53709 10460 61648 10512
rect 53616 10456 61648 10460
rect 0 10373 4666 10378
rect 0 10321 4583 10373
rect 4635 10321 4666 10373
rect 0 10317 4666 10321
rect 55513 10370 61648 10375
rect 55513 10318 55544 10370
rect 55596 10318 61648 10370
rect 55513 10314 61648 10318
rect 0 10230 2794 10236
rect 0 10178 2694 10230
rect 2746 10178 2794 10230
rect 0 10175 2794 10178
rect 57385 10227 61648 10233
rect 57385 10175 57433 10227
rect 57485 10175 61648 10227
rect 57385 10172 61648 10175
rect 0 10089 935 10094
rect 0 10037 806 10089
rect 858 10037 935 10089
rect 0 10033 935 10037
rect 59244 10086 61648 10091
rect 59244 10034 59321 10086
rect 59373 10034 61648 10086
rect 59244 10030 61648 10034
rect 0 9947 1157 9952
rect 0 9895 1033 9947
rect 1085 9895 1157 9947
rect 0 9891 1157 9895
rect 28101 9877 28177 9973
rect 29005 9877 29081 9973
rect 30553 9877 30740 9973
rect 30832 9877 31019 9973
rect 59479 9944 61648 9949
rect 59479 9892 59551 9944
rect 59603 9892 61648 9944
rect 59479 9888 61648 9892
rect 0 9808 3016 9810
rect 0 9756 2920 9808
rect 2972 9756 3016 9808
rect 57620 9805 61648 9807
rect 0 9749 3016 9756
rect 27854 9756 27907 9773
rect 27854 9722 27864 9756
rect 27898 9722 27907 9756
rect 0 9663 4927 9668
rect 0 9611 4809 9663
rect 4861 9611 4927 9663
rect 0 9607 4927 9611
rect 7162 9652 7509 9674
rect 7162 9640 27730 9652
rect 7162 9588 7251 9640
rect 7303 9588 7349 9640
rect 7401 9630 27730 9640
rect 7401 9596 27678 9630
rect 27712 9596 27730 9630
rect 7401 9588 27730 9596
rect 27854 9651 27907 9722
rect 29369 9769 32186 9794
rect 29369 9735 29381 9769
rect 29415 9735 29549 9769
rect 29583 9735 29717 9769
rect 29751 9735 29885 9769
rect 29919 9735 30053 9769
rect 30087 9735 30221 9769
rect 30255 9735 30389 9769
rect 30423 9768 32186 9769
rect 30423 9760 31129 9768
rect 30423 9735 30601 9760
rect 29369 9708 30601 9735
rect 30653 9708 30704 9760
rect 30756 9708 30807 9760
rect 30859 9708 30910 9760
rect 30962 9734 31129 9760
rect 31163 9734 31297 9768
rect 31331 9734 31465 9768
rect 31499 9734 31633 9768
rect 31667 9734 31801 9768
rect 31835 9734 31969 9768
rect 32003 9734 32137 9768
rect 32171 9734 32186 9768
rect 57620 9753 57664 9805
rect 57716 9753 61648 9805
rect 57620 9746 61648 9753
rect 30962 9708 32186 9734
rect 29369 9686 32186 9708
rect 55709 9660 61648 9665
rect 27854 9636 28699 9651
rect 27854 9602 28353 9636
rect 28387 9602 28435 9636
rect 28469 9602 28526 9636
rect 28560 9602 28620 9636
rect 28654 9602 28699 9636
rect 27854 9590 28699 9602
rect 28918 9636 32109 9645
rect 28918 9634 31065 9636
rect 28918 9629 29141 9634
rect 28918 9595 28940 9629
rect 28974 9600 29141 9629
rect 29175 9600 29260 9634
rect 29294 9600 29379 9634
rect 29413 9600 29498 9634
rect 29532 9600 29617 9634
rect 29651 9600 29736 9634
rect 29770 9600 29855 9634
rect 29889 9602 31065 9634
rect 31099 9602 31184 9636
rect 31218 9602 31303 9636
rect 31337 9602 31422 9636
rect 31456 9602 31541 9636
rect 31575 9602 31660 9636
rect 31694 9602 31779 9636
rect 31813 9602 32109 9636
rect 55709 9608 55775 9660
rect 55827 9608 61648 9660
rect 55709 9604 61648 9608
rect 29889 9600 32109 9602
rect 28974 9595 32109 9600
rect 28918 9588 32109 9595
rect 7162 9578 27730 9588
rect 7162 9550 7509 9578
rect 0 9522 6773 9526
rect 0 9470 6698 9522
rect 6750 9470 6773 9522
rect 0 9465 6773 9470
rect 53863 9519 61648 9523
rect 53863 9467 53886 9519
rect 53938 9467 61648 9519
rect 53863 9462 61648 9467
rect 0 9378 8664 9384
rect 0 9326 8585 9378
rect 8637 9326 8664 9378
rect 28101 9333 28177 9429
rect 29005 9332 29081 9428
rect 30553 9333 30740 9429
rect 30832 9333 31019 9429
rect 51972 9375 61648 9381
rect 0 9323 8664 9326
rect 51972 9323 51999 9375
rect 52051 9323 61648 9375
rect 51972 9320 61648 9323
rect 0 9237 10552 9242
rect 0 9185 10473 9237
rect 10525 9185 10552 9237
rect 0 9181 10552 9185
rect 50084 9234 61648 9239
rect 50084 9182 50111 9234
rect 50163 9182 61648 9234
rect 50084 9178 61648 9182
rect 0 9095 12453 9100
rect 0 9043 12362 9095
rect 12414 9043 12453 9095
rect 0 9039 12453 9043
rect 48183 9092 61648 9097
rect 48183 9040 48222 9092
rect 48274 9040 61648 9092
rect 48183 9036 61648 9040
rect 0 8950 14328 8958
rect 0 8898 14250 8950
rect 14302 8898 14328 8950
rect 0 8897 14328 8898
rect 46308 8947 61648 8955
rect 46308 8895 46334 8947
rect 46386 8895 61648 8947
rect 46308 8894 61648 8895
rect 0 8811 16239 8816
rect 0 8759 16128 8811
rect 16180 8759 16239 8811
rect 0 8755 16239 8759
rect 44397 8808 61648 8813
rect 44397 8756 44456 8808
rect 44508 8756 61648 8808
rect 44397 8752 61648 8756
rect 0 8670 18137 8674
rect 0 8618 18019 8670
rect 18071 8618 18137 8670
rect 0 8613 18137 8618
rect 42499 8667 61648 8671
rect 42499 8615 42565 8667
rect 42617 8615 61648 8667
rect 42499 8610 61648 8615
rect 0 8529 20044 8532
rect 0 8477 19904 8529
rect 19956 8477 20044 8529
rect 0 8471 20044 8477
rect 40592 8526 61648 8529
rect 40592 8474 40680 8526
rect 40732 8474 61648 8526
rect 40592 8468 61648 8474
rect 0 8386 21894 8390
rect 0 8334 21795 8386
rect 21847 8334 21894 8386
rect 0 8329 21894 8334
rect 38742 8383 61648 8387
rect 38742 8331 38789 8383
rect 38841 8331 61648 8383
rect 38742 8326 61648 8331
rect 0 8243 23769 8248
rect 0 8191 23685 8243
rect 23737 8191 23769 8243
rect 0 8187 23769 8191
rect 36867 8240 61648 8245
rect 36867 8188 36899 8240
rect 36951 8188 61648 8240
rect 36867 8184 61648 8188
rect 0 8099 25666 8106
rect 0 8047 25568 8099
rect 25620 8047 25666 8099
rect 0 8045 25666 8047
rect 34970 8096 61648 8103
rect 34970 8044 35016 8096
rect 35068 8044 61648 8096
rect 34970 8042 61648 8044
rect 0 7957 27596 7964
rect 0 7905 27458 7957
rect 27510 7905 27596 7957
rect 0 7903 27596 7905
rect 33040 7954 61648 7961
rect 33040 7902 33126 7954
rect 33178 7902 61648 7954
rect 33040 7900 61648 7902
rect 0 7817 29446 7822
rect 0 7765 29350 7817
rect 29402 7765 29446 7817
rect 0 7761 29446 7765
rect 31190 7814 61648 7819
rect 31190 7762 31234 7814
rect 31286 7762 61648 7814
rect 31190 7758 61648 7762
rect 174 6112 955 6127
rect 174 6104 896 6112
rect 174 6052 191 6104
rect 243 6060 896 6104
rect 948 6060 955 6112
rect 243 6052 955 6060
rect 174 6034 955 6052
<< via1 >>
rect 30637 15452 30689 15504
rect 30754 15452 30806 15504
rect 30871 15452 30923 15504
rect 451 13838 503 13890
rect 727 13839 779 13891
rect 29120 12167 29172 12219
rect 31007 12164 31059 12216
rect 27232 12025 27284 12077
rect 32895 12022 32947 12074
rect 25345 11884 25397 11936
rect 34782 11881 34834 11933
rect 23456 11743 23508 11795
rect 36671 11740 36723 11792
rect 21568 11600 21620 11652
rect 38559 11597 38611 11649
rect 19678 11457 19730 11509
rect 40449 11454 40501 11506
rect 17792 11316 17844 11368
rect 42335 11313 42387 11365
rect 15904 11173 15956 11225
rect 44223 11170 44275 11222
rect 14023 11031 14075 11083
rect 46104 11028 46156 11080
rect 12135 10888 12187 10940
rect 47992 10885 48044 10937
rect 10247 10746 10299 10798
rect 49880 10743 49932 10795
rect 8360 10604 8412 10656
rect 51767 10601 51819 10653
rect 6470 10463 6522 10515
rect 53657 10460 53709 10512
rect 4583 10321 4635 10373
rect 55544 10318 55596 10370
rect 2694 10178 2746 10230
rect 57433 10175 57485 10227
rect 806 10037 858 10089
rect 59321 10034 59373 10086
rect 1033 9895 1085 9947
rect 31704 9891 31756 9943
rect 31834 9891 31886 9943
rect 31964 9891 32016 9943
rect 59551 9892 59603 9944
rect 2920 9756 2972 9808
rect 4809 9611 4861 9663
rect 7251 9588 7303 9640
rect 7349 9588 7401 9640
rect 30601 9708 30653 9760
rect 30704 9708 30756 9760
rect 30807 9708 30859 9760
rect 30910 9708 30962 9760
rect 57664 9753 57716 9805
rect 55775 9608 55827 9660
rect 6698 9470 6750 9522
rect 53886 9467 53938 9519
rect 8585 9326 8637 9378
rect 31694 9361 31746 9413
rect 31807 9361 31859 9413
rect 31920 9361 31972 9413
rect 32033 9361 32085 9413
rect 32146 9361 32198 9413
rect 51999 9323 52051 9375
rect 10473 9185 10525 9237
rect 50111 9182 50163 9234
rect 12362 9043 12414 9095
rect 48222 9040 48274 9092
rect 14250 8898 14302 8950
rect 46334 8895 46386 8947
rect 16128 8759 16180 8811
rect 44456 8756 44508 8808
rect 18019 8618 18071 8670
rect 42565 8615 42617 8667
rect 19904 8477 19956 8529
rect 40680 8474 40732 8526
rect 21795 8334 21847 8386
rect 38789 8331 38841 8383
rect 23685 8191 23737 8243
rect 36899 8188 36951 8240
rect 25568 8047 25620 8099
rect 35016 8044 35068 8096
rect 27458 7905 27510 7957
rect 33126 7902 33178 7954
rect 29350 7765 29402 7817
rect 31234 7762 31286 7814
rect 31694 7472 31746 7524
rect 31807 7472 31859 7524
rect 31920 7472 31972 7524
rect 32033 7472 32085 7524
rect 32146 7472 32198 7524
rect 31694 7367 31746 7419
rect 31807 7367 31859 7419
rect 31920 7367 31972 7419
rect 32033 7367 32085 7419
rect 32146 7367 32198 7419
rect 191 6052 243 6104
rect 896 6060 948 6112
rect 30626 3223 30678 3275
rect 30709 3223 30761 3275
rect 30792 3223 30844 3275
rect 30875 3223 30927 3275
<< metal2 >>
rect 2180 19017 2224 20184
rect 4068 19017 4112 19992
rect 5956 19017 6000 19992
rect 7844 19017 7888 19992
rect 9732 19017 9776 19992
rect 11620 19017 11664 19992
rect 13508 19017 13552 19992
rect 15396 19017 15440 19992
rect 17284 19017 17328 19992
rect 19172 19017 19216 19992
rect 21060 19017 21104 19992
rect 22948 19017 22992 19992
rect 24836 19017 24880 19992
rect 26724 19017 26768 19992
rect 28612 19017 28656 19992
rect 30500 19017 30544 19992
rect 32388 19017 32432 19992
rect 34276 19017 34320 19992
rect 36164 19017 36208 19992
rect 38052 19017 38096 19992
rect 39940 19017 39984 19992
rect 41828 19017 41872 19992
rect 43716 19017 43760 19992
rect 45604 19017 45648 19992
rect 47492 19017 47536 19992
rect 49380 19017 49424 20151
rect 51268 19017 51312 19992
rect 53156 19017 53200 19992
rect 55044 19017 55088 19992
rect 56932 19017 56976 19992
rect 58820 19017 58864 19992
rect 60708 19017 60752 19992
rect 61283 18335 61319 18368
rect 182 18299 896 18335
rect 60572 18299 61319 18335
rect 182 6127 218 18299
rect 30573 15559 30969 15588
rect 30573 15503 30604 15559
rect 30660 15504 30713 15559
rect 30769 15504 30822 15559
rect 30878 15504 30969 15559
rect 30689 15503 30713 15504
rect 30806 15503 30822 15504
rect 30573 15457 30637 15503
rect 30689 15457 30754 15503
rect 30806 15457 30871 15503
rect 30573 15401 30604 15457
rect 30689 15452 30713 15457
rect 30806 15452 30822 15457
rect 30923 15452 30969 15504
rect 30660 15401 30713 15452
rect 30769 15401 30822 15452
rect 30878 15401 30969 15452
rect 30573 15380 30969 15401
rect 416 13890 514 13917
rect 416 13838 451 13890
rect 503 13838 514 13890
rect 416 13798 514 13838
rect 714 13891 818 13914
rect 714 13839 727 13891
rect 779 13879 818 13891
rect 61283 13879 61319 18299
rect 779 13843 990 13879
rect 60666 13843 61319 13879
rect 779 13839 818 13843
rect 714 13814 818 13839
rect 181 6104 292 6127
rect 181 6052 191 6104
rect 243 6052 292 6104
rect 181 6012 292 6052
rect 448 1648 484 13798
rect 810 10099 854 13161
rect 2698 10242 2742 13161
rect 4586 10382 4630 13161
rect 6474 10526 6518 13161
rect 8362 10666 8406 13161
rect 10250 10808 10294 12753
rect 12138 10950 12182 12773
rect 14026 11092 14070 12763
rect 15908 11233 15952 12770
rect 17796 11374 17840 12823
rect 19684 11519 19728 12763
rect 21572 11662 21616 12743
rect 23460 11804 23504 12743
rect 25348 11945 25392 12703
rect 27236 12088 27280 12747
rect 29124 12234 29168 12757
rect 29101 12219 29195 12234
rect 31011 12231 31055 12596
rect 29101 12167 29120 12219
rect 29172 12167 29195 12219
rect 29101 12153 29195 12167
rect 30984 12216 31078 12231
rect 30984 12164 31007 12216
rect 31059 12164 31078 12216
rect 29124 12109 29168 12153
rect 30984 12150 31078 12164
rect 31011 12106 31055 12150
rect 27221 12077 27298 12088
rect 32899 12085 32943 12617
rect 27221 12025 27232 12077
rect 27284 12025 27298 12077
rect 27221 12015 27298 12025
rect 32881 12074 32958 12085
rect 32881 12022 32895 12074
rect 32947 12022 32958 12074
rect 27236 11972 27280 12015
rect 32881 12012 32958 12022
rect 32899 11969 32943 12012
rect 25332 11936 25409 11945
rect 34787 11942 34831 12673
rect 25332 11884 25345 11936
rect 25397 11884 25409 11936
rect 25332 11872 25409 11884
rect 34770 11933 34847 11942
rect 34770 11881 34782 11933
rect 34834 11881 34847 11933
rect 25348 11842 25392 11872
rect 34770 11869 34847 11881
rect 34787 11839 34831 11869
rect 23445 11795 23522 11804
rect 36675 11801 36719 12598
rect 23445 11743 23456 11795
rect 23508 11743 23522 11795
rect 23445 11731 23522 11743
rect 36657 11792 36734 11801
rect 36657 11740 36671 11792
rect 36723 11740 36734 11792
rect 23460 11695 23504 11731
rect 36657 11728 36734 11740
rect 36675 11692 36719 11728
rect 21556 11652 21633 11662
rect 38563 11659 38607 12608
rect 21556 11600 21568 11652
rect 21620 11600 21633 11652
rect 21556 11589 21633 11600
rect 38546 11649 38623 11659
rect 38546 11597 38559 11649
rect 38611 11597 38623 11649
rect 21572 11555 21616 11589
rect 38546 11586 38623 11597
rect 38563 11552 38607 11586
rect 19670 11509 19747 11519
rect 40451 11516 40495 12636
rect 19670 11457 19678 11509
rect 19730 11457 19747 11509
rect 19670 11446 19747 11457
rect 40432 11506 40509 11516
rect 40432 11454 40449 11506
rect 40501 11454 40509 11506
rect 19684 11404 19728 11446
rect 40432 11443 40509 11454
rect 40451 11401 40495 11443
rect 17779 11368 17856 11374
rect 42339 11371 42383 12629
rect 17779 11316 17792 11368
rect 17844 11316 17856 11368
rect 17779 11301 17856 11316
rect 42323 11365 42400 11371
rect 42323 11313 42335 11365
rect 42387 11313 42400 11365
rect 17796 11258 17840 11301
rect 42323 11298 42400 11313
rect 42339 11255 42383 11298
rect 15892 11225 15969 11233
rect 44227 11230 44271 12627
rect 15892 11173 15904 11225
rect 15956 11173 15969 11225
rect 15892 11160 15969 11173
rect 44210 11222 44287 11230
rect 44210 11170 44223 11222
rect 44275 11170 44287 11222
rect 15908 11131 15952 11160
rect 44210 11157 44287 11170
rect 44227 11128 44271 11157
rect 14011 11083 14088 11092
rect 46109 11089 46153 12595
rect 14011 11031 14023 11083
rect 14075 11031 14088 11083
rect 14011 11019 14088 11031
rect 46091 11080 46168 11089
rect 46091 11028 46104 11080
rect 46156 11028 46168 11080
rect 14026 10991 14070 11019
rect 46091 11016 46168 11028
rect 46109 10988 46153 11016
rect 12123 10940 12200 10950
rect 47997 10947 48041 12633
rect 12123 10888 12135 10940
rect 12187 10888 12200 10940
rect 12123 10877 12200 10888
rect 47979 10937 48056 10947
rect 47979 10885 47992 10937
rect 48044 10885 48056 10937
rect 12138 10854 12182 10877
rect 47979 10874 48056 10885
rect 47997 10851 48041 10874
rect 10234 10798 10311 10808
rect 49885 10805 49929 12618
rect 10234 10746 10247 10798
rect 10299 10746 10311 10798
rect 10234 10735 10311 10746
rect 49868 10795 49945 10805
rect 49868 10743 49880 10795
rect 49932 10743 49945 10795
rect 10250 10697 10294 10735
rect 49868 10732 49945 10743
rect 49885 10694 49929 10732
rect 8348 10656 8425 10666
rect 51773 10663 51817 12618
rect 8348 10604 8360 10656
rect 8412 10604 8425 10656
rect 8348 10593 8425 10604
rect 51754 10653 51831 10663
rect 51754 10601 51767 10653
rect 51819 10601 51831 10653
rect 8362 10560 8406 10593
rect 51754 10590 51831 10601
rect 51773 10557 51817 10590
rect 6460 10515 6537 10526
rect 53661 10523 53705 12631
rect 6460 10463 6470 10515
rect 6522 10463 6537 10515
rect 6460 10453 6537 10463
rect 53642 10512 53719 10523
rect 53642 10460 53657 10512
rect 53709 10460 53719 10512
rect 6474 10417 6518 10453
rect 53642 10450 53719 10460
rect 4570 10373 4647 10382
rect 4570 10321 4583 10373
rect 4635 10321 4647 10373
rect 4570 10309 4647 10321
rect 30574 10377 30971 10416
rect 53661 10414 53705 10450
rect 55549 10379 55593 12648
rect 30574 10321 30597 10377
rect 30653 10321 30701 10377
rect 30757 10321 30805 10377
rect 30861 10321 30909 10377
rect 30965 10321 30971 10377
rect 4586 10270 4630 10309
rect 30574 10278 30971 10321
rect 55532 10370 55609 10379
rect 55532 10318 55544 10370
rect 55596 10318 55609 10370
rect 55532 10306 55609 10318
rect 2686 10230 2763 10242
rect 2686 10178 2694 10230
rect 2746 10178 2763 10230
rect 2686 10169 2763 10178
rect 30574 10222 30597 10278
rect 30653 10222 30701 10278
rect 30757 10222 30805 10278
rect 30861 10222 30909 10278
rect 30965 10222 30971 10278
rect 55549 10267 55593 10306
rect 57437 10239 57481 12646
rect 2698 10133 2742 10169
rect 793 10089 870 10099
rect 793 10037 806 10089
rect 858 10037 870 10089
rect 793 10026 870 10037
rect 810 10003 854 10026
rect 1039 9958 1083 9988
rect 1022 9947 1101 9958
rect 1022 9895 1033 9947
rect 1085 9895 1101 9947
rect 1022 9882 1101 9895
rect 1039 7250 1083 9882
rect 2927 9817 2971 9861
rect 2908 9808 2987 9817
rect 2908 9756 2920 9808
rect 2972 9756 2987 9808
rect 2908 9741 2987 9756
rect 30574 9760 30971 10222
rect 57416 10227 57493 10239
rect 57416 10175 57433 10227
rect 57485 10175 57493 10227
rect 57416 10166 57493 10175
rect 57437 10130 57481 10166
rect 59325 10096 59369 12644
rect 59309 10086 59386 10096
rect 59309 10034 59321 10086
rect 59373 10034 59386 10086
rect 59309 10023 59386 10034
rect 59325 10000 59369 10023
rect 31665 9947 32066 9972
rect 59553 9955 59597 9985
rect 31665 9891 31704 9947
rect 31760 9891 31833 9947
rect 31889 9891 31962 9947
rect 32018 9891 32066 9947
rect 31665 9878 32066 9891
rect 59535 9944 59614 9955
rect 59535 9892 59551 9944
rect 59603 9892 59614 9944
rect 59535 9879 59614 9892
rect 57665 9814 57709 9858
rect 2927 7204 2971 9741
rect 4815 9671 4859 9744
rect 30574 9708 30601 9760
rect 30653 9708 30704 9760
rect 30756 9708 30807 9760
rect 30859 9708 30910 9760
rect 30962 9708 30971 9760
rect 57649 9805 57728 9814
rect 57649 9753 57664 9805
rect 57716 9753 57728 9805
rect 4790 9663 4869 9671
rect 4790 9611 4809 9663
rect 4861 9611 4869 9663
rect 4790 9595 4869 9611
rect 7162 9644 7509 9674
rect 7162 9640 7252 9644
rect 4815 7167 4859 9595
rect 6703 9530 6747 9604
rect 7162 9588 7251 9640
rect 7308 9588 7349 9644
rect 7405 9588 7509 9644
rect 7162 9550 7509 9588
rect 6685 9522 6764 9530
rect 6685 9470 6698 9522
rect 6750 9470 6764 9522
rect 6685 9454 6764 9470
rect 6703 7216 6747 9454
rect 8591 9389 8635 9438
rect 8574 9378 8653 9389
rect 8574 9326 8585 9378
rect 8637 9326 8653 9378
rect 8574 9313 8653 9326
rect 8591 7253 8635 9313
rect 10479 9247 10523 9292
rect 10462 9237 10541 9247
rect 10462 9185 10473 9237
rect 10525 9185 10541 9237
rect 10462 9171 10541 9185
rect 10479 7216 10523 9171
rect 12367 9104 12411 9145
rect 12351 9095 12430 9104
rect 12351 9043 12362 9095
rect 12414 9043 12430 9095
rect 12351 9028 12430 9043
rect 30574 9048 30971 9708
rect 55777 9668 55821 9741
rect 57649 9738 57728 9753
rect 55767 9660 55846 9668
rect 55767 9608 55775 9660
rect 55827 9608 55846 9660
rect 53889 9527 53933 9601
rect 55767 9592 55846 9608
rect 53872 9519 53951 9527
rect 53872 9467 53886 9519
rect 53938 9467 53951 9519
rect 53872 9451 53951 9467
rect 12367 7192 12411 9028
rect 30574 8992 30610 9048
rect 30666 8992 30698 9048
rect 30754 8992 30786 9048
rect 30842 8992 30874 9048
rect 30930 8992 30971 9048
rect 14255 8959 14299 8986
rect 14239 8950 14318 8959
rect 14239 8898 14250 8950
rect 14302 8898 14318 8950
rect 14239 8883 14318 8898
rect 30574 8953 30971 8992
rect 30574 8897 30610 8953
rect 30666 8897 30698 8953
rect 30754 8897 30786 8953
rect 30842 8897 30874 8953
rect 30930 8897 30971 8953
rect 14255 7216 14299 8883
rect 30574 8866 30971 8897
rect 31639 9413 32306 9430
rect 31639 9361 31694 9413
rect 31746 9361 31807 9413
rect 31859 9361 31920 9413
rect 31972 9361 32033 9413
rect 32085 9361 32146 9413
rect 32198 9361 32306 9413
rect 52001 9386 52045 9435
rect 16137 8821 16181 8863
rect 16117 8811 16196 8821
rect 16117 8759 16128 8811
rect 16180 8759 16196 8811
rect 16117 8745 16196 8759
rect 16137 7161 16181 8745
rect 18025 8679 18069 8735
rect 18007 8670 18086 8679
rect 18007 8618 18019 8670
rect 18071 8618 18086 8670
rect 18007 8603 18086 8618
rect 18025 7192 18069 8603
rect 19913 8538 19957 8594
rect 19893 8529 19972 8538
rect 19893 8477 19904 8529
rect 19956 8477 19972 8529
rect 19893 8462 19972 8477
rect 19913 7234 19957 8462
rect 21801 8396 21845 8453
rect 21783 8386 21862 8396
rect 21783 8334 21795 8386
rect 21847 8334 21862 8386
rect 21783 8320 21862 8334
rect 21801 7210 21845 8320
rect 23689 8253 23733 8319
rect 23673 8243 23752 8253
rect 23673 8191 23685 8243
rect 23737 8191 23752 8243
rect 23673 8177 23752 8191
rect 23689 7161 23733 8177
rect 25577 8112 25621 8166
rect 25555 8099 25634 8112
rect 25555 8047 25568 8099
rect 25620 8047 25634 8099
rect 25555 8036 25634 8047
rect 25577 7192 25621 8036
rect 27465 7970 27509 8007
rect 27449 7957 27528 7970
rect 27449 7905 27458 7957
rect 27510 7905 27528 7957
rect 27449 7894 27528 7905
rect 27465 7192 27509 7894
rect 29353 7828 29397 7903
rect 29339 7817 29418 7828
rect 31239 7825 31283 7900
rect 29339 7765 29350 7817
rect 29402 7765 29418 7817
rect 29339 7752 29418 7765
rect 31218 7814 31297 7825
rect 31218 7762 31234 7814
rect 31286 7762 31297 7814
rect 29353 7198 29397 7752
rect 31218 7749 31297 7762
rect 31239 7293 31283 7749
rect 31639 7524 32306 9361
rect 51983 9375 52062 9386
rect 51983 9323 51999 9375
rect 52051 9323 52062 9375
rect 51983 9310 52062 9323
rect 50113 9244 50157 9289
rect 50095 9234 50174 9244
rect 50095 9182 50111 9234
rect 50163 9182 50174 9234
rect 50095 9168 50174 9182
rect 48225 9101 48269 9142
rect 48206 9092 48285 9101
rect 48206 9040 48222 9092
rect 48274 9040 48285 9092
rect 48206 9025 48285 9040
rect 46337 8956 46381 8983
rect 46318 8947 46397 8956
rect 46318 8895 46334 8947
rect 46386 8895 46397 8947
rect 46318 8880 46397 8895
rect 44455 8818 44499 8860
rect 44440 8808 44519 8818
rect 44440 8756 44456 8808
rect 44508 8756 44519 8808
rect 44440 8742 44519 8756
rect 42567 8676 42611 8732
rect 42550 8667 42629 8676
rect 42550 8615 42565 8667
rect 42617 8615 42629 8667
rect 42550 8600 42629 8615
rect 40679 8535 40723 8591
rect 40664 8526 40743 8535
rect 40664 8474 40680 8526
rect 40732 8474 40743 8526
rect 40664 8459 40743 8474
rect 38791 8393 38835 8450
rect 38774 8383 38853 8393
rect 38774 8331 38789 8383
rect 38841 8331 38853 8383
rect 38774 8317 38853 8331
rect 36903 8250 36947 8316
rect 36884 8240 36963 8250
rect 36884 8188 36899 8240
rect 36951 8188 36963 8240
rect 36884 8174 36963 8188
rect 35015 8109 35059 8163
rect 35002 8096 35081 8109
rect 35002 8044 35016 8096
rect 35068 8044 35081 8096
rect 35002 8033 35081 8044
rect 33127 7967 33171 8004
rect 33108 7954 33187 7967
rect 33108 7902 33126 7954
rect 33178 7902 33187 7954
rect 33108 7891 33187 7902
rect 31639 7472 31694 7524
rect 31746 7472 31807 7524
rect 31859 7472 31920 7524
rect 31972 7472 32033 7524
rect 32085 7472 32146 7524
rect 32198 7472 32306 7524
rect 31639 7419 32306 7472
rect 31639 7367 31694 7419
rect 31746 7367 31807 7419
rect 31859 7367 31920 7419
rect 31972 7367 32033 7419
rect 32085 7367 32146 7419
rect 32198 7367 32306 7419
rect 31639 7319 32306 7367
rect 33127 7340 33171 7891
rect 35015 7302 35059 8033
rect 36903 7299 36947 8174
rect 38791 7293 38835 8317
rect 40679 7319 40723 8459
rect 42567 7244 42611 8600
rect 44455 7287 44499 8742
rect 46337 7306 46381 8880
rect 48225 7270 48269 9025
rect 50113 7259 50157 9168
rect 52001 7285 52045 9310
rect 53889 7310 53933 9451
rect 55777 7268 55821 9592
rect 57665 7329 57709 9738
rect 59553 7299 59597 9879
rect 889 6112 959 6133
rect 889 6060 896 6112
rect 948 6104 959 6112
rect 948 6068 1219 6104
rect 60895 6068 61620 6104
rect 948 6060 959 6068
rect 889 6029 959 6060
rect 30574 3324 30971 3357
rect 30574 3268 30615 3324
rect 30671 3275 30707 3324
rect 30763 3275 30799 3324
rect 30855 3275 30891 3324
rect 30678 3268 30707 3275
rect 30763 3268 30792 3275
rect 30855 3268 30875 3275
rect 30947 3268 30971 3324
rect 30574 3233 30626 3268
rect 30678 3233 30709 3268
rect 30761 3233 30792 3268
rect 30844 3233 30875 3268
rect 30927 3233 30971 3268
rect 30574 3177 30615 3233
rect 30678 3223 30707 3233
rect 30763 3223 30792 3233
rect 30855 3223 30875 3233
rect 30671 3177 30707 3223
rect 30763 3177 30799 3223
rect 30855 3177 30891 3223
rect 30947 3177 30971 3233
rect 30574 3151 30971 3177
rect 61584 1648 61620 6068
rect 448 1612 1125 1648
rect 60801 1612 61620 1648
rect 61584 1601 61620 1612
rect 2409 0 2465 930
rect 4297 0 4353 930
rect 6185 0 6241 930
rect 8073 0 8129 930
rect 9961 0 10017 930
rect 11849 0 11905 930
rect 13737 0 13793 930
rect 15625 0 15681 930
rect 17513 0 17569 930
rect 19401 0 19457 930
rect 21289 0 21345 930
rect 23177 0 23233 930
rect 25065 0 25121 930
rect 26953 0 27009 930
rect 28841 0 28897 930
rect 30729 0 30785 930
rect 32617 0 32673 930
rect 34505 0 34561 930
rect 36393 0 36449 930
rect 38281 0 38337 930
rect 40169 0 40225 930
rect 42057 0 42113 930
rect 43945 0 44001 930
rect 45833 0 45889 930
rect 47721 0 47777 930
rect 49609 0 49665 930
rect 51497 0 51553 930
rect 53385 0 53441 930
rect 55273 0 55329 930
rect 57161 0 57217 930
rect 59049 0 59105 930
rect 60937 0 60993 930
<< via2 >>
rect 30604 15504 30660 15559
rect 30713 15504 30769 15559
rect 30822 15504 30878 15559
rect 30604 15503 30637 15504
rect 30637 15503 30660 15504
rect 30713 15503 30754 15504
rect 30754 15503 30769 15504
rect 30822 15503 30871 15504
rect 30871 15503 30878 15504
rect 30604 15452 30637 15457
rect 30637 15452 30660 15457
rect 30713 15452 30754 15457
rect 30754 15452 30769 15457
rect 30822 15452 30871 15457
rect 30871 15452 30878 15457
rect 30604 15401 30660 15452
rect 30713 15401 30769 15452
rect 30822 15401 30878 15452
rect 30597 10321 30653 10377
rect 30701 10321 30757 10377
rect 30805 10321 30861 10377
rect 30909 10321 30965 10377
rect 30597 10222 30653 10278
rect 30701 10222 30757 10278
rect 30805 10222 30861 10278
rect 30909 10222 30965 10278
rect 31704 9943 31760 9947
rect 31704 9891 31756 9943
rect 31756 9891 31760 9943
rect 31833 9943 31889 9947
rect 31833 9891 31834 9943
rect 31834 9891 31886 9943
rect 31886 9891 31889 9943
rect 31962 9943 32018 9947
rect 31962 9891 31964 9943
rect 31964 9891 32016 9943
rect 32016 9891 32018 9943
rect 7252 9640 7308 9644
rect 7252 9588 7303 9640
rect 7303 9588 7308 9640
rect 7349 9640 7405 9644
rect 7349 9588 7401 9640
rect 7401 9588 7405 9640
rect 30610 8992 30666 9048
rect 30698 8992 30754 9048
rect 30786 8992 30842 9048
rect 30874 8992 30930 9048
rect 30610 8897 30666 8953
rect 30698 8897 30754 8953
rect 30786 8897 30842 8953
rect 30874 8897 30930 8953
rect 30615 3275 30671 3324
rect 30707 3275 30763 3324
rect 30799 3275 30855 3324
rect 30891 3275 30947 3324
rect 30615 3268 30626 3275
rect 30626 3268 30671 3275
rect 30707 3268 30709 3275
rect 30709 3268 30761 3275
rect 30761 3268 30763 3275
rect 30799 3268 30844 3275
rect 30844 3268 30855 3275
rect 30891 3268 30927 3275
rect 30927 3268 30947 3275
rect 30615 3223 30626 3233
rect 30626 3223 30671 3233
rect 30707 3223 30709 3233
rect 30709 3223 30761 3233
rect 30761 3223 30763 3233
rect 30799 3223 30844 3233
rect 30844 3223 30855 3233
rect 30891 3223 30927 3233
rect 30927 3223 30947 3233
rect 30615 3177 30671 3223
rect 30707 3177 30763 3223
rect 30799 3177 30855 3223
rect 30891 3177 30947 3223
<< metal3 >>
rect 20135 19764 20241 19781
rect 20135 19700 20156 19764
rect 20220 19700 20241 19764
rect 20135 19684 20241 19700
rect 20135 19620 20156 19684
rect 20220 19620 20241 19684
rect 20135 19603 20241 19620
rect 20309 19764 20415 19781
rect 20309 19700 20330 19764
rect 20394 19700 20415 19764
rect 20309 19684 20415 19700
rect 20309 19620 20330 19684
rect 20394 19620 20415 19684
rect 20309 19603 20415 19620
rect 20483 19764 20589 19781
rect 20483 19700 20504 19764
rect 20568 19700 20589 19764
rect 20483 19684 20589 19700
rect 20483 19620 20504 19684
rect 20568 19620 20589 19684
rect 20483 19603 20589 19620
rect 35110 19741 35216 19758
rect 35110 19677 35131 19741
rect 35195 19677 35216 19741
rect 35110 19661 35216 19677
rect 35110 19597 35131 19661
rect 35195 19597 35216 19661
rect 35110 19580 35216 19597
rect 35293 19741 35399 19758
rect 35293 19677 35314 19741
rect 35378 19677 35399 19741
rect 35293 19661 35399 19677
rect 35293 19597 35314 19661
rect 35378 19597 35399 19661
rect 35293 19580 35399 19597
rect 35476 19741 35582 19758
rect 35476 19677 35497 19741
rect 35561 19677 35582 19741
rect 35476 19661 35582 19677
rect 35476 19597 35497 19661
rect 35561 19597 35582 19661
rect 35476 19580 35582 19597
rect 50608 19754 50714 19771
rect 50608 19690 50629 19754
rect 50693 19690 50714 19754
rect 50608 19674 50714 19690
rect 50608 19610 50629 19674
rect 50693 19610 50714 19674
rect 50608 19593 50714 19610
rect 50791 19754 50897 19771
rect 50791 19690 50812 19754
rect 50876 19690 50897 19754
rect 50791 19674 50897 19690
rect 50791 19610 50812 19674
rect 50876 19610 50897 19674
rect 50791 19593 50897 19610
rect 50974 19754 51080 19771
rect 50974 19690 50995 19754
rect 51059 19690 51080 19754
rect 50974 19674 51080 19690
rect 50974 19610 50995 19674
rect 51059 19610 51080 19674
rect 50974 19593 51080 19610
rect 18612 17620 18718 17637
rect 18612 17556 18633 17620
rect 18697 17556 18718 17620
rect 18612 17540 18718 17556
rect 18612 17476 18633 17540
rect 18697 17476 18718 17540
rect 18612 17459 18718 17476
rect 18786 17620 18892 17637
rect 18786 17556 18807 17620
rect 18871 17556 18892 17620
rect 18786 17540 18892 17556
rect 18786 17476 18807 17540
rect 18871 17476 18892 17540
rect 18786 17459 18892 17476
rect 18960 17620 19066 17637
rect 18960 17556 18981 17620
rect 19045 17556 19066 17620
rect 18960 17540 19066 17556
rect 18960 17476 18981 17540
rect 19045 17476 19066 17540
rect 18960 17459 19066 17476
rect 33589 17625 33695 17642
rect 33589 17561 33610 17625
rect 33674 17561 33695 17625
rect 33589 17545 33695 17561
rect 33589 17481 33610 17545
rect 33674 17481 33695 17545
rect 33589 17464 33695 17481
rect 33772 17625 33878 17642
rect 33772 17561 33793 17625
rect 33857 17561 33878 17625
rect 33772 17545 33878 17561
rect 33772 17481 33793 17545
rect 33857 17481 33878 17545
rect 33772 17464 33878 17481
rect 33955 17625 34061 17642
rect 33955 17561 33976 17625
rect 34040 17561 34061 17625
rect 33955 17545 34061 17561
rect 33955 17481 33976 17545
rect 34040 17481 34061 17545
rect 33955 17464 34061 17481
rect 49083 17616 49189 17633
rect 49083 17552 49104 17616
rect 49168 17552 49189 17616
rect 49083 17536 49189 17552
rect 49083 17472 49104 17536
rect 49168 17472 49189 17536
rect 49083 17455 49189 17472
rect 49266 17616 49372 17633
rect 49266 17552 49287 17616
rect 49351 17552 49372 17616
rect 49266 17536 49372 17552
rect 49266 17472 49287 17536
rect 49351 17472 49372 17536
rect 49266 17455 49372 17472
rect 49449 17616 49555 17633
rect 49449 17552 49470 17616
rect 49534 17552 49555 17616
rect 49449 17536 49555 17552
rect 49449 17472 49470 17536
rect 49534 17472 49555 17536
rect 49449 17455 49555 17472
rect 30573 15559 30968 15588
rect 30573 15503 30604 15559
rect 30660 15514 30713 15559
rect 30660 15503 30663 15514
rect 30769 15503 30822 15559
rect 30878 15503 30968 15559
rect 30573 15457 30663 15503
rect 30727 15457 30968 15503
rect 30573 15401 30604 15457
rect 30660 15450 30663 15457
rect 30660 15401 30713 15450
rect 30769 15401 30822 15457
rect 30878 15401 30968 15457
rect 30573 15380 30968 15401
rect 18625 14692 18731 14709
rect 18625 14628 18646 14692
rect 18710 14628 18731 14692
rect 18625 14612 18731 14628
rect 18625 14548 18646 14612
rect 18710 14548 18731 14612
rect 18625 14531 18731 14548
rect 18799 14692 18905 14709
rect 18799 14628 18820 14692
rect 18884 14628 18905 14692
rect 18799 14612 18905 14628
rect 18799 14548 18820 14612
rect 18884 14548 18905 14612
rect 18799 14531 18905 14548
rect 18973 14692 19079 14709
rect 18973 14628 18994 14692
rect 19058 14628 19079 14692
rect 18973 14612 19079 14628
rect 18973 14548 18994 14612
rect 19058 14548 19079 14612
rect 18973 14531 19079 14548
rect 31710 14689 31834 14700
rect 31710 14625 31740 14689
rect 31804 14625 31834 14689
rect 31710 14609 31834 14625
rect 31710 14545 31740 14609
rect 31804 14545 31834 14609
rect 31710 14534 31834 14545
rect 31909 14689 32033 14700
rect 31909 14625 31939 14689
rect 32003 14625 32033 14689
rect 31909 14609 32033 14625
rect 31909 14545 31939 14609
rect 32003 14545 32033 14609
rect 31909 14534 32033 14545
rect 33575 14690 33681 14707
rect 33575 14626 33596 14690
rect 33660 14626 33681 14690
rect 33575 14610 33681 14626
rect 33575 14546 33596 14610
rect 33660 14546 33681 14610
rect 33575 14529 33681 14546
rect 33758 14690 33864 14707
rect 33758 14626 33779 14690
rect 33843 14626 33864 14690
rect 33758 14610 33864 14626
rect 33758 14546 33779 14610
rect 33843 14546 33864 14610
rect 33758 14529 33864 14546
rect 33941 14690 34047 14707
rect 33941 14626 33962 14690
rect 34026 14626 34047 14690
rect 33941 14610 34047 14626
rect 33941 14546 33962 14610
rect 34026 14546 34047 14610
rect 33941 14529 34047 14546
rect 49114 14687 49220 14704
rect 49114 14623 49135 14687
rect 49199 14623 49220 14687
rect 49114 14607 49220 14623
rect 49114 14543 49135 14607
rect 49199 14543 49220 14607
rect 49114 14526 49220 14543
rect 49297 14687 49403 14704
rect 49297 14623 49318 14687
rect 49382 14623 49403 14687
rect 49297 14607 49403 14623
rect 49297 14543 49318 14607
rect 49382 14543 49403 14607
rect 49297 14526 49403 14543
rect 49480 14687 49586 14704
rect 49480 14623 49501 14687
rect 49565 14623 49586 14687
rect 49480 14607 49586 14623
rect 49480 14543 49501 14607
rect 49565 14543 49586 14607
rect 49480 14526 49586 14543
rect 20135 12556 20241 12573
rect 20135 12492 20156 12556
rect 20220 12492 20241 12556
rect 20135 12476 20241 12492
rect 20135 12412 20156 12476
rect 20220 12412 20241 12476
rect 20135 12395 20241 12412
rect 20309 12556 20415 12573
rect 20309 12492 20330 12556
rect 20394 12492 20415 12556
rect 20309 12476 20415 12492
rect 20309 12412 20330 12476
rect 20394 12412 20415 12476
rect 20309 12395 20415 12412
rect 20483 12556 20589 12573
rect 20483 12492 20504 12556
rect 20568 12492 20589 12556
rect 20483 12476 20589 12492
rect 20483 12412 20504 12476
rect 20568 12412 20589 12476
rect 20483 12395 20589 12412
rect 35125 12567 35231 12584
rect 35125 12503 35146 12567
rect 35210 12503 35231 12567
rect 35125 12487 35231 12503
rect 35125 12423 35146 12487
rect 35210 12423 35231 12487
rect 35125 12406 35231 12423
rect 35308 12567 35414 12584
rect 35308 12503 35329 12567
rect 35393 12503 35414 12567
rect 35308 12487 35414 12503
rect 35308 12423 35329 12487
rect 35393 12423 35414 12487
rect 35308 12406 35414 12423
rect 35491 12567 35597 12584
rect 35491 12503 35512 12567
rect 35576 12503 35597 12567
rect 35491 12487 35597 12503
rect 35491 12423 35512 12487
rect 35576 12423 35597 12487
rect 35491 12406 35597 12423
rect 50583 12558 50689 12575
rect 50583 12494 50604 12558
rect 50668 12494 50689 12558
rect 50583 12478 50689 12494
rect 50583 12414 50604 12478
rect 50668 12414 50689 12478
rect 50583 12397 50689 12414
rect 50766 12558 50872 12575
rect 50766 12494 50787 12558
rect 50851 12494 50872 12558
rect 50766 12478 50872 12494
rect 50766 12414 50787 12478
rect 50851 12414 50872 12478
rect 50766 12397 50872 12414
rect 50949 12558 51055 12575
rect 50949 12494 50970 12558
rect 51034 12494 51055 12558
rect 50949 12478 51055 12494
rect 50949 12414 50970 12478
rect 51034 12414 51055 12478
rect 50949 12397 51055 12414
rect 30573 10377 30970 10419
rect 30573 10321 30597 10377
rect 30653 10330 30701 10377
rect 30653 10321 30654 10330
rect 30757 10321 30805 10377
rect 30861 10330 30909 10377
rect 30900 10321 30909 10330
rect 30965 10321 30970 10377
rect 30573 10278 30654 10321
rect 30718 10278 30836 10321
rect 30900 10278 30970 10321
rect 30573 10222 30597 10278
rect 30653 10266 30654 10278
rect 30653 10222 30701 10266
rect 30757 10222 30805 10278
rect 30900 10266 30909 10278
rect 30861 10222 30909 10266
rect 30965 10222 30970 10278
rect 30573 10195 30970 10222
rect 31665 9961 32066 9972
rect 31665 9947 31801 9961
rect 31865 9947 31881 9961
rect 31945 9947 32066 9961
rect 31665 9891 31704 9947
rect 31760 9897 31801 9947
rect 31945 9897 31962 9947
rect 31760 9891 31833 9897
rect 31889 9891 31962 9897
rect 32018 9891 32066 9947
rect 31665 9878 32066 9891
rect 7162 9660 7509 9674
rect 61 9644 7509 9660
rect 61 9588 7252 9644
rect 7308 9588 7349 9644
rect 7405 9588 7509 9644
rect 61 9570 7509 9588
rect 7162 9550 7509 9570
rect 30574 9048 30971 9106
rect 30574 8992 30610 9048
rect 30666 9007 30698 9048
rect 30754 8992 30786 9048
rect 30842 9007 30874 9048
rect 30930 8992 30971 9048
rect 30574 8953 30646 8992
rect 30710 8953 30836 8992
rect 30900 8953 30971 8992
rect 30574 8897 30610 8953
rect 30666 8897 30698 8943
rect 30754 8897 30786 8953
rect 30842 8897 30874 8943
rect 30930 8897 30971 8953
rect 30574 8866 30971 8897
rect 3333 7515 3439 7532
rect 3333 7451 3354 7515
rect 3418 7451 3439 7515
rect 3333 7435 3439 7451
rect 3333 7371 3354 7435
rect 3418 7371 3439 7435
rect 3333 7354 3439 7371
rect 3584 7515 3690 7532
rect 3584 7451 3605 7515
rect 3669 7451 3690 7515
rect 3584 7435 3690 7451
rect 3584 7371 3605 7435
rect 3669 7371 3690 7435
rect 3584 7354 3690 7371
rect 3835 7515 3941 7532
rect 3835 7451 3856 7515
rect 3920 7451 3941 7515
rect 3835 7435 3941 7451
rect 3835 7371 3856 7435
rect 3920 7371 3941 7435
rect 3835 7354 3941 7371
rect 20113 7518 20219 7535
rect 20113 7454 20134 7518
rect 20198 7454 20219 7518
rect 20113 7438 20219 7454
rect 20113 7374 20134 7438
rect 20198 7374 20219 7438
rect 20113 7357 20219 7374
rect 20287 7518 20393 7535
rect 20287 7454 20308 7518
rect 20372 7454 20393 7518
rect 20287 7438 20393 7454
rect 20287 7374 20308 7438
rect 20372 7374 20393 7438
rect 20287 7357 20393 7374
rect 20461 7518 20567 7535
rect 20461 7454 20482 7518
rect 20546 7454 20567 7518
rect 20461 7438 20567 7454
rect 20461 7374 20482 7438
rect 20546 7374 20567 7438
rect 20461 7357 20567 7374
rect 35080 7525 35186 7542
rect 35080 7461 35101 7525
rect 35165 7461 35186 7525
rect 35080 7445 35186 7461
rect 35080 7381 35101 7445
rect 35165 7381 35186 7445
rect 35080 7364 35186 7381
rect 35263 7525 35369 7542
rect 35263 7461 35284 7525
rect 35348 7461 35369 7525
rect 35263 7445 35369 7461
rect 35263 7381 35284 7445
rect 35348 7381 35369 7445
rect 35263 7364 35369 7381
rect 35446 7525 35552 7542
rect 35446 7461 35467 7525
rect 35531 7461 35552 7525
rect 35446 7445 35552 7461
rect 35446 7381 35467 7445
rect 35531 7381 35552 7445
rect 35446 7364 35552 7381
rect 50585 7517 50691 7534
rect 50585 7453 50606 7517
rect 50670 7453 50691 7517
rect 50585 7437 50691 7453
rect 50585 7373 50606 7437
rect 50670 7373 50691 7437
rect 50585 7356 50691 7373
rect 50768 7517 50874 7534
rect 50768 7453 50789 7517
rect 50853 7453 50874 7517
rect 50768 7437 50874 7453
rect 50768 7373 50789 7437
rect 50853 7373 50874 7437
rect 50768 7356 50874 7373
rect 50951 7517 51057 7534
rect 50951 7453 50972 7517
rect 51036 7453 51057 7517
rect 50951 7437 51057 7453
rect 50951 7373 50972 7437
rect 51036 7373 51057 7437
rect 50951 7356 51057 7373
rect 2108 5386 2214 5403
rect 2108 5322 2129 5386
rect 2193 5322 2214 5386
rect 2108 5306 2214 5322
rect 2108 5242 2129 5306
rect 2193 5242 2214 5306
rect 2108 5225 2214 5242
rect 2284 5386 2390 5403
rect 2284 5322 2305 5386
rect 2369 5322 2390 5386
rect 2284 5306 2390 5322
rect 2284 5242 2305 5306
rect 2369 5242 2390 5306
rect 2284 5225 2390 5242
rect 2460 5386 2566 5403
rect 2460 5322 2481 5386
rect 2545 5322 2566 5386
rect 2460 5306 2566 5322
rect 2460 5242 2481 5306
rect 2545 5242 2566 5306
rect 2460 5225 2566 5242
rect 18611 5392 18717 5409
rect 18611 5328 18632 5392
rect 18696 5328 18717 5392
rect 18611 5312 18717 5328
rect 18611 5248 18632 5312
rect 18696 5248 18717 5312
rect 18611 5231 18717 5248
rect 18785 5392 18891 5409
rect 18785 5328 18806 5392
rect 18870 5328 18891 5392
rect 18785 5312 18891 5328
rect 18785 5248 18806 5312
rect 18870 5248 18891 5312
rect 18785 5231 18891 5248
rect 18959 5392 19065 5409
rect 18959 5328 18980 5392
rect 19044 5328 19065 5392
rect 18959 5312 19065 5328
rect 18959 5248 18980 5312
rect 19044 5248 19065 5312
rect 18959 5231 19065 5248
rect 33587 5393 33693 5410
rect 33587 5329 33608 5393
rect 33672 5329 33693 5393
rect 33587 5313 33693 5329
rect 33587 5249 33608 5313
rect 33672 5249 33693 5313
rect 33587 5232 33693 5249
rect 33770 5393 33876 5410
rect 33770 5329 33791 5393
rect 33855 5329 33876 5393
rect 33770 5313 33876 5329
rect 33770 5249 33791 5313
rect 33855 5249 33876 5313
rect 33770 5232 33876 5249
rect 33953 5393 34059 5410
rect 33953 5329 33974 5393
rect 34038 5329 34059 5393
rect 33953 5313 34059 5329
rect 33953 5249 33974 5313
rect 34038 5249 34059 5313
rect 33953 5232 34059 5249
rect 49082 5389 49188 5406
rect 49082 5325 49103 5389
rect 49167 5325 49188 5389
rect 49082 5309 49188 5325
rect 49082 5245 49103 5309
rect 49167 5245 49188 5309
rect 49082 5228 49188 5245
rect 49265 5389 49371 5406
rect 49265 5325 49286 5389
rect 49350 5325 49371 5389
rect 49265 5309 49371 5325
rect 49265 5245 49286 5309
rect 49350 5245 49371 5309
rect 49265 5228 49371 5245
rect 49448 5389 49554 5406
rect 49448 5325 49469 5389
rect 49533 5325 49554 5389
rect 49448 5309 49554 5325
rect 49448 5245 49469 5309
rect 49533 5245 49554 5309
rect 49448 5228 49554 5245
rect 30574 3324 30971 3357
rect 30574 3268 30615 3324
rect 30671 3278 30707 3324
rect 30763 3268 30799 3324
rect 30855 3279 30891 3324
rect 30947 3268 30971 3324
rect 30574 3233 30658 3268
rect 30722 3233 30832 3268
rect 30896 3233 30971 3268
rect 30574 3177 30615 3233
rect 30671 3177 30707 3214
rect 30763 3177 30799 3233
rect 30855 3177 30891 3215
rect 30947 3177 30971 3233
rect 30574 3151 30971 3177
rect 2104 2453 2210 2470
rect 2104 2389 2125 2453
rect 2189 2389 2210 2453
rect 2104 2373 2210 2389
rect 2104 2309 2125 2373
rect 2189 2309 2210 2373
rect 2104 2292 2210 2309
rect 2280 2453 2386 2470
rect 2280 2389 2301 2453
rect 2365 2389 2386 2453
rect 2280 2373 2386 2389
rect 2280 2309 2301 2373
rect 2365 2309 2386 2373
rect 2280 2292 2386 2309
rect 2456 2453 2562 2470
rect 2456 2389 2477 2453
rect 2541 2389 2562 2453
rect 2456 2373 2562 2389
rect 2456 2309 2477 2373
rect 2541 2309 2562 2373
rect 2456 2292 2562 2309
rect 18608 2456 18714 2473
rect 18608 2392 18629 2456
rect 18693 2392 18714 2456
rect 18608 2376 18714 2392
rect 18608 2312 18629 2376
rect 18693 2312 18714 2376
rect 18608 2295 18714 2312
rect 18782 2456 18888 2473
rect 18782 2392 18803 2456
rect 18867 2392 18888 2456
rect 18782 2376 18888 2392
rect 18782 2312 18803 2376
rect 18867 2312 18888 2376
rect 18782 2295 18888 2312
rect 18956 2456 19062 2473
rect 18956 2392 18977 2456
rect 19041 2392 19062 2456
rect 18956 2376 19062 2392
rect 18956 2312 18977 2376
rect 19041 2312 19062 2376
rect 18956 2295 19062 2312
rect 33599 2452 33705 2469
rect 33599 2388 33620 2452
rect 33684 2388 33705 2452
rect 33599 2372 33705 2388
rect 33599 2308 33620 2372
rect 33684 2308 33705 2372
rect 33599 2291 33705 2308
rect 33782 2452 33888 2469
rect 33782 2388 33803 2452
rect 33867 2388 33888 2452
rect 33782 2372 33888 2388
rect 33782 2308 33803 2372
rect 33867 2308 33888 2372
rect 33782 2291 33888 2308
rect 33965 2452 34071 2469
rect 33965 2388 33986 2452
rect 34050 2388 34071 2452
rect 33965 2372 34071 2388
rect 33965 2308 33986 2372
rect 34050 2308 34071 2372
rect 33965 2291 34071 2308
rect 49090 2456 49196 2473
rect 49090 2392 49111 2456
rect 49175 2392 49196 2456
rect 49090 2376 49196 2392
rect 49090 2312 49111 2376
rect 49175 2312 49196 2376
rect 49090 2295 49196 2312
rect 49273 2456 49379 2473
rect 49273 2392 49294 2456
rect 49358 2392 49379 2456
rect 49273 2376 49379 2392
rect 49273 2312 49294 2376
rect 49358 2312 49379 2376
rect 49273 2295 49379 2312
rect 49456 2456 49562 2473
rect 49456 2392 49477 2456
rect 49541 2392 49562 2456
rect 49456 2376 49562 2392
rect 49456 2312 49477 2376
rect 49541 2312 49562 2376
rect 49456 2295 49562 2312
rect 3367 331 3473 348
rect 3367 267 3388 331
rect 3452 267 3473 331
rect 3367 251 3473 267
rect 3367 187 3388 251
rect 3452 187 3473 251
rect 3367 170 3473 187
rect 3618 331 3724 348
rect 3618 267 3639 331
rect 3703 267 3724 331
rect 3618 251 3724 267
rect 3618 187 3639 251
rect 3703 187 3724 251
rect 3618 170 3724 187
rect 3869 331 3975 348
rect 3869 267 3890 331
rect 3954 267 3975 331
rect 3869 251 3975 267
rect 3869 187 3890 251
rect 3954 187 3975 251
rect 3869 170 3975 187
rect 20117 334 20223 351
rect 20117 270 20138 334
rect 20202 270 20223 334
rect 20117 254 20223 270
rect 20117 190 20138 254
rect 20202 190 20223 254
rect 20117 173 20223 190
rect 20291 334 20397 351
rect 20291 270 20312 334
rect 20376 270 20397 334
rect 20291 254 20397 270
rect 20291 190 20312 254
rect 20376 190 20397 254
rect 20291 173 20397 190
rect 20465 334 20571 351
rect 20465 270 20486 334
rect 20550 270 20571 334
rect 20465 254 20571 270
rect 20465 190 20486 254
rect 20550 190 20571 254
rect 20465 173 20571 190
rect 35126 345 35232 362
rect 35126 281 35147 345
rect 35211 281 35232 345
rect 35126 265 35232 281
rect 35126 201 35147 265
rect 35211 201 35232 265
rect 35126 184 35232 201
rect 35309 345 35415 362
rect 35309 281 35330 345
rect 35394 281 35415 345
rect 35309 265 35415 281
rect 35309 201 35330 265
rect 35394 201 35415 265
rect 35309 184 35415 201
rect 35492 345 35598 362
rect 35492 281 35513 345
rect 35577 281 35598 345
rect 35492 265 35598 281
rect 35492 201 35513 265
rect 35577 201 35598 265
rect 35492 184 35598 201
rect 50626 337 50732 354
rect 50626 273 50647 337
rect 50711 273 50732 337
rect 50626 257 50732 273
rect 50626 193 50647 257
rect 50711 193 50732 257
rect 50626 176 50732 193
rect 50809 337 50915 354
rect 50809 273 50830 337
rect 50894 273 50915 337
rect 50809 257 50915 273
rect 50809 193 50830 257
rect 50894 193 50915 257
rect 50809 176 50915 193
rect 50992 337 51098 354
rect 50992 273 51013 337
rect 51077 273 51098 337
rect 50992 257 51098 273
rect 50992 193 51013 257
rect 51077 193 51098 257
rect 50992 176 51098 193
<< via3 >>
rect 20156 19700 20220 19764
rect 20156 19620 20220 19684
rect 20330 19700 20394 19764
rect 20330 19620 20394 19684
rect 20504 19700 20568 19764
rect 20504 19620 20568 19684
rect 35131 19677 35195 19741
rect 35131 19597 35195 19661
rect 35314 19677 35378 19741
rect 35314 19597 35378 19661
rect 35497 19677 35561 19741
rect 35497 19597 35561 19661
rect 50629 19690 50693 19754
rect 50629 19610 50693 19674
rect 50812 19690 50876 19754
rect 50812 19610 50876 19674
rect 50995 19690 51059 19754
rect 50995 19610 51059 19674
rect 18633 17556 18697 17620
rect 18633 17476 18697 17540
rect 18807 17556 18871 17620
rect 18807 17476 18871 17540
rect 18981 17556 19045 17620
rect 18981 17476 19045 17540
rect 33610 17561 33674 17625
rect 33610 17481 33674 17545
rect 33793 17561 33857 17625
rect 33793 17481 33857 17545
rect 33976 17561 34040 17625
rect 33976 17481 34040 17545
rect 49104 17552 49168 17616
rect 49104 17472 49168 17536
rect 49287 17552 49351 17616
rect 49287 17472 49351 17536
rect 49470 17552 49534 17616
rect 49470 17472 49534 17536
rect 30663 15503 30713 15514
rect 30713 15503 30727 15514
rect 30663 15457 30727 15503
rect 30663 15450 30713 15457
rect 30713 15450 30727 15457
rect 18646 14628 18710 14692
rect 18646 14548 18710 14612
rect 18820 14628 18884 14692
rect 18820 14548 18884 14612
rect 18994 14628 19058 14692
rect 18994 14548 19058 14612
rect 31740 14625 31804 14689
rect 31740 14545 31804 14609
rect 31939 14625 32003 14689
rect 31939 14545 32003 14609
rect 33596 14626 33660 14690
rect 33596 14546 33660 14610
rect 33779 14626 33843 14690
rect 33779 14546 33843 14610
rect 33962 14626 34026 14690
rect 33962 14546 34026 14610
rect 49135 14623 49199 14687
rect 49135 14543 49199 14607
rect 49318 14623 49382 14687
rect 49318 14543 49382 14607
rect 49501 14623 49565 14687
rect 49501 14543 49565 14607
rect 20156 12492 20220 12556
rect 20156 12412 20220 12476
rect 20330 12492 20394 12556
rect 20330 12412 20394 12476
rect 20504 12492 20568 12556
rect 20504 12412 20568 12476
rect 35146 12503 35210 12567
rect 35146 12423 35210 12487
rect 35329 12503 35393 12567
rect 35329 12423 35393 12487
rect 35512 12503 35576 12567
rect 35512 12423 35576 12487
rect 50604 12494 50668 12558
rect 50604 12414 50668 12478
rect 50787 12494 50851 12558
rect 50787 12414 50851 12478
rect 50970 12494 51034 12558
rect 50970 12414 51034 12478
rect 30654 10321 30701 10330
rect 30701 10321 30718 10330
rect 30836 10321 30861 10330
rect 30861 10321 30900 10330
rect 30654 10278 30718 10321
rect 30836 10278 30900 10321
rect 30654 10266 30701 10278
rect 30701 10266 30718 10278
rect 30836 10266 30861 10278
rect 30861 10266 30900 10278
rect 31801 9947 31865 9961
rect 31881 9947 31945 9961
rect 31801 9897 31833 9947
rect 31833 9897 31865 9947
rect 31881 9897 31889 9947
rect 31889 9897 31945 9947
rect 30646 8992 30666 9007
rect 30666 8992 30698 9007
rect 30698 8992 30710 9007
rect 30836 8992 30842 9007
rect 30842 8992 30874 9007
rect 30874 8992 30900 9007
rect 30646 8953 30710 8992
rect 30836 8953 30900 8992
rect 30646 8943 30666 8953
rect 30666 8943 30698 8953
rect 30698 8943 30710 8953
rect 30836 8943 30842 8953
rect 30842 8943 30874 8953
rect 30874 8943 30900 8953
rect 3354 7451 3418 7515
rect 3354 7371 3418 7435
rect 3605 7451 3669 7515
rect 3605 7371 3669 7435
rect 3856 7451 3920 7515
rect 3856 7371 3920 7435
rect 20134 7454 20198 7518
rect 20134 7374 20198 7438
rect 20308 7454 20372 7518
rect 20308 7374 20372 7438
rect 20482 7454 20546 7518
rect 20482 7374 20546 7438
rect 35101 7461 35165 7525
rect 35101 7381 35165 7445
rect 35284 7461 35348 7525
rect 35284 7381 35348 7445
rect 35467 7461 35531 7525
rect 35467 7381 35531 7445
rect 50606 7453 50670 7517
rect 50606 7373 50670 7437
rect 50789 7453 50853 7517
rect 50789 7373 50853 7437
rect 50972 7453 51036 7517
rect 50972 7373 51036 7437
rect 2129 5322 2193 5386
rect 2129 5242 2193 5306
rect 2305 5322 2369 5386
rect 2305 5242 2369 5306
rect 2481 5322 2545 5386
rect 2481 5242 2545 5306
rect 18632 5328 18696 5392
rect 18632 5248 18696 5312
rect 18806 5328 18870 5392
rect 18806 5248 18870 5312
rect 18980 5328 19044 5392
rect 18980 5248 19044 5312
rect 33608 5329 33672 5393
rect 33608 5249 33672 5313
rect 33791 5329 33855 5393
rect 33791 5249 33855 5313
rect 33974 5329 34038 5393
rect 33974 5249 34038 5313
rect 49103 5325 49167 5389
rect 49103 5245 49167 5309
rect 49286 5325 49350 5389
rect 49286 5245 49350 5309
rect 49469 5325 49533 5389
rect 49469 5245 49533 5309
rect 30658 3268 30671 3278
rect 30671 3268 30707 3278
rect 30707 3268 30722 3278
rect 30832 3268 30855 3279
rect 30855 3268 30891 3279
rect 30891 3268 30896 3279
rect 30658 3233 30722 3268
rect 30832 3233 30896 3268
rect 30658 3214 30671 3233
rect 30671 3214 30707 3233
rect 30707 3214 30722 3233
rect 30832 3215 30855 3233
rect 30855 3215 30891 3233
rect 30891 3215 30896 3233
rect 2125 2389 2189 2453
rect 2125 2309 2189 2373
rect 2301 2389 2365 2453
rect 2301 2309 2365 2373
rect 2477 2389 2541 2453
rect 2477 2309 2541 2373
rect 18629 2392 18693 2456
rect 18629 2312 18693 2376
rect 18803 2392 18867 2456
rect 18803 2312 18867 2376
rect 18977 2392 19041 2456
rect 18977 2312 19041 2376
rect 33620 2388 33684 2452
rect 33620 2308 33684 2372
rect 33803 2388 33867 2452
rect 33803 2308 33867 2372
rect 33986 2388 34050 2452
rect 33986 2308 34050 2372
rect 49111 2392 49175 2456
rect 49111 2312 49175 2376
rect 49294 2392 49358 2456
rect 49294 2312 49358 2376
rect 49477 2392 49541 2456
rect 49477 2312 49541 2376
rect 3388 267 3452 331
rect 3388 187 3452 251
rect 3639 267 3703 331
rect 3639 187 3703 251
rect 3890 267 3954 331
rect 3890 187 3954 251
rect 20138 270 20202 334
rect 20138 190 20202 254
rect 20312 270 20376 334
rect 20312 190 20376 254
rect 20486 270 20550 334
rect 20486 190 20550 254
rect 35147 281 35211 345
rect 35147 201 35211 265
rect 35330 281 35394 345
rect 35330 201 35394 265
rect 35513 281 35577 345
rect 35513 201 35577 265
rect 50647 273 50711 337
rect 50647 193 50711 257
rect 50830 273 50894 337
rect 50830 193 50894 257
rect 51013 273 51077 337
rect 51013 193 51077 257
<< metal4 >>
rect 2024 5386 2642 20087
rect 2024 5322 2129 5386
rect 2193 5322 2305 5386
rect 2369 5322 2481 5386
rect 2545 5322 2642 5386
rect 2024 5306 2642 5322
rect 2024 5242 2129 5306
rect 2193 5242 2305 5306
rect 2369 5242 2481 5306
rect 2545 5242 2642 5306
rect 2024 2453 2642 5242
rect 2024 2389 2125 2453
rect 2189 2389 2301 2453
rect 2365 2389 2477 2453
rect 2541 2389 2642 2453
rect 2024 2373 2642 2389
rect 2024 2309 2125 2373
rect 2189 2309 2301 2373
rect 2365 2309 2477 2373
rect 2541 2309 2642 2373
rect 2024 38 2642 2309
rect 3257 7515 4041 20087
rect 3257 7451 3354 7515
rect 3418 7451 3605 7515
rect 3669 7451 3856 7515
rect 3920 7451 4041 7515
rect 3257 7435 4041 7451
rect 3257 7371 3354 7435
rect 3418 7371 3605 7435
rect 3669 7371 3856 7435
rect 3920 7371 4041 7435
rect 3257 331 4041 7371
rect 3257 267 3388 331
rect 3452 267 3639 331
rect 3703 267 3890 331
rect 3954 267 4041 331
rect 3257 251 4041 267
rect 3257 187 3388 251
rect 3452 187 3639 251
rect 3703 187 3890 251
rect 3954 187 4041 251
rect 3257 74 4041 187
rect 18524 17620 19142 20087
rect 18524 17556 18633 17620
rect 18697 17556 18807 17620
rect 18871 17556 18981 17620
rect 19045 17556 19142 17620
rect 18524 17540 19142 17556
rect 18524 17476 18633 17540
rect 18697 17476 18807 17540
rect 18871 17476 18981 17540
rect 19045 17476 19142 17540
rect 18524 14692 19142 17476
rect 18524 14628 18646 14692
rect 18710 14628 18820 14692
rect 18884 14628 18994 14692
rect 19058 14628 19142 14692
rect 18524 14612 19142 14628
rect 18524 14548 18646 14612
rect 18710 14548 18820 14612
rect 18884 14548 18994 14612
rect 19058 14548 19142 14612
rect 18524 5392 19142 14548
rect 18524 5328 18632 5392
rect 18696 5328 18806 5392
rect 18870 5328 18980 5392
rect 19044 5328 19142 5392
rect 18524 5312 19142 5328
rect 18524 5248 18632 5312
rect 18696 5248 18806 5312
rect 18870 5248 18980 5312
rect 19044 5248 19142 5312
rect 18524 2456 19142 5248
rect 18524 2392 18629 2456
rect 18693 2392 18803 2456
rect 18867 2392 18977 2456
rect 19041 2392 19142 2456
rect 18524 2376 19142 2392
rect 18524 2312 18629 2376
rect 18693 2312 18803 2376
rect 18867 2312 18977 2376
rect 19041 2312 19142 2376
rect 18524 38 19142 2312
rect 20024 19764 20642 20087
rect 20024 19700 20156 19764
rect 20220 19700 20330 19764
rect 20394 19700 20504 19764
rect 20568 19700 20642 19764
rect 20024 19684 20642 19700
rect 20024 19620 20156 19684
rect 20220 19620 20330 19684
rect 20394 19620 20504 19684
rect 20568 19620 20642 19684
rect 20024 12556 20642 19620
rect 33524 17625 34142 20087
rect 33524 17561 33610 17625
rect 33674 17561 33793 17625
rect 33857 17561 33976 17625
rect 34040 17561 34142 17625
rect 33524 17545 34142 17561
rect 33524 17481 33610 17545
rect 33674 17481 33793 17545
rect 33857 17481 33976 17545
rect 34040 17481 34142 17545
rect 20024 12492 20156 12556
rect 20220 12492 20330 12556
rect 20394 12492 20504 12556
rect 20568 12492 20642 12556
rect 20024 12476 20642 12492
rect 20024 12412 20156 12476
rect 20220 12412 20330 12476
rect 20394 12412 20504 12476
rect 20568 12412 20642 12476
rect 20024 7518 20642 12412
rect 30573 15514 30970 15648
rect 30573 15450 30663 15514
rect 30727 15450 30970 15514
rect 30573 10856 30970 15450
rect 30572 10495 30970 10856
rect 30573 10330 30970 10495
rect 30573 10266 30654 10330
rect 30718 10266 30836 10330
rect 30900 10266 30970 10330
rect 30573 10195 30970 10266
rect 31658 14689 32062 14819
rect 31658 14625 31740 14689
rect 31804 14625 31939 14689
rect 32003 14625 32062 14689
rect 31658 14609 32062 14625
rect 31658 14545 31740 14609
rect 31804 14545 31939 14609
rect 32003 14545 32062 14609
rect 31658 9989 32062 14545
rect 33524 14690 34142 17481
rect 33524 14626 33596 14690
rect 33660 14626 33779 14690
rect 33843 14626 33962 14690
rect 34026 14626 34142 14690
rect 33524 14610 34142 14626
rect 33524 14546 33596 14610
rect 33660 14546 33779 14610
rect 33843 14546 33962 14610
rect 34026 14546 34142 14610
rect 31658 9967 32066 9989
rect 31665 9961 32066 9967
rect 31665 9897 31801 9961
rect 31865 9897 31881 9961
rect 31945 9897 32066 9961
rect 31665 9878 32066 9897
rect 20024 7454 20134 7518
rect 20198 7454 20308 7518
rect 20372 7454 20482 7518
rect 20546 7454 20642 7518
rect 20024 7438 20642 7454
rect 20024 7374 20134 7438
rect 20198 7374 20308 7438
rect 20372 7374 20482 7438
rect 20546 7374 20642 7438
rect 20024 334 20642 7374
rect 30575 9007 30971 9105
rect 30575 8943 30646 9007
rect 30710 8943 30836 9007
rect 30900 8943 30971 9007
rect 30575 3279 30971 8943
rect 30575 3278 30832 3279
rect 30575 3214 30658 3278
rect 30722 3215 30832 3278
rect 30896 3215 30971 3279
rect 30722 3214 30971 3215
rect 30575 3089 30971 3214
rect 33524 5393 34142 14546
rect 33524 5329 33608 5393
rect 33672 5329 33791 5393
rect 33855 5329 33974 5393
rect 34038 5329 34142 5393
rect 33524 5313 34142 5329
rect 33524 5249 33608 5313
rect 33672 5249 33791 5313
rect 33855 5249 33974 5313
rect 34038 5249 34142 5313
rect 20024 270 20138 334
rect 20202 270 20312 334
rect 20376 270 20486 334
rect 20550 270 20642 334
rect 20024 254 20642 270
rect 20024 190 20138 254
rect 20202 190 20312 254
rect 20376 190 20486 254
rect 20550 190 20642 254
rect 20024 38 20642 190
rect 33524 2452 34142 5249
rect 33524 2388 33620 2452
rect 33684 2388 33803 2452
rect 33867 2388 33986 2452
rect 34050 2388 34142 2452
rect 33524 2372 34142 2388
rect 33524 2308 33620 2372
rect 33684 2308 33803 2372
rect 33867 2308 33986 2372
rect 34050 2308 34142 2372
rect 33524 38 34142 2308
rect 35024 19741 35642 20087
rect 35024 19677 35131 19741
rect 35195 19677 35314 19741
rect 35378 19677 35497 19741
rect 35561 19677 35642 19741
rect 35024 19661 35642 19677
rect 35024 19597 35131 19661
rect 35195 19597 35314 19661
rect 35378 19597 35497 19661
rect 35561 19597 35642 19661
rect 35024 12567 35642 19597
rect 35024 12503 35146 12567
rect 35210 12503 35329 12567
rect 35393 12503 35512 12567
rect 35576 12503 35642 12567
rect 35024 12487 35642 12503
rect 35024 12423 35146 12487
rect 35210 12423 35329 12487
rect 35393 12423 35512 12487
rect 35576 12423 35642 12487
rect 35024 7525 35642 12423
rect 35024 7461 35101 7525
rect 35165 7461 35284 7525
rect 35348 7461 35467 7525
rect 35531 7461 35642 7525
rect 35024 7445 35642 7461
rect 35024 7381 35101 7445
rect 35165 7381 35284 7445
rect 35348 7381 35467 7445
rect 35531 7381 35642 7445
rect 35024 345 35642 7381
rect 35024 281 35147 345
rect 35211 281 35330 345
rect 35394 281 35513 345
rect 35577 281 35642 345
rect 35024 265 35642 281
rect 35024 201 35147 265
rect 35211 201 35330 265
rect 35394 201 35513 265
rect 35577 201 35642 265
rect 35024 38 35642 201
rect 49024 17616 49642 20087
rect 49024 17552 49104 17616
rect 49168 17552 49287 17616
rect 49351 17552 49470 17616
rect 49534 17552 49642 17616
rect 49024 17536 49642 17552
rect 49024 17472 49104 17536
rect 49168 17472 49287 17536
rect 49351 17472 49470 17536
rect 49534 17472 49642 17536
rect 49024 14687 49642 17472
rect 49024 14623 49135 14687
rect 49199 14623 49318 14687
rect 49382 14623 49501 14687
rect 49565 14623 49642 14687
rect 49024 14607 49642 14623
rect 49024 14543 49135 14607
rect 49199 14543 49318 14607
rect 49382 14543 49501 14607
rect 49565 14543 49642 14607
rect 49024 5389 49642 14543
rect 49024 5325 49103 5389
rect 49167 5325 49286 5389
rect 49350 5325 49469 5389
rect 49533 5325 49642 5389
rect 49024 5309 49642 5325
rect 49024 5245 49103 5309
rect 49167 5245 49286 5309
rect 49350 5245 49469 5309
rect 49533 5245 49642 5309
rect 49024 2456 49642 5245
rect 49024 2392 49111 2456
rect 49175 2392 49294 2456
rect 49358 2392 49477 2456
rect 49541 2392 49642 2456
rect 49024 2376 49642 2392
rect 49024 2312 49111 2376
rect 49175 2312 49294 2376
rect 49358 2312 49477 2376
rect 49541 2312 49642 2376
rect 49024 38 49642 2312
rect 50524 19754 51142 20087
rect 50524 19690 50629 19754
rect 50693 19690 50812 19754
rect 50876 19690 50995 19754
rect 51059 19690 51142 19754
rect 50524 19674 51142 19690
rect 50524 19610 50629 19674
rect 50693 19610 50812 19674
rect 50876 19610 50995 19674
rect 51059 19610 51142 19674
rect 50524 12558 51142 19610
rect 50524 12494 50604 12558
rect 50668 12494 50787 12558
rect 50851 12494 50970 12558
rect 51034 12494 51142 12558
rect 50524 12478 51142 12494
rect 50524 12414 50604 12478
rect 50668 12414 50787 12478
rect 50851 12414 50970 12478
rect 51034 12414 51142 12478
rect 50524 7517 51142 12414
rect 50524 7453 50606 7517
rect 50670 7453 50789 7517
rect 50853 7453 50972 7517
rect 51036 7453 51142 7517
rect 50524 7437 51142 7453
rect 50524 7373 50606 7437
rect 50670 7373 50789 7437
rect 50853 7373 50972 7437
rect 51036 7373 51142 7437
rect 50524 337 51142 7373
rect 50524 273 50647 337
rect 50711 273 50830 337
rect 50894 273 51013 337
rect 51077 273 51142 337
rect 50524 257 51142 273
rect 50524 193 50647 257
rect 50711 193 50830 257
rect 50894 193 51013 257
rect 51077 193 51142 257
rect 50524 38 51142 193
use BR128half  BR128half_0
timestamp 1483428465
transform 1 0 790 0 1 12369
box -430 -58 60604 7443
use BR128half  BR128half_1
timestamp 1483428465
transform -1 0 61001 0 1 138
box -430 -58 60604 7443
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0
timestamp 1483428465
transform 1 0 27641 0 1 9381
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0
timestamp 1483428465
transform 1 0 28177 0 1 9381
box -38 -48 866 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0
timestamp 1483428465
transform 1 0 29081 0 1 9381
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1483428465
transform 1 0 30997 0 1 9381
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1483428465
transform 1 0 30740 0 1 9381
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1483428465
transform 1 0 28009 0 1 9381
box -38 -48 130 592
<< labels >>
flabel metal1 s 61150 13149 61394 13227 1 FreeSans 1000 0 0 0 OUT
port 1 nsew
flabel metal1 s 61176 10030 61648 10091 1 FreeSans 1000 0 0 0 C[127]
port 2 nsew
flabel metal1 s 61176 10172 61648 10233 1 FreeSans 1000 0 0 0 C[126]
port 3 nsew
flabel metal1 s 61176 10314 61648 10375 1 FreeSans 1000 0 0 0 C[125]
port 4 nsew
flabel metal1 s 61176 10456 61648 10517 1 FreeSans 1000 0 0 0 C[124]
port 5 nsew
flabel metal1 s 61176 10598 61648 10659 1 FreeSans 1000 0 0 0 C[123]
port 6 nsew
flabel metal1 s 61176 10740 61648 10801 1 FreeSans 1000 0 0 0 C[122]
port 7 nsew
flabel metal1 s 61176 10882 61648 10943 1 FreeSans 1000 0 0 0 C[121]
port 8 nsew
flabel metal1 s 61176 11024 61648 11085 1 FreeSans 1000 0 0 0 C[120]
port 9 nsew
flabel metal1 s 61176 11166 61648 11227 1 FreeSans 1000 0 0 0 C[119]
port 10 nsew
flabel metal1 s 61176 11308 61648 11369 1 FreeSans 1000 0 0 0 C[118]
port 11 nsew
flabel metal1 s 61176 11450 61648 11511 1 FreeSans 1000 0 0 0 C[117]
port 12 nsew
flabel metal1 s 61176 11592 61648 11653 1 FreeSans 1000 0 0 0 C[116]
port 13 nsew
flabel metal1 s 61176 11734 61648 11795 1 FreeSans 1000 0 0 0 C[115]
port 14 nsew
flabel metal1 s 61176 11876 61648 11937 1 FreeSans 1000 0 0 0 C[114]
port 15 nsew
flabel metal1 s 61176 12018 61648 12079 1 FreeSans 1000 0 0 0 C[113]
port 16 nsew
flabel metal1 s 61176 12160 61648 12221 1 FreeSans 1000 0 0 0 C[112]
port 17 nsew
flabel metal1 s 61176 9888 61648 9949 1 FreeSans 1000 0 0 0 C[63]
port 18 nsew
flabel metal1 s 61176 9746 61648 9807 1 FreeSans 1000 0 0 0 C[62]
port 19 nsew
flabel metal1 s 61176 9604 61648 9665 1 FreeSans 1000 0 0 0 C[61]
port 20 nsew
flabel metal1 s 61176 9462 61648 9523 1 FreeSans 1000 0 0 0 C[60]
port 21 nsew
flabel metal1 s 61176 9320 61648 9381 1 FreeSans 1000 0 0 0 C[59]
port 22 nsew
flabel metal1 s 61176 9178 61648 9239 1 FreeSans 1000 0 0 0 C[58]
port 23 nsew
flabel metal1 s 61176 9036 61648 9097 1 FreeSans 1000 0 0 0 C[57]
port 24 nsew
flabel metal1 s 61176 8894 61648 8955 1 FreeSans 1000 0 0 0 C[56]
port 25 nsew
flabel metal1 s 61176 8752 61648 8813 1 FreeSans 1000 0 0 0 C[55]
port 26 nsew
flabel metal1 s 61176 8610 61648 8671 1 FreeSans 1000 0 0 0 C[54]
port 27 nsew
flabel metal1 s 61176 8468 61648 8529 1 FreeSans 1000 0 0 0 C[53]
port 28 nsew
flabel metal1 s 61176 8326 61648 8387 1 FreeSans 1000 0 0 0 C[52]
port 29 nsew
flabel metal1 s 61176 8184 61648 8245 1 FreeSans 1000 0 0 0 C[51]
port 30 nsew
flabel metal1 s 61176 8042 61648 8103 1 FreeSans 1000 0 0 0 C[50]
port 31 nsew
flabel metal1 s 61176 7900 61648 7961 1 FreeSans 1000 0 0 0 C[49]
port 32 nsew
flabel metal1 s 61176 7758 61648 7819 1 FreeSans 1000 0 0 0 C[48]
port 33 nsew
flabel metal3 s 61 9570 307 9660 1 FreeSans 500 0 0 0 RESET
port 34 nsew
flabel metal4 s 2024 38 2642 20087 1 FreeSans 2000 0 0 0 VDD
port 35 nsew
flabel metal4 s 18524 38 19142 20087 1 FreeSans 2000 0 0 0 VDD
port 35 nsew
flabel metal4 s 33524 38 34142 20087 1 FreeSans 2000 0 0 0 VDD
port 35 nsew
flabel metal4 s 49024 38 49642 20087 1 FreeSans 2000 0 0 0 VDD
port 35 nsew
flabel metal4 s 3257 74 4041 20087 1 FreeSans 2000 0 0 0 VSS
port 36 nsew
flabel metal4 s 20024 38 20642 20087 1 FreeSans 2000 0 0 0 VSS
port 36 nsew
flabel metal4 s 35024 38 35642 20087 1 FreeSans 2000 0 0 0 VSS
port 36 nsew
flabel metal4 s 50524 38 51142 20087 1 FreeSans 2000 0 0 0 VSS
port 36 nsew
flabel metal1 s 0 12163 460 12224 1 FreeSans 1500 0 0 0 C[111]
port 37 nsew
flabel metal1 s 0 12021 460 12082 1 FreeSans 1500 0 0 0 C[110]
port 38 nsew
flabel metal1 s 0 11879 460 11940 1 FreeSans 1500 0 0 0 C[109]
port 39 nsew
flabel metal1 s 0 11737 460 11798 1 FreeSans 1500 0 0 0 C[108]
port 40 nsew
flabel metal1 s 0 11595 460 11656 1 FreeSans 1500 0 0 0 C[107]
port 41 nsew
flabel metal1 s 0 11453 460 11514 1 FreeSans 1500 0 0 0 C[106]
port 42 nsew
flabel metal1 s 0 11311 460 11372 1 FreeSans 1500 0 0 0 C[105]
port 43 nsew
flabel metal1 s 0 11169 460 11230 1 FreeSans 1500 0 0 0 C[104]
port 44 nsew
flabel metal1 s 0 11027 460 11088 1 FreeSans 1500 0 0 0 C[103]
port 45 nsew
flabel metal1 s 0 10885 460 10946 1 FreeSans 1500 0 0 0 C[102]
port 46 nsew
flabel metal1 s 0 10743 460 10804 1 FreeSans 1500 0 0 0 C[101]
port 47 nsew
flabel metal1 s 0 10601 460 10662 1 FreeSans 1500 0 0 0 C[100]
port 48 nsew
flabel metal1 s 0 10459 460 10520 1 FreeSans 1500 0 0 0 C[99]
port 49 nsew
flabel metal1 s 0 10317 460 10378 1 FreeSans 1500 0 0 0 C[98]
port 50 nsew
flabel metal1 s 0 10175 460 10236 1 FreeSans 1500 0 0 0 C[97]
port 51 nsew
flabel metal1 s 0 10033 460 10094 1 FreeSans 1500 0 0 0 C[96]
port 52 nsew
flabel metal1 s 0 9891 460 9952 1 FreeSans 1500 0 0 0 C[32]
port 53 nsew
flabel metal1 s 0 9749 460 9810 1 FreeSans 1500 0 0 0 C[33]
port 54 nsew
flabel metal1 s 0 9607 460 9668 1 FreeSans 1500 0 0 0 C[34]
port 55 nsew
flabel metal1 s 0 9465 460 9526 1 FreeSans 1500 0 0 0 C[35]
port 56 nsew
flabel metal1 s 0 9323 460 9384 1 FreeSans 1500 0 0 0 C[36]
port 57 nsew
flabel metal1 s 0 9181 460 9242 1 FreeSans 1500 0 0 0 C[37]
port 58 nsew
flabel metal1 s 0 9039 460 9100 1 FreeSans 1500 0 0 0 C[38]
port 59 nsew
flabel metal1 s 0 8897 460 8958 1 FreeSans 1500 0 0 0 C[39]
port 60 nsew
flabel metal1 s 0 8755 460 8816 1 FreeSans 1500 0 0 0 C[40]
port 61 nsew
flabel metal1 s 0 8613 460 8674 1 FreeSans 1500 0 0 0 C[41]
port 62 nsew
flabel metal1 s 0 8471 460 8532 1 FreeSans 1500 0 0 0 C[42]
port 63 nsew
flabel metal1 s 0 8329 460 8390 1 FreeSans 1500 0 0 0 C[43]
port 64 nsew
flabel metal1 s 0 8187 460 8248 1 FreeSans 1500 0 0 0 C[44]
port 65 nsew
flabel metal1 s 0 8045 460 8106 1 FreeSans 1500 0 0 0 C[45]
port 66 nsew
flabel metal1 s 0 7903 460 7964 1 FreeSans 1500 0 0 0 C[46]
port 67 nsew
flabel metal1 s 0 7761 460 7822 1 FreeSans 1500 0 0 0 C[47]
port 68 nsew
flabel metal2 s 60708 19017 60752 19992 1 FreeSans 2000 0 0 0 C[0]
port 69 nsew
flabel metal2 s 58820 19017 58864 19992 1 FreeSans 2000 0 0 0 C[1]
port 70 nsew
flabel metal2 s 56932 19017 56976 19992 1 FreeSans 2000 0 0 0 C[2]
port 71 nsew
flabel metal2 s 55044 19017 55088 19992 1 FreeSans 2000 0 0 0 C[3]
port 72 nsew
flabel metal2 s 53156 19017 53200 19992 1 FreeSans 2000 0 0 0 C[4]
port 73 nsew
flabel metal2 s 51268 19017 51312 19992 1 FreeSans 2000 0 0 0 C[5]
port 74 nsew
flabel metal2 s 47492 19017 47536 19992 1 FreeSans 2000 0 0 0 C[7]
port 75 nsew
flabel metal2 s 45604 19017 45648 19992 1 FreeSans 2000 0 0 0 C[8]
port 76 nsew
flabel metal2 s 43716 19017 43760 19992 1 FreeSans 2000 0 0 0 C[9]
port 77 nsew
flabel metal2 s 41828 19017 41872 19992 1 FreeSans 2000 0 0 0 C[10]
port 78 nsew
flabel metal2 s 39940 19017 39984 19992 1 FreeSans 2000 0 0 0 C[11]
port 79 nsew
flabel metal2 s 38052 19017 38096 19992 1 FreeSans 2000 0 0 0 C[12]
port 80 nsew
flabel metal2 s 36164 19017 36208 19992 1 FreeSans 2000 0 0 0 C[13]
port 81 nsew
flabel metal2 s 34276 19017 34320 19992 1 FreeSans 2000 0 0 0 C[14]
port 82 nsew
flabel metal2 s 32388 19017 32432 19992 1 FreeSans 2000 0 0 0 C[15]
port 83 nsew
flabel metal2 s 30500 19017 30544 19992 1 FreeSans 2000 0 0 0 C[16]
port 84 nsew
flabel metal2 s 28612 19017 28656 19992 1 FreeSans 2000 0 0 0 C[17]
port 85 nsew
flabel metal2 s 26724 19017 26768 19992 1 FreeSans 2000 0 0 0 C[18]
port 86 nsew
flabel metal2 s 24836 19017 24880 19992 1 FreeSans 2000 0 0 0 C[19]
port 87 nsew
flabel metal2 s 22948 19017 22992 19992 1 FreeSans 2000 0 0 0 C[20]
port 88 nsew
flabel metal2 s 21060 19017 21104 19992 1 FreeSans 2000 0 0 0 C[21]
port 89 nsew
flabel metal2 s 19172 19017 19216 19992 1 FreeSans 2000 0 0 0 C[22]
port 90 nsew
flabel metal2 s 17284 19017 17328 19992 1 FreeSans 2000 0 0 0 C[23]
port 91 nsew
flabel metal2 s 15396 19017 15440 19992 1 FreeSans 2000 0 0 0 C[24]
port 92 nsew
flabel metal2 s 13508 19017 13552 19992 1 FreeSans 2000 0 0 0 C[25]
port 93 nsew
flabel metal2 s 11620 19017 11664 19992 1 FreeSans 2000 0 0 0 C[26]
port 94 nsew
flabel metal2 s 9732 19017 9776 19992 1 FreeSans 2000 0 0 0 C[27]
port 95 nsew
flabel metal2 s 7844 19017 7888 19992 1 FreeSans 2000 0 0 0 C[28]
port 96 nsew
flabel metal2 s 5956 19017 6000 19992 1 FreeSans 2000 0 0 0 C[29]
port 97 nsew
flabel metal2 s 4068 19017 4112 19992 1 FreeSans 2000 0 0 0 C[30]
port 98 nsew
flabel metal2 s 49380 19017 49424 20151 1 FreeSans 1000 0 0 0 C[6]
port 99 nsew
flabel metal2 s 2180 19017 2224 20184 1 FreeSans 2000 0 0 0 C[31]
port 100 nsew
flabel metal2 s 2409 0 2465 930 1 FreeSans 2000 0 0 0 C[95]
port 101 nsew
flabel metal2 s 4297 0 4353 930 1 FreeSans 2000 0 0 0 C[94]
port 102 nsew
flabel metal2 s 6185 0 6241 930 1 FreeSans 2000 0 0 0 C[93]
port 103 nsew
flabel metal2 s 8073 0 8129 930 1 FreeSans 2000 0 0 0 C[92]
port 104 nsew
flabel metal2 s 9961 0 10017 930 1 FreeSans 2000 0 0 0 C[91]
port 105 nsew
flabel metal2 s 11849 0 11905 930 1 FreeSans 2000 0 0 0 C[90]
port 106 nsew
flabel metal2 s 13737 0 13793 930 1 FreeSans 2000 0 0 0 C[89]
port 107 nsew
flabel metal2 s 15625 0 15681 930 1 FreeSans 2000 0 0 0 C[88]
port 108 nsew
flabel metal2 s 17513 0 17569 930 1 FreeSans 2000 0 0 0 C[87]
port 109 nsew
flabel metal2 s 19401 0 19457 930 1 FreeSans 2000 0 0 0 C[86]
port 110 nsew
flabel metal2 s 21289 0 21345 930 1 FreeSans 2000 0 0 0 C[85]
port 111 nsew
flabel metal2 s 23177 0 23233 930 1 FreeSans 2000 0 0 0 C[84]
port 112 nsew
flabel metal2 s 25065 0 25121 930 1 FreeSans 2000 0 0 0 C[83]
port 113 nsew
flabel metal2 s 26953 0 27009 930 1 FreeSans 2000 0 0 0 C[82]
port 114 nsew
flabel metal2 s 28841 0 28897 930 1 FreeSans 2000 0 0 0 C[81]
port 115 nsew
flabel metal2 s 30729 0 30785 930 1 FreeSans 2000 0 0 0 C[80]
port 116 nsew
flabel metal2 s 32617 0 32673 930 1 FreeSans 2000 0 0 0 C[79]
port 117 nsew
flabel metal2 s 34505 0 34561 930 1 FreeSans 2000 0 0 0 C[78]
port 118 nsew
flabel metal2 s 36393 0 36449 930 1 FreeSans 2000 0 0 0 C[77]
port 119 nsew
flabel metal2 s 38281 0 38337 930 1 FreeSans 2000 0 0 0 C[76]
port 120 nsew
flabel metal2 s 40169 0 40225 930 1 FreeSans 2000 0 0 0 C[75]
port 121 nsew
flabel metal2 s 42057 0 42113 930 1 FreeSans 2000 0 0 0 C[74]
port 122 nsew
flabel metal2 s 43945 0 44001 930 1 FreeSans 2000 0 0 0 C[73]
port 123 nsew
flabel metal2 s 45833 0 45889 930 1 FreeSans 2000 0 0 0 C[72]
port 124 nsew
flabel metal2 s 47721 0 47777 930 1 FreeSans 2000 0 0 0 C[71]
port 125 nsew
flabel metal2 s 49609 0 49665 930 1 FreeSans 2000 0 0 0 C[70]
port 126 nsew
flabel metal2 s 51497 0 51553 930 1 FreeSans 2000 0 0 0 C[69]
port 127 nsew
flabel metal2 s 53385 0 53441 930 1 FreeSans 2000 0 0 0 C[68]
port 128 nsew
flabel metal2 s 55273 0 55329 930 1 FreeSans 2000 0 0 0 C[67]
port 129 nsew
flabel metal2 s 57161 0 57217 930 1 FreeSans 2000 0 0 0 C[66]
port 130 nsew
flabel metal2 s 59049 0 59105 930 1 FreeSans 2000 0 0 0 C[65]
port 131 nsew
flabel metal2 s 60937 0 60993 930 1 FreeSans 2000 0 0 0 C[64]
port 132 nsew
<< end >>
