magic
tech sky130A
timestamp 1656729169
<< metal3 >>
rect -90 76 90 90
rect -90 -76 -76 76
rect 76 -76 90 76
rect -90 -90 90 -76
<< via3 >>
rect -76 -76 76 76
<< metal4 >>
rect -90 76 90 90
rect -90 -76 -76 76
rect 76 -76 90 76
rect -90 -90 90 -76
<< properties >>
string GDS_END 9339418
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/merge/design_merged.gds
string GDS_START 9338262
<< end >>
