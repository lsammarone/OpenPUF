magic
tech sky130A
magscale 1 2
timestamp 1654736712
<< metal4 >>
rect -180 598 180 737
rect -180 362 -118 598
rect 118 362 180 598
rect -180 278 180 362
rect -180 42 -118 278
rect 118 42 180 278
rect -180 -42 180 42
rect -180 -278 -118 -42
rect 118 -278 180 -42
rect -180 -362 180 -278
rect -180 -598 -118 -362
rect 118 -598 180 -362
rect -180 -737 180 -598
<< via4 >>
rect -118 362 118 598
rect -118 42 118 278
rect -118 -278 118 -42
rect -118 -598 118 -362
<< metal5 >>
rect -180 598 180 737
rect -180 362 -118 598
rect 118 362 180 598
rect -180 278 180 362
rect -180 42 -118 278
rect 118 42 180 278
rect -180 -42 180 42
rect -180 -278 -118 -42
rect 118 -278 180 -42
rect -180 -362 180 -278
rect -180 -598 -118 -362
rect 118 -598 180 -362
rect -180 -737 180 -598
<< end >>
