magic
tech sky130A
magscale 1 2
timestamp 1656729169
<< nwell >>
rect 15089 3413 15613 3591
<< pwell >>
rect 9527 3441 9757 3559
rect 24565 3445 24793 3571
<< psubdiff >>
rect 9553 3517 9731 3533
rect 24591 3525 24767 3545
rect 9553 3483 9591 3517
rect 9625 3483 9659 3517
rect 9693 3483 9731 3517
rect 9553 3467 9731 3483
rect 24591 3491 24628 3525
rect 24662 3491 24696 3525
rect 24730 3491 24767 3525
rect 24591 3471 24767 3491
<< nsubdiff >>
rect 15181 3508 15389 3525
rect 15181 3474 15234 3508
rect 15268 3474 15302 3508
rect 15336 3474 15389 3508
rect 15181 3457 15389 3474
<< psubdiffcont >>
rect 9591 3483 9625 3517
rect 9659 3483 9693 3517
rect 24628 3491 24662 3525
rect 24696 3491 24730 3525
<< nsubdiffcont >>
rect 15234 3474 15268 3508
rect 15302 3474 15336 3508
<< locali >>
rect 9425 3517 9723 3533
rect 24599 3532 24759 3545
rect 24520 3525 24759 3532
rect 9425 3483 9591 3517
rect 9625 3483 9659 3517
rect 9693 3483 9723 3517
rect 9425 3467 9723 3483
rect 15189 3508 15381 3525
rect 15189 3474 15234 3508
rect 15268 3474 15302 3508
rect 15336 3474 15381 3508
rect 24520 3491 24628 3525
rect 24662 3491 24696 3525
rect 24730 3491 24759 3525
rect 24520 3488 24759 3491
rect 15189 3429 15381 3474
rect 24599 3471 24759 3488
rect 15259 3213 15297 3217
rect 15259 3179 15261 3213
rect 15295 3179 15297 3213
rect 15259 3175 15297 3179
rect 16615 3126 16661 3129
rect 16615 3092 16621 3126
rect 16655 3092 16661 3126
rect 16615 3089 16661 3092
<< viali >>
rect 15261 3179 15295 3213
rect 16621 3092 16655 3126
rect 19160 3088 19194 3122
<< metal1 >>
rect 22909 3645 22969 3677
rect 9773 3642 11032 3643
rect 9773 3597 11503 3642
rect 9396 3275 10170 3352
rect 9396 3159 9485 3275
rect 9793 3159 10170 3275
rect 9396 2898 10170 3159
rect 11443 3161 11503 3597
rect 22909 3599 24650 3645
rect 15167 3441 15411 3459
rect 15167 3389 15199 3441
rect 15251 3389 15263 3441
rect 15315 3389 15327 3441
rect 15379 3389 15411 3441
rect 15167 3371 15411 3389
rect 18933 3453 19177 3461
rect 18933 3443 19201 3453
rect 18933 3391 18965 3443
rect 19017 3391 19029 3443
rect 19081 3391 19093 3443
rect 19145 3391 19201 3443
rect 18933 3381 19201 3391
rect 18933 3373 19177 3381
rect 19213 3367 19413 3463
rect 15253 3213 15309 3229
rect 15253 3179 15261 3213
rect 15295 3179 15309 3213
rect 15253 3161 15309 3179
rect 11443 3101 15309 3161
rect 16599 3135 16673 3145
rect 11443 2660 11503 3101
rect 16599 3083 16611 3135
rect 16663 3083 16673 3135
rect 16599 3077 16673 3083
rect 19148 3135 19230 3146
rect 22909 3135 22969 3599
rect 19148 3122 22969 3135
rect 19148 3088 19160 3122
rect 19194 3088 22969 3122
rect 19148 3075 22969 3088
rect 19148 3064 19230 3075
rect 17031 2899 17315 2917
rect 17031 2847 17051 2899
rect 17103 2847 17115 2899
rect 17167 2847 17179 2899
rect 17231 2847 17243 2899
rect 17295 2847 17315 2899
rect 17031 2829 17315 2847
rect 19219 2823 19419 2919
rect 10764 2604 11503 2660
rect 22909 2661 22969 3075
rect 24450 3317 25206 3374
rect 24450 3201 24573 3317
rect 24881 3201 25206 3317
rect 24450 2880 25206 3201
rect 22909 2615 24760 2661
rect 22909 2583 22969 2615
rect 32393 782 32622 859
<< via1 >>
rect 9485 3159 9793 3275
rect 15199 3389 15251 3441
rect 15263 3389 15315 3441
rect 15327 3389 15379 3441
rect 18965 3391 19017 3443
rect 19029 3391 19081 3443
rect 19093 3391 19145 3443
rect 16611 3126 16663 3135
rect 16611 3092 16621 3126
rect 16621 3092 16655 3126
rect 16655 3092 16663 3126
rect 16611 3083 16663 3092
rect 17051 2847 17103 2899
rect 17115 2847 17167 2899
rect 17179 2847 17231 2899
rect 17243 2847 17295 2899
rect 24573 3201 24881 3317
<< metal2 >>
rect 3730 5465 3774 6257
rect 5618 5465 5662 6257
rect 7506 5465 7550 6257
rect 9394 5465 9438 6257
rect 11282 5465 11326 6257
rect 13170 5465 13214 6257
rect 15058 5465 15102 6257
rect 16946 5465 16990 6257
rect 18834 5465 18878 6257
rect 20722 5465 20766 6257
rect 22610 5465 22654 6257
rect 24498 5465 24542 6257
rect 26386 5465 26430 6257
rect 28274 5465 28318 6257
rect 30162 5465 30206 6257
rect 0 5226 1947 5262
rect 0 1036 36 5226
rect 30088 5224 32830 5260
rect 169 4747 1959 4783
rect 30177 4747 32667 4783
rect 169 1511 205 4747
rect 15177 3443 15401 3469
rect 15177 3387 15181 3443
rect 15237 3441 15261 3443
rect 15317 3441 15341 3443
rect 15251 3389 15261 3441
rect 15317 3389 15327 3441
rect 15237 3387 15261 3389
rect 15317 3387 15341 3389
rect 15397 3387 15401 3443
rect 15177 3361 15401 3387
rect 18943 3445 19167 3471
rect 18943 3389 18947 3445
rect 19003 3443 19027 3445
rect 19083 3443 19107 3445
rect 19017 3391 19027 3443
rect 19083 3391 19093 3443
rect 19003 3389 19027 3391
rect 19083 3389 19107 3391
rect 19163 3389 19167 3445
rect 18943 3363 19167 3389
rect 24573 3317 24881 3327
rect 9485 3275 9793 3285
rect 24573 3191 24881 3201
rect 9485 3149 9793 3159
rect 16605 3135 16669 3145
rect 429 3111 569 3131
rect 429 3055 463 3111
rect 519 3103 569 3111
rect 16605 3103 16611 3135
rect 519 3083 16611 3103
rect 16663 3083 16669 3135
rect 519 3071 16669 3083
rect 519 3055 569 3071
rect 429 3035 569 3055
rect 17041 2901 17305 2927
rect 17041 2899 17065 2901
rect 17121 2899 17145 2901
rect 17201 2899 17225 2901
rect 17281 2899 17305 2901
rect 17041 2847 17051 2899
rect 17295 2847 17305 2899
rect 17041 2845 17065 2847
rect 17121 2845 17145 2847
rect 17201 2845 17225 2847
rect 17281 2845 17305 2847
rect 17041 2819 17305 2845
rect 613 2555 1639 2556
rect 2503 2555 3529 2556
rect 393 2367 4355 2555
rect 613 2110 1639 2367
rect 2503 2110 3529 2367
rect 393 2001 4276 2110
rect 32631 1511 32667 4747
rect 169 1475 437 1511
rect 32417 1475 32669 1511
rect 0 1000 514 1036
rect 32794 1020 32830 5224
rect 32446 984 32830 1020
rect 413 1 457 793
rect 2301 1 2345 793
rect 4189 1 4233 793
rect 6077 1 6121 793
rect 7965 1 8009 793
rect 9853 1 9897 793
rect 11741 1 11785 793
rect 13629 1 13673 793
rect 15517 1 15561 793
rect 17405 1 17449 793
rect 19293 1 19337 793
rect 21181 1 21225 793
rect 23069 1 23113 793
rect 24957 1 25001 793
rect 26845 1 26889 793
rect 28733 1 28777 793
rect 30621 1 30665 793
<< via2 >>
rect 15181 3441 15237 3443
rect 15261 3441 15317 3443
rect 15341 3441 15397 3443
rect 15181 3389 15199 3441
rect 15199 3389 15237 3441
rect 15261 3389 15263 3441
rect 15263 3389 15315 3441
rect 15315 3389 15317 3441
rect 15341 3389 15379 3441
rect 15379 3389 15397 3441
rect 15181 3387 15237 3389
rect 15261 3387 15317 3389
rect 15341 3387 15397 3389
rect 18947 3443 19003 3445
rect 19027 3443 19083 3445
rect 19107 3443 19163 3445
rect 18947 3391 18965 3443
rect 18965 3391 19003 3443
rect 19027 3391 19029 3443
rect 19029 3391 19081 3443
rect 19081 3391 19083 3443
rect 19107 3391 19145 3443
rect 19145 3391 19163 3443
rect 18947 3389 19003 3391
rect 19027 3389 19083 3391
rect 19107 3389 19163 3391
rect 9491 3189 9547 3245
rect 9571 3189 9627 3245
rect 9651 3189 9707 3245
rect 9731 3189 9787 3245
rect 24579 3231 24635 3287
rect 24659 3231 24715 3287
rect 24739 3231 24795 3287
rect 24819 3231 24875 3287
rect 463 3055 519 3111
rect 17065 2899 17121 2901
rect 17145 2899 17201 2901
rect 17225 2899 17281 2901
rect 17065 2847 17103 2899
rect 17103 2847 17115 2899
rect 17115 2847 17121 2899
rect 17145 2847 17167 2899
rect 17167 2847 17179 2899
rect 17179 2847 17201 2899
rect 17225 2847 17231 2899
rect 17231 2847 17243 2899
rect 17243 2847 17281 2899
rect 17065 2845 17121 2847
rect 17145 2845 17201 2847
rect 17225 2845 17281 2847
<< metal3 >>
rect 1948 6167 2276 6193
rect 1948 6103 1960 6167
rect 2024 6103 2040 6167
rect 2104 6103 2120 6167
rect 2184 6103 2200 6167
rect 2264 6103 2276 6167
rect 1948 6077 2276 6103
rect 5724 6167 6052 6193
rect 5724 6103 5736 6167
rect 5800 6103 5816 6167
rect 5880 6103 5896 6167
rect 5960 6103 5976 6167
rect 6040 6103 6052 6167
rect 5724 6077 6052 6103
rect 9500 6167 9828 6193
rect 9500 6103 9512 6167
rect 9576 6103 9592 6167
rect 9656 6103 9672 6167
rect 9736 6103 9752 6167
rect 9816 6103 9828 6167
rect 9500 6077 9828 6103
rect 13276 6167 13604 6193
rect 13276 6103 13288 6167
rect 13352 6103 13368 6167
rect 13432 6103 13448 6167
rect 13512 6103 13528 6167
rect 13592 6103 13604 6167
rect 13276 6077 13604 6103
rect 17046 6167 17374 6193
rect 17046 6103 17058 6167
rect 17122 6103 17138 6167
rect 17202 6103 17218 6167
rect 17282 6103 17298 6167
rect 17362 6103 17374 6167
rect 17046 6077 17374 6103
rect 20822 6167 21150 6193
rect 20822 6103 20834 6167
rect 20898 6103 20914 6167
rect 20978 6103 20994 6167
rect 21058 6103 21074 6167
rect 21138 6103 21150 6167
rect 20822 6077 21150 6103
rect 24598 6167 24926 6193
rect 24598 6103 24610 6167
rect 24674 6103 24690 6167
rect 24754 6103 24770 6167
rect 24834 6103 24850 6167
rect 24914 6103 24926 6167
rect 24598 6077 24926 6103
rect 28374 6167 28702 6193
rect 28374 6103 28386 6167
rect 28450 6103 28466 6167
rect 28530 6103 28546 6167
rect 28610 6103 28626 6167
rect 28690 6103 28702 6167
rect 28374 6077 28702 6103
rect 3836 4043 4164 4069
rect 3836 3979 3848 4043
rect 3912 3979 3928 4043
rect 3992 3979 4008 4043
rect 4072 3979 4088 4043
rect 4152 3979 4164 4043
rect 3836 3953 4164 3979
rect 7612 4043 7940 4069
rect 7612 3979 7624 4043
rect 7688 3979 7704 4043
rect 7768 3979 7784 4043
rect 7848 3979 7864 4043
rect 7928 3979 7940 4043
rect 7612 3953 7940 3979
rect 11388 4043 11716 4069
rect 11388 3979 11400 4043
rect 11464 3979 11480 4043
rect 11544 3979 11560 4043
rect 11624 3979 11640 4043
rect 11704 3979 11716 4043
rect 11388 3953 11716 3979
rect 15164 4043 15492 4069
rect 15164 3979 15176 4043
rect 15240 3979 15256 4043
rect 15320 3979 15336 4043
rect 15400 3979 15416 4043
rect 15480 3979 15492 4043
rect 15164 3953 15492 3979
rect 18934 4043 19262 4069
rect 18934 3979 18946 4043
rect 19010 3979 19026 4043
rect 19090 3979 19106 4043
rect 19170 3979 19186 4043
rect 19250 3979 19262 4043
rect 18934 3953 19262 3979
rect 22710 4043 23038 4069
rect 22710 3979 22722 4043
rect 22786 3979 22802 4043
rect 22866 3979 22882 4043
rect 22946 3979 22962 4043
rect 23026 3979 23038 4043
rect 22710 3953 23038 3979
rect 26486 4043 26814 4069
rect 26486 3979 26498 4043
rect 26562 3979 26578 4043
rect 26642 3979 26658 4043
rect 26722 3979 26738 4043
rect 26802 3979 26814 4043
rect 26486 3953 26814 3979
rect 15167 3447 15411 3464
rect 15167 3383 15177 3447
rect 15241 3383 15257 3447
rect 15321 3383 15337 3447
rect 15401 3383 15411 3447
rect 15167 3366 15411 3383
rect 18933 3449 19177 3466
rect 18933 3385 18943 3449
rect 19007 3385 19023 3449
rect 19087 3385 19103 3449
rect 19167 3385 19177 3449
rect 18933 3368 19177 3385
rect 24563 3291 24891 3322
rect 9475 3249 9803 3280
rect 9475 3185 9487 3249
rect 9551 3185 9567 3249
rect 9631 3185 9647 3249
rect 9711 3185 9727 3249
rect 9791 3185 9803 3249
rect 24563 3227 24575 3291
rect 24639 3227 24655 3291
rect 24719 3227 24735 3291
rect 24799 3227 24815 3291
rect 24879 3227 24891 3291
rect 24563 3196 24891 3227
rect 9475 3154 9803 3185
rect 18 3111 554 3129
rect 18 3055 463 3111
rect 519 3055 554 3111
rect 18 3036 554 3055
rect 17031 2905 17315 2922
rect 17031 2841 17061 2905
rect 17125 2841 17141 2905
rect 17205 2841 17221 2905
rect 17285 2841 17315 2905
rect 17031 2824 17315 2841
rect 3806 2279 4134 2305
rect 3806 2215 3818 2279
rect 3882 2215 3898 2279
rect 3962 2215 3978 2279
rect 4042 2215 4058 2279
rect 4122 2215 4134 2279
rect 3806 2189 4134 2215
rect 7582 2279 7910 2305
rect 7582 2215 7594 2279
rect 7658 2215 7674 2279
rect 7738 2215 7754 2279
rect 7818 2215 7834 2279
rect 7898 2215 7910 2279
rect 7582 2189 7910 2215
rect 11358 2279 11686 2305
rect 11358 2215 11370 2279
rect 11434 2215 11450 2279
rect 11514 2215 11530 2279
rect 11594 2215 11610 2279
rect 11674 2215 11686 2279
rect 11358 2189 11686 2215
rect 15134 2279 15462 2305
rect 15134 2215 15146 2279
rect 15210 2215 15226 2279
rect 15290 2215 15306 2279
rect 15370 2215 15386 2279
rect 15450 2215 15462 2279
rect 15134 2189 15462 2215
rect 18904 2279 19232 2305
rect 18904 2215 18916 2279
rect 18980 2215 18996 2279
rect 19060 2215 19076 2279
rect 19140 2215 19156 2279
rect 19220 2215 19232 2279
rect 18904 2189 19232 2215
rect 22680 2279 23008 2305
rect 22680 2215 22692 2279
rect 22756 2215 22772 2279
rect 22836 2215 22852 2279
rect 22916 2215 22932 2279
rect 22996 2215 23008 2279
rect 22680 2189 23008 2215
rect 26456 2279 26784 2305
rect 26456 2215 26468 2279
rect 26532 2215 26548 2279
rect 26612 2215 26628 2279
rect 26692 2215 26708 2279
rect 26772 2215 26784 2279
rect 26456 2189 26784 2215
rect 1918 155 2246 181
rect 1918 91 1930 155
rect 1994 91 2010 155
rect 2074 91 2090 155
rect 2154 91 2170 155
rect 2234 91 2246 155
rect 1918 65 2246 91
rect 5694 155 6022 181
rect 5694 91 5706 155
rect 5770 91 5786 155
rect 5850 91 5866 155
rect 5930 91 5946 155
rect 6010 91 6022 155
rect 5694 65 6022 91
rect 9470 155 9798 181
rect 9470 91 9482 155
rect 9546 91 9562 155
rect 9626 91 9642 155
rect 9706 91 9722 155
rect 9786 91 9798 155
rect 9470 65 9798 91
rect 13246 155 13574 181
rect 13246 91 13258 155
rect 13322 91 13338 155
rect 13402 91 13418 155
rect 13482 91 13498 155
rect 13562 91 13574 155
rect 13246 65 13574 91
rect 17022 155 17350 181
rect 17022 91 17034 155
rect 17098 91 17114 155
rect 17178 91 17194 155
rect 17258 91 17274 155
rect 17338 91 17350 155
rect 17022 65 17350 91
rect 20792 155 21120 181
rect 20792 91 20804 155
rect 20868 91 20884 155
rect 20948 91 20964 155
rect 21028 91 21044 155
rect 21108 91 21120 155
rect 20792 65 21120 91
rect 24568 155 24896 181
rect 24568 91 24580 155
rect 24644 91 24660 155
rect 24724 91 24740 155
rect 24804 91 24820 155
rect 24884 91 24896 155
rect 24568 65 24896 91
rect 28344 155 28672 181
rect 28344 91 28356 155
rect 28420 91 28436 155
rect 28500 91 28516 155
rect 28580 91 28596 155
rect 28660 91 28672 155
rect 28344 65 28672 91
<< via3 >>
rect 1960 6103 2024 6167
rect 2040 6103 2104 6167
rect 2120 6103 2184 6167
rect 2200 6103 2264 6167
rect 5736 6103 5800 6167
rect 5816 6103 5880 6167
rect 5896 6103 5960 6167
rect 5976 6103 6040 6167
rect 9512 6103 9576 6167
rect 9592 6103 9656 6167
rect 9672 6103 9736 6167
rect 9752 6103 9816 6167
rect 13288 6103 13352 6167
rect 13368 6103 13432 6167
rect 13448 6103 13512 6167
rect 13528 6103 13592 6167
rect 17058 6103 17122 6167
rect 17138 6103 17202 6167
rect 17218 6103 17282 6167
rect 17298 6103 17362 6167
rect 20834 6103 20898 6167
rect 20914 6103 20978 6167
rect 20994 6103 21058 6167
rect 21074 6103 21138 6167
rect 24610 6103 24674 6167
rect 24690 6103 24754 6167
rect 24770 6103 24834 6167
rect 24850 6103 24914 6167
rect 28386 6103 28450 6167
rect 28466 6103 28530 6167
rect 28546 6103 28610 6167
rect 28626 6103 28690 6167
rect 3848 3979 3912 4043
rect 3928 3979 3992 4043
rect 4008 3979 4072 4043
rect 4088 3979 4152 4043
rect 7624 3979 7688 4043
rect 7704 3979 7768 4043
rect 7784 3979 7848 4043
rect 7864 3979 7928 4043
rect 11400 3979 11464 4043
rect 11480 3979 11544 4043
rect 11560 3979 11624 4043
rect 11640 3979 11704 4043
rect 15176 3979 15240 4043
rect 15256 3979 15320 4043
rect 15336 3979 15400 4043
rect 15416 3979 15480 4043
rect 18946 3979 19010 4043
rect 19026 3979 19090 4043
rect 19106 3979 19170 4043
rect 19186 3979 19250 4043
rect 22722 3979 22786 4043
rect 22802 3979 22866 4043
rect 22882 3979 22946 4043
rect 22962 3979 23026 4043
rect 26498 3979 26562 4043
rect 26578 3979 26642 4043
rect 26658 3979 26722 4043
rect 26738 3979 26802 4043
rect 15177 3443 15241 3447
rect 15177 3387 15181 3443
rect 15181 3387 15237 3443
rect 15237 3387 15241 3443
rect 15177 3383 15241 3387
rect 15257 3443 15321 3447
rect 15257 3387 15261 3443
rect 15261 3387 15317 3443
rect 15317 3387 15321 3443
rect 15257 3383 15321 3387
rect 15337 3443 15401 3447
rect 15337 3387 15341 3443
rect 15341 3387 15397 3443
rect 15397 3387 15401 3443
rect 15337 3383 15401 3387
rect 18943 3445 19007 3449
rect 18943 3389 18947 3445
rect 18947 3389 19003 3445
rect 19003 3389 19007 3445
rect 18943 3385 19007 3389
rect 19023 3445 19087 3449
rect 19023 3389 19027 3445
rect 19027 3389 19083 3445
rect 19083 3389 19087 3445
rect 19023 3385 19087 3389
rect 19103 3445 19167 3449
rect 19103 3389 19107 3445
rect 19107 3389 19163 3445
rect 19163 3389 19167 3445
rect 19103 3385 19167 3389
rect 9487 3245 9551 3249
rect 9487 3189 9491 3245
rect 9491 3189 9547 3245
rect 9547 3189 9551 3245
rect 9487 3185 9551 3189
rect 9567 3245 9631 3249
rect 9567 3189 9571 3245
rect 9571 3189 9627 3245
rect 9627 3189 9631 3245
rect 9567 3185 9631 3189
rect 9647 3245 9711 3249
rect 9647 3189 9651 3245
rect 9651 3189 9707 3245
rect 9707 3189 9711 3245
rect 9647 3185 9711 3189
rect 9727 3245 9791 3249
rect 9727 3189 9731 3245
rect 9731 3189 9787 3245
rect 9787 3189 9791 3245
rect 9727 3185 9791 3189
rect 24575 3287 24639 3291
rect 24575 3231 24579 3287
rect 24579 3231 24635 3287
rect 24635 3231 24639 3287
rect 24575 3227 24639 3231
rect 24655 3287 24719 3291
rect 24655 3231 24659 3287
rect 24659 3231 24715 3287
rect 24715 3231 24719 3287
rect 24655 3227 24719 3231
rect 24735 3287 24799 3291
rect 24735 3231 24739 3287
rect 24739 3231 24795 3287
rect 24795 3231 24799 3287
rect 24735 3227 24799 3231
rect 24815 3287 24879 3291
rect 24815 3231 24819 3287
rect 24819 3231 24875 3287
rect 24875 3231 24879 3287
rect 24815 3227 24879 3231
rect 17061 2901 17125 2905
rect 17061 2845 17065 2901
rect 17065 2845 17121 2901
rect 17121 2845 17125 2901
rect 17061 2841 17125 2845
rect 17141 2901 17205 2905
rect 17141 2845 17145 2901
rect 17145 2845 17201 2901
rect 17201 2845 17205 2901
rect 17141 2841 17205 2845
rect 17221 2901 17285 2905
rect 17221 2845 17225 2901
rect 17225 2845 17281 2901
rect 17281 2845 17285 2901
rect 17221 2841 17285 2845
rect 3818 2215 3882 2279
rect 3898 2215 3962 2279
rect 3978 2215 4042 2279
rect 4058 2215 4122 2279
rect 7594 2215 7658 2279
rect 7674 2215 7738 2279
rect 7754 2215 7818 2279
rect 7834 2215 7898 2279
rect 11370 2215 11434 2279
rect 11450 2215 11514 2279
rect 11530 2215 11594 2279
rect 11610 2215 11674 2279
rect 15146 2215 15210 2279
rect 15226 2215 15290 2279
rect 15306 2215 15370 2279
rect 15386 2215 15450 2279
rect 18916 2215 18980 2279
rect 18996 2215 19060 2279
rect 19076 2215 19140 2279
rect 19156 2215 19220 2279
rect 22692 2215 22756 2279
rect 22772 2215 22836 2279
rect 22852 2215 22916 2279
rect 22932 2215 22996 2279
rect 26468 2215 26532 2279
rect 26548 2215 26612 2279
rect 26628 2215 26692 2279
rect 26708 2215 26772 2279
rect 1930 91 1994 155
rect 2010 91 2074 155
rect 2090 91 2154 155
rect 2170 91 2234 155
rect 5706 91 5770 155
rect 5786 91 5850 155
rect 5866 91 5930 155
rect 5946 91 6010 155
rect 9482 91 9546 155
rect 9562 91 9626 155
rect 9642 91 9706 155
rect 9722 91 9786 155
rect 13258 91 13322 155
rect 13338 91 13402 155
rect 13418 91 13482 155
rect 13498 91 13562 155
rect 17034 91 17098 155
rect 17114 91 17178 155
rect 17194 91 17258 155
rect 17274 91 17338 155
rect 20804 91 20868 155
rect 20884 91 20948 155
rect 20964 91 21028 155
rect 21044 91 21108 155
rect 24580 91 24644 155
rect 24660 91 24724 155
rect 24740 91 24804 155
rect 24820 91 24884 155
rect 28356 91 28420 155
rect 28436 91 28500 155
rect 28516 91 28580 155
rect 28596 91 28660 155
<< metal4 >>
rect 1915 6194 2253 6259
rect 1915 6167 2267 6194
rect 1915 6103 1960 6167
rect 2024 6103 2040 6167
rect 2104 6103 2120 6167
rect 2184 6103 2200 6167
rect 2264 6103 2267 6167
rect 1915 6076 2267 6103
rect 1915 155 2253 6076
rect 1915 91 1930 155
rect 1994 91 2010 155
rect 2074 91 2090 155
rect 2154 91 2170 155
rect 2234 91 2253 155
rect 1915 1 2253 91
rect 3813 4070 4151 6257
rect 5699 6194 6037 6258
rect 5699 6167 6043 6194
rect 5699 6103 5736 6167
rect 5800 6103 5816 6167
rect 5880 6103 5896 6167
rect 5960 6103 5976 6167
rect 6040 6103 6043 6167
rect 5699 6076 6043 6103
rect 3813 4043 4155 4070
rect 3813 3979 3848 4043
rect 3912 3979 3928 4043
rect 3992 3979 4008 4043
rect 4072 3979 4088 4043
rect 4152 3979 4155 4043
rect 3813 3952 4155 3979
rect 3813 2279 4151 3952
rect 3813 2215 3818 2279
rect 3882 2215 3898 2279
rect 3962 2215 3978 2279
rect 4042 2215 4058 2279
rect 4122 2215 4151 2279
rect 3813 1 4151 2215
rect 5699 155 6037 6076
rect 5699 91 5706 155
rect 5770 91 5786 155
rect 5850 91 5866 155
rect 5930 91 5946 155
rect 6010 91 6037 155
rect 5699 0 6037 91
rect 7589 4070 7927 6257
rect 9473 6194 9811 6259
rect 9473 6167 9819 6194
rect 9473 6103 9512 6167
rect 9576 6103 9592 6167
rect 9656 6103 9672 6167
rect 9736 6103 9752 6167
rect 9816 6103 9819 6167
rect 9473 6076 9819 6103
rect 7589 4043 7931 4070
rect 7589 3979 7624 4043
rect 7688 3979 7704 4043
rect 7768 3979 7784 4043
rect 7848 3979 7864 4043
rect 7928 3979 7931 4043
rect 7589 3952 7931 3979
rect 7589 2279 7927 3952
rect 7589 2215 7594 2279
rect 7658 2215 7674 2279
rect 7738 2215 7754 2279
rect 7818 2215 7834 2279
rect 7898 2215 7927 2279
rect 7589 1 7927 2215
rect 9473 3249 9811 6076
rect 9473 3185 9487 3249
rect 9551 3185 9567 3249
rect 9631 3185 9647 3249
rect 9711 3185 9727 3249
rect 9791 3185 9811 3249
rect 9473 155 9811 3185
rect 9473 91 9482 155
rect 9546 91 9562 155
rect 9626 91 9642 155
rect 9706 91 9722 155
rect 9786 91 9811 155
rect 9473 1 9811 91
rect 11359 4070 11697 6257
rect 13251 6194 13589 6259
rect 13251 6167 13595 6194
rect 13251 6103 13288 6167
rect 13352 6103 13368 6167
rect 13432 6103 13448 6167
rect 13512 6103 13528 6167
rect 13592 6103 13595 6167
rect 13251 6076 13595 6103
rect 11359 4043 11707 4070
rect 11359 3979 11400 4043
rect 11464 3979 11480 4043
rect 11544 3979 11560 4043
rect 11624 3979 11640 4043
rect 11704 3979 11707 4043
rect 11359 3952 11707 3979
rect 11359 2279 11697 3952
rect 11359 2215 11370 2279
rect 11434 2215 11450 2279
rect 11514 2215 11530 2279
rect 11594 2215 11610 2279
rect 11674 2215 11697 2279
rect 11359 1 11697 2215
rect 13251 155 13589 6076
rect 13251 91 13258 155
rect 13322 91 13338 155
rect 13402 91 13418 155
rect 13482 91 13498 155
rect 13562 91 13589 155
rect 13251 1 13589 91
rect 15127 4070 15465 6257
rect 17019 6194 17357 6259
rect 17019 6167 17365 6194
rect 17019 6103 17058 6167
rect 17122 6103 17138 6167
rect 17202 6103 17218 6167
rect 17282 6103 17298 6167
rect 17362 6103 17365 6167
rect 17019 6076 17365 6103
rect 15127 4043 15483 4070
rect 15127 3979 15176 4043
rect 15240 3979 15256 4043
rect 15320 3979 15336 4043
rect 15400 3979 15416 4043
rect 15480 3979 15483 4043
rect 15127 3952 15483 3979
rect 15127 3447 15465 3952
rect 15127 3383 15177 3447
rect 15241 3383 15257 3447
rect 15321 3383 15337 3447
rect 15401 3383 15465 3447
rect 15127 2279 15465 3383
rect 15127 2215 15146 2279
rect 15210 2215 15226 2279
rect 15290 2215 15306 2279
rect 15370 2215 15386 2279
rect 15450 2215 15465 2279
rect 15127 1 15465 2215
rect 17019 2905 17357 6076
rect 17019 2841 17061 2905
rect 17125 2841 17141 2905
rect 17205 2841 17221 2905
rect 17285 2841 17357 2905
rect 17019 155 17357 2841
rect 17019 91 17034 155
rect 17098 91 17114 155
rect 17178 91 17194 155
rect 17258 91 17274 155
rect 17338 91 17357 155
rect 17019 1 17357 91
rect 18899 4070 19237 6257
rect 20791 6194 21129 6259
rect 20791 6167 21141 6194
rect 20791 6103 20834 6167
rect 20898 6103 20914 6167
rect 20978 6103 20994 6167
rect 21058 6103 21074 6167
rect 21138 6103 21141 6167
rect 20791 6076 21141 6103
rect 18899 4043 19253 4070
rect 18899 3979 18946 4043
rect 19010 3979 19026 4043
rect 19090 3979 19106 4043
rect 19170 3979 19186 4043
rect 19250 3979 19253 4043
rect 18899 3952 19253 3979
rect 18899 3449 19237 3952
rect 18899 3385 18943 3449
rect 19007 3385 19023 3449
rect 19087 3385 19103 3449
rect 19167 3385 19237 3449
rect 18899 2279 19237 3385
rect 18899 2215 18916 2279
rect 18980 2215 18996 2279
rect 19060 2215 19076 2279
rect 19140 2215 19156 2279
rect 19220 2215 19237 2279
rect 18899 1 19237 2215
rect 20791 155 21129 6076
rect 20791 91 20804 155
rect 20868 91 20884 155
rect 20948 91 20964 155
rect 21028 91 21044 155
rect 21108 91 21129 155
rect 20791 1 21129 91
rect 22667 4070 23005 6257
rect 24561 6194 24899 6259
rect 24561 6167 24917 6194
rect 24561 6103 24610 6167
rect 24674 6103 24690 6167
rect 24754 6103 24770 6167
rect 24834 6103 24850 6167
rect 24914 6103 24917 6167
rect 24561 6076 24917 6103
rect 22667 4043 23029 4070
rect 22667 3979 22722 4043
rect 22786 3979 22802 4043
rect 22866 3979 22882 4043
rect 22946 3979 22962 4043
rect 23026 3979 23029 4043
rect 22667 3952 23029 3979
rect 22667 2279 23005 3952
rect 22667 2215 22692 2279
rect 22756 2215 22772 2279
rect 22836 2215 22852 2279
rect 22916 2215 22932 2279
rect 22996 2215 23005 2279
rect 22667 1 23005 2215
rect 24561 3291 24899 6076
rect 24561 3227 24575 3291
rect 24639 3227 24655 3291
rect 24719 3227 24735 3291
rect 24799 3227 24815 3291
rect 24879 3227 24899 3291
rect 24561 155 24899 3227
rect 24561 91 24580 155
rect 24644 91 24660 155
rect 24724 91 24740 155
rect 24804 91 24820 155
rect 24884 91 24899 155
rect 24561 1 24899 91
rect 26463 4070 26801 6257
rect 28349 6194 28687 6258
rect 28349 6167 28693 6194
rect 28349 6103 28386 6167
rect 28450 6103 28466 6167
rect 28530 6103 28546 6167
rect 28610 6103 28626 6167
rect 28690 6103 28693 6167
rect 28349 6076 28693 6103
rect 26463 4043 26805 4070
rect 26463 3979 26498 4043
rect 26562 3979 26578 4043
rect 26642 3979 26658 4043
rect 26722 3979 26738 4043
rect 26802 3979 26805 4043
rect 26463 3952 26805 3979
rect 26463 2279 26801 3952
rect 26463 2215 26468 2279
rect 26532 2215 26548 2279
rect 26612 2215 26628 2279
rect 26692 2215 26708 2279
rect 26772 2215 26801 2279
rect 26463 1 26801 2215
rect 28349 155 28687 6076
rect 28349 91 28356 155
rect 28420 91 28436 155
rect 28500 91 28516 155
rect 28580 91 28596 155
rect 28660 91 28687 155
rect 28349 0 28687 91
use invcell  invcell_0
timestamp 1656729169
transform 1 0 6097 0 1 -4063
box 8992 6886 13272 7528
use nbrhalf_32  nbrhalf_32_0
timestamp 1656729169
transform -1 0 28562 0 -1 8785
box -1666 2527 26658 5448
use nbrhalf_32  nbrhalf_32_1
timestamp 1656729169
transform 1 0 5833 0 1 -2527
box -1666 2527 26658 5448
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1656729169
transform 1 0 19407 0 1 2871
box -38 -48 130 592
use unitcell_nbr  unitcell_nbr_0
timestamp 1656729169
transform 1 0 967 0 1 1185
box -574 -1185 1322 1192
use unitcell_nbr  unitcell_nbr_1
timestamp 1656729169
transform 1 0 2855 0 1 1185
box -574 -1185 1322 1192
<< labels >>
flabel metal2 s 30621 1 30665 793 1 FreeSans 2000 0 0 0 C[31]
port 1 nsew
flabel metal2 s 28733 1 28777 793 1 FreeSans 2000 0 0 0 C[30]
port 2 nsew
flabel metal2 s 26845 1 26889 793 1 FreeSans 2000 0 0 0 C[29]
port 3 nsew
flabel metal2 s 24957 1 25001 793 1 FreeSans 2000 0 0 0 C[28]
port 4 nsew
flabel metal2 s 23069 1 23113 793 1 FreeSans 2000 0 0 0 C[27]
port 5 nsew
flabel metal2 s 21181 1 21225 793 1 FreeSans 2000 0 0 0 C[26]
port 6 nsew
flabel metal2 s 19293 1 19337 793 1 FreeSans 2000 0 0 0 C[25]
port 7 nsew
flabel metal2 s 17405 1 17449 793 1 FreeSans 2000 0 0 0 C[24]
port 8 nsew
flabel metal2 s 15517 1 15561 793 1 FreeSans 2000 0 0 0 C[23]
port 9 nsew
flabel metal2 s 13629 1 13673 793 1 FreeSans 2000 0 0 0 C[22]
port 10 nsew
flabel metal2 s 11741 1 11785 793 1 FreeSans 2000 0 0 0 C[21]
port 11 nsew
flabel metal2 s 9853 1 9897 793 1 FreeSans 2000 0 0 0 C[20]
port 12 nsew
flabel metal2 s 7965 1 8009 793 1 FreeSans 2000 0 0 0 C[19]
port 13 nsew
flabel metal2 s 6077 1 6121 793 1 FreeSans 2000 0 0 0 C[18]
port 14 nsew
flabel metal2 s 4189 1 4233 793 1 FreeSans 2000 0 0 0 C[17]
port 15 nsew
flabel metal2 s 2301 1 2345 793 1 FreeSans 2000 0 0 0 C[16]
port 16 nsew
flabel metal2 s 413 1 457 793 1 FreeSans 2000 0 0 0 C[15]
port 17 nsew
flabel metal2 s 3730 5465 3774 6257 1 FreeSans 2000 0 0 0 C[14]
port 18 nsew
flabel metal2 s 5618 5465 5662 6257 1 FreeSans 2000 0 0 0 C[13]
port 19 nsew
flabel metal2 s 7506 5465 7550 6257 1 FreeSans 2000 0 0 0 C[12]
port 20 nsew
flabel metal2 s 9394 5465 9438 6257 1 FreeSans 2000 0 0 0 C[11]
port 21 nsew
flabel metal2 s 11282 5465 11326 6257 1 FreeSans 2000 0 0 0 C[10]
port 22 nsew
flabel metal2 s 13170 5465 13214 6257 1 FreeSans 2000 0 0 0 C[9]
port 23 nsew
flabel metal2 s 15058 5465 15102 6257 1 FreeSans 2000 0 0 0 C[8]
port 24 nsew
flabel metal2 s 16946 5465 16990 6257 1 FreeSans 2000 0 0 0 C[7]
port 25 nsew
flabel metal2 s 18834 5465 18878 6257 1 FreeSans 2000 0 0 0 C[6]
port 26 nsew
flabel metal2 s 20722 5465 20766 6257 1 FreeSans 2000 0 0 0 C[5]
port 27 nsew
flabel metal2 s 22610 5465 22654 6257 1 FreeSans 2000 0 0 0 C[4]
port 28 nsew
flabel metal2 s 24498 5465 24542 6257 1 FreeSans 2000 0 0 0 C[3]
port 29 nsew
flabel metal2 s 26386 5465 26430 6257 1 FreeSans 2000 0 0 0 C[2]
port 30 nsew
flabel metal2 s 28274 5465 28318 6257 1 FreeSans 2000 0 0 0 C[1]
port 31 nsew
flabel metal2 s 30162 5465 30206 6257 1 FreeSans 2000 0 0 0 C[0]
port 32 nsew
flabel metal4 s 1915 1 2253 6259 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 5699 0 6037 6258 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 9473 1 9811 6259 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 13251 1 13589 6259 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 17019 1 17357 6259 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 20791 1 21129 6259 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 24561 1 24899 6259 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 28349 0 28687 6258 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 3813 1 4151 6257 1 FreeSans 2000 0 0 0 VDD
port 34 nsew
flabel metal4 s 7589 1 7927 6257 1 FreeSans 2000 0 0 0 VDD
port 34 nsew
flabel metal4 s 11359 1 11697 6257 1 FreeSans 2000 0 0 0 VDD
port 34 nsew
flabel metal4 s 15127 1 15465 6257 1 FreeSans 2000 0 0 0 VDD
port 34 nsew
flabel metal4 s 18899 1 19237 6257 1 FreeSans 2000 0 0 0 VDD
port 34 nsew
flabel metal4 s 22667 1 23005 6257 1 FreeSans 2000 0 0 0 VDD
port 34 nsew
flabel metal4 s 26463 1 26801 6257 1 FreeSans 2000 0 0 0 VDD
port 34 nsew
flabel metal3 s 18 3036 554 3129 1 FreeSans 1000 0 0 0 RESET
port 35 nsew
flabel metal1 s 32393 782 32622 859 1 FreeSans 1000 0 0 0 OUT
port 36 nsew
<< properties >>
string GDS_END 9106022
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/merge/design_merged.gds
string GDS_START 9075298
<< end >>
