magic
tech sky130A
magscale 1 2
timestamp 1655322987
<< nwell >>
rect 15071 3413 15595 3591
<< pwell >>
rect 9509 3441 9739 3559
rect 24547 3445 24775 3571
<< psubdiff >>
rect 9535 3517 9713 3533
rect 24573 3525 24749 3545
rect 9535 3483 9573 3517
rect 9607 3483 9641 3517
rect 9675 3483 9713 3517
rect 9535 3467 9713 3483
rect 24573 3491 24610 3525
rect 24644 3491 24678 3525
rect 24712 3491 24749 3525
rect 24573 3471 24749 3491
<< nsubdiff >>
rect 15163 3508 15371 3525
rect 15163 3474 15216 3508
rect 15250 3474 15284 3508
rect 15318 3474 15371 3508
rect 15163 3457 15371 3474
<< psubdiffcont >>
rect 9573 3483 9607 3517
rect 9641 3483 9675 3517
rect 24610 3491 24644 3525
rect 24678 3491 24712 3525
<< nsubdiffcont >>
rect 15216 3474 15250 3508
rect 15284 3474 15318 3508
<< locali >>
rect 9407 3517 9705 3533
rect 24581 3532 24741 3545
rect 24502 3525 24741 3532
rect 9407 3483 9573 3517
rect 9607 3483 9641 3517
rect 9675 3483 9705 3517
rect 9407 3467 9705 3483
rect 15171 3508 15363 3525
rect 15171 3474 15216 3508
rect 15250 3474 15284 3508
rect 15318 3474 15363 3508
rect 24502 3491 24610 3525
rect 24644 3491 24678 3525
rect 24712 3491 24741 3525
rect 24502 3488 24741 3491
rect 15171 3429 15363 3474
rect 24581 3471 24741 3488
rect 15241 3213 15279 3217
rect 15241 3179 15243 3213
rect 15277 3179 15279 3213
rect 15241 3175 15279 3179
rect 16597 3126 16643 3129
rect 16597 3092 16603 3126
rect 16637 3092 16643 3126
rect 16597 3089 16643 3092
<< viali >>
rect 15243 3179 15277 3213
rect 16603 3092 16637 3126
rect 19142 3088 19176 3122
<< metal1 >>
rect 22891 3645 22951 3677
rect 9755 3642 11014 3643
rect 9755 3597 11485 3642
rect 9378 3275 10152 3352
rect 9378 3159 9467 3275
rect 9775 3159 10152 3275
rect 9378 2898 10152 3159
rect 11425 3161 11485 3597
rect 22891 3599 24632 3645
rect 15149 3441 15393 3459
rect 15149 3389 15181 3441
rect 15233 3389 15245 3441
rect 15297 3389 15309 3441
rect 15361 3389 15393 3441
rect 15149 3371 15393 3389
rect 18915 3453 19159 3461
rect 18915 3443 19183 3453
rect 18915 3391 18947 3443
rect 18999 3391 19011 3443
rect 19063 3391 19075 3443
rect 19127 3391 19183 3443
rect 18915 3381 19183 3391
rect 18915 3373 19159 3381
rect 19195 3367 19395 3463
rect 15235 3213 15291 3229
rect 15235 3179 15243 3213
rect 15277 3179 15291 3213
rect 15235 3161 15291 3179
rect 11425 3101 15291 3161
rect 16581 3135 16655 3145
rect 11425 2660 11485 3101
rect 16581 3083 16593 3135
rect 16645 3083 16655 3135
rect 16581 3077 16655 3083
rect 19130 3135 19212 3146
rect 22891 3135 22951 3599
rect 19130 3122 22951 3135
rect 19130 3088 19142 3122
rect 19176 3088 22951 3122
rect 19130 3075 22951 3088
rect 19130 3064 19212 3075
rect 17013 2899 17297 2917
rect 17013 2847 17033 2899
rect 17085 2847 17097 2899
rect 17149 2847 17161 2899
rect 17213 2847 17225 2899
rect 17277 2847 17297 2899
rect 17013 2829 17297 2847
rect 19201 2823 19401 2919
rect 10746 2604 11485 2660
rect 22891 2661 22951 3075
rect 24432 3317 25188 3374
rect 24432 3201 24555 3317
rect 24863 3201 25188 3317
rect 24432 2880 25188 3201
rect 22891 2615 24742 2661
rect 22891 2583 22951 2615
rect 32375 782 32604 859
<< via1 >>
rect 9467 3159 9775 3275
rect 15181 3389 15233 3441
rect 15245 3389 15297 3441
rect 15309 3389 15361 3441
rect 18947 3391 18999 3443
rect 19011 3391 19063 3443
rect 19075 3391 19127 3443
rect 16593 3126 16645 3135
rect 16593 3092 16603 3126
rect 16603 3092 16637 3126
rect 16637 3092 16645 3126
rect 16593 3083 16645 3092
rect 17033 2847 17085 2899
rect 17097 2847 17149 2899
rect 17161 2847 17213 2899
rect 17225 2847 17277 2899
rect 24555 3201 24863 3317
<< metal2 >>
rect 3712 5465 3756 6257
rect 5600 5465 5644 6257
rect 7488 5465 7532 6257
rect 9376 5465 9420 6257
rect 11264 5465 11308 6257
rect 13152 5465 13196 6257
rect 15040 5465 15084 6257
rect 16928 5465 16972 6257
rect 18816 5465 18860 6257
rect 20704 5465 20748 6257
rect 22592 5465 22636 6257
rect 24480 5465 24524 6257
rect 26368 5465 26412 6257
rect 28256 5465 28300 6257
rect 30144 5465 30188 6257
rect 151 4747 1941 4783
rect 30159 4747 32649 4783
rect 151 1511 187 4747
rect 15159 3443 15383 3469
rect 15159 3387 15163 3443
rect 15219 3441 15243 3443
rect 15299 3441 15323 3443
rect 15233 3389 15243 3441
rect 15299 3389 15309 3441
rect 15219 3387 15243 3389
rect 15299 3387 15323 3389
rect 15379 3387 15383 3443
rect 15159 3361 15383 3387
rect 18925 3445 19149 3471
rect 18925 3389 18929 3445
rect 18985 3443 19009 3445
rect 19065 3443 19089 3445
rect 18999 3391 19009 3443
rect 19065 3391 19075 3443
rect 18985 3389 19009 3391
rect 19065 3389 19089 3391
rect 19145 3389 19149 3445
rect 18925 3363 19149 3389
rect 24555 3317 24863 3327
rect 9467 3275 9775 3285
rect 24555 3191 24863 3201
rect 9467 3149 9775 3159
rect 16587 3135 16651 3145
rect 411 3111 551 3131
rect 411 3055 445 3111
rect 501 3103 551 3111
rect 16587 3103 16593 3135
rect 501 3083 16593 3103
rect 16645 3083 16651 3135
rect 501 3071 16651 3083
rect 501 3055 551 3071
rect 411 3035 551 3055
rect 17023 2901 17287 2927
rect 17023 2899 17047 2901
rect 17103 2899 17127 2901
rect 17183 2899 17207 2901
rect 17263 2899 17287 2901
rect 17023 2847 17033 2899
rect 17277 2847 17287 2899
rect 17023 2845 17047 2847
rect 17103 2845 17127 2847
rect 17183 2845 17207 2847
rect 17263 2845 17287 2847
rect 17023 2819 17287 2845
rect 595 2555 1621 2556
rect 2485 2555 3511 2556
rect 375 2367 4337 2555
rect 595 2110 1621 2367
rect 2485 2110 3511 2367
rect 375 2001 4258 2110
rect 32613 1511 32649 4747
rect 151 1475 419 1511
rect 32399 1475 32651 1511
rect 395 1 439 793
rect 2283 1 2327 793
rect 4171 1 4215 793
rect 6059 1 6103 793
rect 7947 1 7991 793
rect 9835 1 9879 793
rect 11723 1 11767 793
rect 13611 1 13655 793
rect 15499 1 15543 793
rect 17387 1 17431 793
rect 19275 1 19319 793
rect 21163 1 21207 793
rect 23051 1 23095 793
rect 24939 1 24983 793
rect 26827 1 26871 793
rect 28715 1 28759 793
rect 30603 1 30647 793
<< via2 >>
rect 15163 3441 15219 3443
rect 15243 3441 15299 3443
rect 15323 3441 15379 3443
rect 15163 3389 15181 3441
rect 15181 3389 15219 3441
rect 15243 3389 15245 3441
rect 15245 3389 15297 3441
rect 15297 3389 15299 3441
rect 15323 3389 15361 3441
rect 15361 3389 15379 3441
rect 15163 3387 15219 3389
rect 15243 3387 15299 3389
rect 15323 3387 15379 3389
rect 18929 3443 18985 3445
rect 19009 3443 19065 3445
rect 19089 3443 19145 3445
rect 18929 3391 18947 3443
rect 18947 3391 18985 3443
rect 19009 3391 19011 3443
rect 19011 3391 19063 3443
rect 19063 3391 19065 3443
rect 19089 3391 19127 3443
rect 19127 3391 19145 3443
rect 18929 3389 18985 3391
rect 19009 3389 19065 3391
rect 19089 3389 19145 3391
rect 9473 3189 9529 3245
rect 9553 3189 9609 3245
rect 9633 3189 9689 3245
rect 9713 3189 9769 3245
rect 24561 3231 24617 3287
rect 24641 3231 24697 3287
rect 24721 3231 24777 3287
rect 24801 3231 24857 3287
rect 445 3055 501 3111
rect 17047 2899 17103 2901
rect 17127 2899 17183 2901
rect 17207 2899 17263 2901
rect 17047 2847 17085 2899
rect 17085 2847 17097 2899
rect 17097 2847 17103 2899
rect 17127 2847 17149 2899
rect 17149 2847 17161 2899
rect 17161 2847 17183 2899
rect 17207 2847 17213 2899
rect 17213 2847 17225 2899
rect 17225 2847 17263 2899
rect 17047 2845 17103 2847
rect 17127 2845 17183 2847
rect 17207 2845 17263 2847
<< metal3 >>
rect 1930 6167 2258 6193
rect 1930 6103 1942 6167
rect 2006 6103 2022 6167
rect 2086 6103 2102 6167
rect 2166 6103 2182 6167
rect 2246 6103 2258 6167
rect 1930 6077 2258 6103
rect 5706 6167 6034 6193
rect 5706 6103 5718 6167
rect 5782 6103 5798 6167
rect 5862 6103 5878 6167
rect 5942 6103 5958 6167
rect 6022 6103 6034 6167
rect 5706 6077 6034 6103
rect 9482 6167 9810 6193
rect 9482 6103 9494 6167
rect 9558 6103 9574 6167
rect 9638 6103 9654 6167
rect 9718 6103 9734 6167
rect 9798 6103 9810 6167
rect 9482 6077 9810 6103
rect 13258 6167 13586 6193
rect 13258 6103 13270 6167
rect 13334 6103 13350 6167
rect 13414 6103 13430 6167
rect 13494 6103 13510 6167
rect 13574 6103 13586 6167
rect 13258 6077 13586 6103
rect 17028 6167 17356 6193
rect 17028 6103 17040 6167
rect 17104 6103 17120 6167
rect 17184 6103 17200 6167
rect 17264 6103 17280 6167
rect 17344 6103 17356 6167
rect 17028 6077 17356 6103
rect 20804 6167 21132 6193
rect 20804 6103 20816 6167
rect 20880 6103 20896 6167
rect 20960 6103 20976 6167
rect 21040 6103 21056 6167
rect 21120 6103 21132 6167
rect 20804 6077 21132 6103
rect 24580 6167 24908 6193
rect 24580 6103 24592 6167
rect 24656 6103 24672 6167
rect 24736 6103 24752 6167
rect 24816 6103 24832 6167
rect 24896 6103 24908 6167
rect 24580 6077 24908 6103
rect 28356 6167 28684 6193
rect 28356 6103 28368 6167
rect 28432 6103 28448 6167
rect 28512 6103 28528 6167
rect 28592 6103 28608 6167
rect 28672 6103 28684 6167
rect 28356 6077 28684 6103
rect 3818 4043 4146 4069
rect 3818 3979 3830 4043
rect 3894 3979 3910 4043
rect 3974 3979 3990 4043
rect 4054 3979 4070 4043
rect 4134 3979 4146 4043
rect 3818 3953 4146 3979
rect 7594 4043 7922 4069
rect 7594 3979 7606 4043
rect 7670 3979 7686 4043
rect 7750 3979 7766 4043
rect 7830 3979 7846 4043
rect 7910 3979 7922 4043
rect 7594 3953 7922 3979
rect 11370 4043 11698 4069
rect 11370 3979 11382 4043
rect 11446 3979 11462 4043
rect 11526 3979 11542 4043
rect 11606 3979 11622 4043
rect 11686 3979 11698 4043
rect 11370 3953 11698 3979
rect 15146 4043 15474 4069
rect 15146 3979 15158 4043
rect 15222 3979 15238 4043
rect 15302 3979 15318 4043
rect 15382 3979 15398 4043
rect 15462 3979 15474 4043
rect 15146 3953 15474 3979
rect 18916 4043 19244 4069
rect 18916 3979 18928 4043
rect 18992 3979 19008 4043
rect 19072 3979 19088 4043
rect 19152 3979 19168 4043
rect 19232 3979 19244 4043
rect 18916 3953 19244 3979
rect 22692 4043 23020 4069
rect 22692 3979 22704 4043
rect 22768 3979 22784 4043
rect 22848 3979 22864 4043
rect 22928 3979 22944 4043
rect 23008 3979 23020 4043
rect 22692 3953 23020 3979
rect 26468 4043 26796 4069
rect 26468 3979 26480 4043
rect 26544 3979 26560 4043
rect 26624 3979 26640 4043
rect 26704 3979 26720 4043
rect 26784 3979 26796 4043
rect 26468 3953 26796 3979
rect 15149 3447 15393 3464
rect 15149 3383 15159 3447
rect 15223 3383 15239 3447
rect 15303 3383 15319 3447
rect 15383 3383 15393 3447
rect 15149 3366 15393 3383
rect 18915 3449 19159 3466
rect 18915 3385 18925 3449
rect 18989 3385 19005 3449
rect 19069 3385 19085 3449
rect 19149 3385 19159 3449
rect 18915 3368 19159 3385
rect 24545 3291 24873 3322
rect 9457 3249 9785 3280
rect 9457 3185 9469 3249
rect 9533 3185 9549 3249
rect 9613 3185 9629 3249
rect 9693 3185 9709 3249
rect 9773 3185 9785 3249
rect 24545 3227 24557 3291
rect 24621 3227 24637 3291
rect 24701 3227 24717 3291
rect 24781 3227 24797 3291
rect 24861 3227 24873 3291
rect 24545 3196 24873 3227
rect 9457 3154 9785 3185
rect 0 3111 536 3129
rect 0 3055 445 3111
rect 501 3055 536 3111
rect 0 3036 536 3055
rect 17013 2905 17297 2922
rect 17013 2841 17043 2905
rect 17107 2841 17123 2905
rect 17187 2841 17203 2905
rect 17267 2841 17297 2905
rect 17013 2824 17297 2841
rect 3788 2279 4116 2305
rect 3788 2215 3800 2279
rect 3864 2215 3880 2279
rect 3944 2215 3960 2279
rect 4024 2215 4040 2279
rect 4104 2215 4116 2279
rect 3788 2189 4116 2215
rect 7564 2279 7892 2305
rect 7564 2215 7576 2279
rect 7640 2215 7656 2279
rect 7720 2215 7736 2279
rect 7800 2215 7816 2279
rect 7880 2215 7892 2279
rect 7564 2189 7892 2215
rect 11340 2279 11668 2305
rect 11340 2215 11352 2279
rect 11416 2215 11432 2279
rect 11496 2215 11512 2279
rect 11576 2215 11592 2279
rect 11656 2215 11668 2279
rect 11340 2189 11668 2215
rect 15116 2279 15444 2305
rect 15116 2215 15128 2279
rect 15192 2215 15208 2279
rect 15272 2215 15288 2279
rect 15352 2215 15368 2279
rect 15432 2215 15444 2279
rect 15116 2189 15444 2215
rect 18886 2279 19214 2305
rect 18886 2215 18898 2279
rect 18962 2215 18978 2279
rect 19042 2215 19058 2279
rect 19122 2215 19138 2279
rect 19202 2215 19214 2279
rect 18886 2189 19214 2215
rect 22662 2279 22990 2305
rect 22662 2215 22674 2279
rect 22738 2215 22754 2279
rect 22818 2215 22834 2279
rect 22898 2215 22914 2279
rect 22978 2215 22990 2279
rect 22662 2189 22990 2215
rect 26438 2279 26766 2305
rect 26438 2215 26450 2279
rect 26514 2215 26530 2279
rect 26594 2215 26610 2279
rect 26674 2215 26690 2279
rect 26754 2215 26766 2279
rect 26438 2189 26766 2215
rect 1900 155 2228 181
rect 1900 91 1912 155
rect 1976 91 1992 155
rect 2056 91 2072 155
rect 2136 91 2152 155
rect 2216 91 2228 155
rect 1900 65 2228 91
rect 5676 155 6004 181
rect 5676 91 5688 155
rect 5752 91 5768 155
rect 5832 91 5848 155
rect 5912 91 5928 155
rect 5992 91 6004 155
rect 5676 65 6004 91
rect 9452 155 9780 181
rect 9452 91 9464 155
rect 9528 91 9544 155
rect 9608 91 9624 155
rect 9688 91 9704 155
rect 9768 91 9780 155
rect 9452 65 9780 91
rect 13228 155 13556 181
rect 13228 91 13240 155
rect 13304 91 13320 155
rect 13384 91 13400 155
rect 13464 91 13480 155
rect 13544 91 13556 155
rect 13228 65 13556 91
rect 17004 155 17332 181
rect 17004 91 17016 155
rect 17080 91 17096 155
rect 17160 91 17176 155
rect 17240 91 17256 155
rect 17320 91 17332 155
rect 17004 65 17332 91
rect 20774 155 21102 181
rect 20774 91 20786 155
rect 20850 91 20866 155
rect 20930 91 20946 155
rect 21010 91 21026 155
rect 21090 91 21102 155
rect 20774 65 21102 91
rect 24550 155 24878 181
rect 24550 91 24562 155
rect 24626 91 24642 155
rect 24706 91 24722 155
rect 24786 91 24802 155
rect 24866 91 24878 155
rect 24550 65 24878 91
rect 28326 155 28654 181
rect 28326 91 28338 155
rect 28402 91 28418 155
rect 28482 91 28498 155
rect 28562 91 28578 155
rect 28642 91 28654 155
rect 28326 65 28654 91
<< via3 >>
rect 1942 6103 2006 6167
rect 2022 6103 2086 6167
rect 2102 6103 2166 6167
rect 2182 6103 2246 6167
rect 5718 6103 5782 6167
rect 5798 6103 5862 6167
rect 5878 6103 5942 6167
rect 5958 6103 6022 6167
rect 9494 6103 9558 6167
rect 9574 6103 9638 6167
rect 9654 6103 9718 6167
rect 9734 6103 9798 6167
rect 13270 6103 13334 6167
rect 13350 6103 13414 6167
rect 13430 6103 13494 6167
rect 13510 6103 13574 6167
rect 17040 6103 17104 6167
rect 17120 6103 17184 6167
rect 17200 6103 17264 6167
rect 17280 6103 17344 6167
rect 20816 6103 20880 6167
rect 20896 6103 20960 6167
rect 20976 6103 21040 6167
rect 21056 6103 21120 6167
rect 24592 6103 24656 6167
rect 24672 6103 24736 6167
rect 24752 6103 24816 6167
rect 24832 6103 24896 6167
rect 28368 6103 28432 6167
rect 28448 6103 28512 6167
rect 28528 6103 28592 6167
rect 28608 6103 28672 6167
rect 3830 3979 3894 4043
rect 3910 3979 3974 4043
rect 3990 3979 4054 4043
rect 4070 3979 4134 4043
rect 7606 3979 7670 4043
rect 7686 3979 7750 4043
rect 7766 3979 7830 4043
rect 7846 3979 7910 4043
rect 11382 3979 11446 4043
rect 11462 3979 11526 4043
rect 11542 3979 11606 4043
rect 11622 3979 11686 4043
rect 15158 3979 15222 4043
rect 15238 3979 15302 4043
rect 15318 3979 15382 4043
rect 15398 3979 15462 4043
rect 18928 3979 18992 4043
rect 19008 3979 19072 4043
rect 19088 3979 19152 4043
rect 19168 3979 19232 4043
rect 22704 3979 22768 4043
rect 22784 3979 22848 4043
rect 22864 3979 22928 4043
rect 22944 3979 23008 4043
rect 26480 3979 26544 4043
rect 26560 3979 26624 4043
rect 26640 3979 26704 4043
rect 26720 3979 26784 4043
rect 15159 3443 15223 3447
rect 15159 3387 15163 3443
rect 15163 3387 15219 3443
rect 15219 3387 15223 3443
rect 15159 3383 15223 3387
rect 15239 3443 15303 3447
rect 15239 3387 15243 3443
rect 15243 3387 15299 3443
rect 15299 3387 15303 3443
rect 15239 3383 15303 3387
rect 15319 3443 15383 3447
rect 15319 3387 15323 3443
rect 15323 3387 15379 3443
rect 15379 3387 15383 3443
rect 15319 3383 15383 3387
rect 18925 3445 18989 3449
rect 18925 3389 18929 3445
rect 18929 3389 18985 3445
rect 18985 3389 18989 3445
rect 18925 3385 18989 3389
rect 19005 3445 19069 3449
rect 19005 3389 19009 3445
rect 19009 3389 19065 3445
rect 19065 3389 19069 3445
rect 19005 3385 19069 3389
rect 19085 3445 19149 3449
rect 19085 3389 19089 3445
rect 19089 3389 19145 3445
rect 19145 3389 19149 3445
rect 19085 3385 19149 3389
rect 9469 3245 9533 3249
rect 9469 3189 9473 3245
rect 9473 3189 9529 3245
rect 9529 3189 9533 3245
rect 9469 3185 9533 3189
rect 9549 3245 9613 3249
rect 9549 3189 9553 3245
rect 9553 3189 9609 3245
rect 9609 3189 9613 3245
rect 9549 3185 9613 3189
rect 9629 3245 9693 3249
rect 9629 3189 9633 3245
rect 9633 3189 9689 3245
rect 9689 3189 9693 3245
rect 9629 3185 9693 3189
rect 9709 3245 9773 3249
rect 9709 3189 9713 3245
rect 9713 3189 9769 3245
rect 9769 3189 9773 3245
rect 9709 3185 9773 3189
rect 24557 3287 24621 3291
rect 24557 3231 24561 3287
rect 24561 3231 24617 3287
rect 24617 3231 24621 3287
rect 24557 3227 24621 3231
rect 24637 3287 24701 3291
rect 24637 3231 24641 3287
rect 24641 3231 24697 3287
rect 24697 3231 24701 3287
rect 24637 3227 24701 3231
rect 24717 3287 24781 3291
rect 24717 3231 24721 3287
rect 24721 3231 24777 3287
rect 24777 3231 24781 3287
rect 24717 3227 24781 3231
rect 24797 3287 24861 3291
rect 24797 3231 24801 3287
rect 24801 3231 24857 3287
rect 24857 3231 24861 3287
rect 24797 3227 24861 3231
rect 17043 2901 17107 2905
rect 17043 2845 17047 2901
rect 17047 2845 17103 2901
rect 17103 2845 17107 2901
rect 17043 2841 17107 2845
rect 17123 2901 17187 2905
rect 17123 2845 17127 2901
rect 17127 2845 17183 2901
rect 17183 2845 17187 2901
rect 17123 2841 17187 2845
rect 17203 2901 17267 2905
rect 17203 2845 17207 2901
rect 17207 2845 17263 2901
rect 17263 2845 17267 2901
rect 17203 2841 17267 2845
rect 3800 2215 3864 2279
rect 3880 2215 3944 2279
rect 3960 2215 4024 2279
rect 4040 2215 4104 2279
rect 7576 2215 7640 2279
rect 7656 2215 7720 2279
rect 7736 2215 7800 2279
rect 7816 2215 7880 2279
rect 11352 2215 11416 2279
rect 11432 2215 11496 2279
rect 11512 2215 11576 2279
rect 11592 2215 11656 2279
rect 15128 2215 15192 2279
rect 15208 2215 15272 2279
rect 15288 2215 15352 2279
rect 15368 2215 15432 2279
rect 18898 2215 18962 2279
rect 18978 2215 19042 2279
rect 19058 2215 19122 2279
rect 19138 2215 19202 2279
rect 22674 2215 22738 2279
rect 22754 2215 22818 2279
rect 22834 2215 22898 2279
rect 22914 2215 22978 2279
rect 26450 2215 26514 2279
rect 26530 2215 26594 2279
rect 26610 2215 26674 2279
rect 26690 2215 26754 2279
rect 1912 91 1976 155
rect 1992 91 2056 155
rect 2072 91 2136 155
rect 2152 91 2216 155
rect 5688 91 5752 155
rect 5768 91 5832 155
rect 5848 91 5912 155
rect 5928 91 5992 155
rect 9464 91 9528 155
rect 9544 91 9608 155
rect 9624 91 9688 155
rect 9704 91 9768 155
rect 13240 91 13304 155
rect 13320 91 13384 155
rect 13400 91 13464 155
rect 13480 91 13544 155
rect 17016 91 17080 155
rect 17096 91 17160 155
rect 17176 91 17240 155
rect 17256 91 17320 155
rect 20786 91 20850 155
rect 20866 91 20930 155
rect 20946 91 21010 155
rect 21026 91 21090 155
rect 24562 91 24626 155
rect 24642 91 24706 155
rect 24722 91 24786 155
rect 24802 91 24866 155
rect 28338 91 28402 155
rect 28418 91 28482 155
rect 28498 91 28562 155
rect 28578 91 28642 155
<< metal4 >>
rect 1897 6194 2235 6259
rect 1897 6167 2249 6194
rect 1897 6103 1942 6167
rect 2006 6103 2022 6167
rect 2086 6103 2102 6167
rect 2166 6103 2182 6167
rect 2246 6103 2249 6167
rect 1897 6076 2249 6103
rect 1897 155 2235 6076
rect 1897 91 1912 155
rect 1976 91 1992 155
rect 2056 91 2072 155
rect 2136 91 2152 155
rect 2216 91 2235 155
rect 1897 1 2235 91
rect 3795 4070 4133 6257
rect 5681 6194 6019 6258
rect 5681 6167 6025 6194
rect 5681 6103 5718 6167
rect 5782 6103 5798 6167
rect 5862 6103 5878 6167
rect 5942 6103 5958 6167
rect 6022 6103 6025 6167
rect 5681 6076 6025 6103
rect 3795 4043 4137 4070
rect 3795 3979 3830 4043
rect 3894 3979 3910 4043
rect 3974 3979 3990 4043
rect 4054 3979 4070 4043
rect 4134 3979 4137 4043
rect 3795 3952 4137 3979
rect 3795 2279 4133 3952
rect 3795 2215 3800 2279
rect 3864 2215 3880 2279
rect 3944 2215 3960 2279
rect 4024 2215 4040 2279
rect 4104 2215 4133 2279
rect 3795 1 4133 2215
rect 5681 155 6019 6076
rect 5681 91 5688 155
rect 5752 91 5768 155
rect 5832 91 5848 155
rect 5912 91 5928 155
rect 5992 91 6019 155
rect 5681 0 6019 91
rect 7571 4070 7909 6257
rect 9455 6194 9793 6259
rect 9455 6167 9801 6194
rect 9455 6103 9494 6167
rect 9558 6103 9574 6167
rect 9638 6103 9654 6167
rect 9718 6103 9734 6167
rect 9798 6103 9801 6167
rect 9455 6076 9801 6103
rect 7571 4043 7913 4070
rect 7571 3979 7606 4043
rect 7670 3979 7686 4043
rect 7750 3979 7766 4043
rect 7830 3979 7846 4043
rect 7910 3979 7913 4043
rect 7571 3952 7913 3979
rect 7571 2279 7909 3952
rect 7571 2215 7576 2279
rect 7640 2215 7656 2279
rect 7720 2215 7736 2279
rect 7800 2215 7816 2279
rect 7880 2215 7909 2279
rect 7571 1 7909 2215
rect 9455 3249 9793 6076
rect 9455 3185 9469 3249
rect 9533 3185 9549 3249
rect 9613 3185 9629 3249
rect 9693 3185 9709 3249
rect 9773 3185 9793 3249
rect 9455 155 9793 3185
rect 9455 91 9464 155
rect 9528 91 9544 155
rect 9608 91 9624 155
rect 9688 91 9704 155
rect 9768 91 9793 155
rect 9455 1 9793 91
rect 11341 4070 11679 6257
rect 13233 6194 13571 6259
rect 13233 6167 13577 6194
rect 13233 6103 13270 6167
rect 13334 6103 13350 6167
rect 13414 6103 13430 6167
rect 13494 6103 13510 6167
rect 13574 6103 13577 6167
rect 13233 6076 13577 6103
rect 11341 4043 11689 4070
rect 11341 3979 11382 4043
rect 11446 3979 11462 4043
rect 11526 3979 11542 4043
rect 11606 3979 11622 4043
rect 11686 3979 11689 4043
rect 11341 3952 11689 3979
rect 11341 2279 11679 3952
rect 11341 2215 11352 2279
rect 11416 2215 11432 2279
rect 11496 2215 11512 2279
rect 11576 2215 11592 2279
rect 11656 2215 11679 2279
rect 11341 1 11679 2215
rect 13233 155 13571 6076
rect 13233 91 13240 155
rect 13304 91 13320 155
rect 13384 91 13400 155
rect 13464 91 13480 155
rect 13544 91 13571 155
rect 13233 1 13571 91
rect 15109 4070 15447 6257
rect 17001 6194 17339 6259
rect 17001 6167 17347 6194
rect 17001 6103 17040 6167
rect 17104 6103 17120 6167
rect 17184 6103 17200 6167
rect 17264 6103 17280 6167
rect 17344 6103 17347 6167
rect 17001 6076 17347 6103
rect 15109 4043 15465 4070
rect 15109 3979 15158 4043
rect 15222 3979 15238 4043
rect 15302 3979 15318 4043
rect 15382 3979 15398 4043
rect 15462 3979 15465 4043
rect 15109 3952 15465 3979
rect 15109 3447 15447 3952
rect 15109 3383 15159 3447
rect 15223 3383 15239 3447
rect 15303 3383 15319 3447
rect 15383 3383 15447 3447
rect 15109 2279 15447 3383
rect 15109 2215 15128 2279
rect 15192 2215 15208 2279
rect 15272 2215 15288 2279
rect 15352 2215 15368 2279
rect 15432 2215 15447 2279
rect 15109 1 15447 2215
rect 17001 2905 17339 6076
rect 17001 2841 17043 2905
rect 17107 2841 17123 2905
rect 17187 2841 17203 2905
rect 17267 2841 17339 2905
rect 17001 155 17339 2841
rect 17001 91 17016 155
rect 17080 91 17096 155
rect 17160 91 17176 155
rect 17240 91 17256 155
rect 17320 91 17339 155
rect 17001 1 17339 91
rect 18881 4070 19219 6257
rect 20773 6194 21111 6259
rect 20773 6167 21123 6194
rect 20773 6103 20816 6167
rect 20880 6103 20896 6167
rect 20960 6103 20976 6167
rect 21040 6103 21056 6167
rect 21120 6103 21123 6167
rect 20773 6076 21123 6103
rect 18881 4043 19235 4070
rect 18881 3979 18928 4043
rect 18992 3979 19008 4043
rect 19072 3979 19088 4043
rect 19152 3979 19168 4043
rect 19232 3979 19235 4043
rect 18881 3952 19235 3979
rect 18881 3449 19219 3952
rect 18881 3385 18925 3449
rect 18989 3385 19005 3449
rect 19069 3385 19085 3449
rect 19149 3385 19219 3449
rect 18881 2279 19219 3385
rect 18881 2215 18898 2279
rect 18962 2215 18978 2279
rect 19042 2215 19058 2279
rect 19122 2215 19138 2279
rect 19202 2215 19219 2279
rect 18881 1 19219 2215
rect 20773 155 21111 6076
rect 20773 91 20786 155
rect 20850 91 20866 155
rect 20930 91 20946 155
rect 21010 91 21026 155
rect 21090 91 21111 155
rect 20773 1 21111 91
rect 22649 4070 22987 6257
rect 24543 6194 24881 6259
rect 24543 6167 24899 6194
rect 24543 6103 24592 6167
rect 24656 6103 24672 6167
rect 24736 6103 24752 6167
rect 24816 6103 24832 6167
rect 24896 6103 24899 6167
rect 24543 6076 24899 6103
rect 22649 4043 23011 4070
rect 22649 3979 22704 4043
rect 22768 3979 22784 4043
rect 22848 3979 22864 4043
rect 22928 3979 22944 4043
rect 23008 3979 23011 4043
rect 22649 3952 23011 3979
rect 22649 2279 22987 3952
rect 22649 2215 22674 2279
rect 22738 2215 22754 2279
rect 22818 2215 22834 2279
rect 22898 2215 22914 2279
rect 22978 2215 22987 2279
rect 22649 1 22987 2215
rect 24543 3291 24881 6076
rect 24543 3227 24557 3291
rect 24621 3227 24637 3291
rect 24701 3227 24717 3291
rect 24781 3227 24797 3291
rect 24861 3227 24881 3291
rect 24543 155 24881 3227
rect 24543 91 24562 155
rect 24626 91 24642 155
rect 24706 91 24722 155
rect 24786 91 24802 155
rect 24866 91 24881 155
rect 24543 1 24881 91
rect 26445 4070 26783 6257
rect 28331 6194 28669 6258
rect 28331 6167 28675 6194
rect 28331 6103 28368 6167
rect 28432 6103 28448 6167
rect 28512 6103 28528 6167
rect 28592 6103 28608 6167
rect 28672 6103 28675 6167
rect 28331 6076 28675 6103
rect 26445 4043 26787 4070
rect 26445 3979 26480 4043
rect 26544 3979 26560 4043
rect 26624 3979 26640 4043
rect 26704 3979 26720 4043
rect 26784 3979 26787 4043
rect 26445 3952 26787 3979
rect 26445 2279 26783 3952
rect 26445 2215 26450 2279
rect 26514 2215 26530 2279
rect 26594 2215 26610 2279
rect 26674 2215 26690 2279
rect 26754 2215 26783 2279
rect 26445 1 26783 2215
rect 28331 155 28669 6076
rect 28331 91 28338 155
rect 28402 91 28418 155
rect 28482 91 28498 155
rect 28562 91 28578 155
rect 28642 91 28669 155
rect 28331 0 28669 91
use brbufhalf_32  brbufhalf_32_0
timestamp 1655322987
transform 1 0 5815 0 1 -2527
box -1666 2527 26658 5448
use brbufhalf_32  brbufhalf_32_1
timestamp 1655322987
transform -1 0 28544 0 -1 8785
box -1666 2527 26658 5448
use invcell  invcell_0
timestamp 1655322987
transform 1 0 6079 0 1 -4063
box 8992 6886 13272 7528
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1655322987
transform 1 0 19389 0 1 2871
box -38 -48 130 592
use unitcell2buf_32  unitcell2buf_32_0
timestamp 1655322987
transform 1 0 949 0 1 1185
box -574 -1185 1322 1192
use unitcell2buf_32  unitcell2buf_32_1
timestamp 1655322987
transform 1 0 2837 0 1 1185
box -574 -1185 1322 1192
<< labels >>
flabel metal2 s 30603 1 30647 793 1 FreeSans 2000 0 0 0 C[31]
port 1 nsew
flabel metal2 s 28715 1 28759 793 1 FreeSans 2000 0 0 0 C[30]
port 2 nsew
flabel metal2 s 26827 1 26871 793 1 FreeSans 2000 0 0 0 C[29]
port 3 nsew
flabel metal2 s 24939 1 24983 793 1 FreeSans 2000 0 0 0 C[28]
port 4 nsew
flabel metal2 s 23051 1 23095 793 1 FreeSans 2000 0 0 0 C[27]
port 5 nsew
flabel metal2 s 21163 1 21207 793 1 FreeSans 2000 0 0 0 C[26]
port 6 nsew
flabel metal2 s 19275 1 19319 793 1 FreeSans 2000 0 0 0 C[25]
port 7 nsew
flabel metal2 s 17387 1 17431 793 1 FreeSans 2000 0 0 0 C[24]
port 8 nsew
flabel metal2 s 15499 1 15543 793 1 FreeSans 2000 0 0 0 C[23]
port 9 nsew
flabel metal2 s 13611 1 13655 793 1 FreeSans 2000 0 0 0 C[22]
port 10 nsew
flabel metal2 s 11723 1 11767 793 1 FreeSans 2000 0 0 0 C[21]
port 11 nsew
flabel metal2 s 9835 1 9879 793 1 FreeSans 2000 0 0 0 C[20]
port 12 nsew
flabel metal2 s 7947 1 7991 793 1 FreeSans 2000 0 0 0 C[19]
port 13 nsew
flabel metal2 s 6059 1 6103 793 1 FreeSans 2000 0 0 0 C[18]
port 14 nsew
flabel metal2 s 4171 1 4215 793 1 FreeSans 2000 0 0 0 C[17]
port 15 nsew
flabel metal2 s 2283 1 2327 793 1 FreeSans 2000 0 0 0 C[16]
port 16 nsew
flabel metal2 s 395 1 439 793 1 FreeSans 2000 0 0 0 C[15]
port 17 nsew
flabel metal2 s 3712 5465 3756 6257 1 FreeSans 2000 0 0 0 C[14]
port 18 nsew
flabel metal2 s 5600 5465 5644 6257 1 FreeSans 2000 0 0 0 C[13]
port 19 nsew
flabel metal2 s 7488 5465 7532 6257 1 FreeSans 2000 0 0 0 C[12]
port 20 nsew
flabel metal2 s 9376 5465 9420 6257 1 FreeSans 2000 0 0 0 C[11]
port 21 nsew
flabel metal2 s 11264 5465 11308 6257 1 FreeSans 2000 0 0 0 C[10]
port 22 nsew
flabel metal2 s 13152 5465 13196 6257 1 FreeSans 2000 0 0 0 C[9]
port 23 nsew
flabel metal2 s 15040 5465 15084 6257 1 FreeSans 2000 0 0 0 C[8]
port 24 nsew
flabel metal2 s 16928 5465 16972 6257 1 FreeSans 2000 0 0 0 C[7]
port 25 nsew
flabel metal2 s 18816 5465 18860 6257 1 FreeSans 2000 0 0 0 C[6]
port 26 nsew
flabel metal2 s 20704 5465 20748 6257 1 FreeSans 2000 0 0 0 C[5]
port 27 nsew
flabel metal2 s 22592 5465 22636 6257 1 FreeSans 2000 0 0 0 C[4]
port 28 nsew
flabel metal2 s 24480 5465 24524 6257 1 FreeSans 2000 0 0 0 C[3]
port 29 nsew
flabel metal2 s 26368 5465 26412 6257 1 FreeSans 2000 0 0 0 C[2]
port 30 nsew
flabel metal2 s 28256 5465 28300 6257 1 FreeSans 2000 0 0 0 C[1]
port 31 nsew
flabel metal2 s 30144 5465 30188 6257 1 FreeSans 2000 0 0 0 C[0]
port 32 nsew
flabel metal4 s 1897 1 2235 6259 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 5681 0 6019 6258 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 9455 1 9793 6259 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 13233 1 13571 6259 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 17001 1 17339 6259 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 20773 1 21111 6259 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 24543 1 24881 6259 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 28331 0 28669 6258 1 FreeSans 2000 0 0 0 VSS
port 33 nsew
flabel metal4 s 3795 1 4133 6257 1 FreeSans 2000 0 0 0 VDD
port 34 nsew
flabel metal4 s 7571 1 7909 6257 1 FreeSans 2000 0 0 0 VDD
port 34 nsew
flabel metal4 s 11341 1 11679 6257 1 FreeSans 2000 0 0 0 VDD
port 34 nsew
flabel metal4 s 15109 1 15447 6257 1 FreeSans 2000 0 0 0 VDD
port 34 nsew
flabel metal4 s 18881 1 19219 6257 1 FreeSans 2000 0 0 0 VDD
port 34 nsew
flabel metal4 s 22649 1 22987 6257 1 FreeSans 2000 0 0 0 VDD
port 34 nsew
flabel metal4 s 26445 1 26783 6257 1 FreeSans 2000 0 0 0 VDD
port 34 nsew
flabel metal3 s 0 3036 536 3129 1 FreeSans 1000 0 0 0 RESET
port 35 nsew
flabel metal1 s 32375 782 32604 859 1 FreeSans 1000 0 0 0 OUT
port 36 nsew
<< end >>
