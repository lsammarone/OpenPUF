magic
tech sky130A
magscale 1 2
timestamp 1656307017
<< locali >>
rect 560520 582856 560827 582916
rect 560520 581430 560580 582856
rect 574316 582752 574638 582792
rect 565923 581536 566340 581596
rect 560362 581428 560908 581430
rect 560406 581370 560908 581428
rect 574316 581270 574356 582752
rect 579714 581372 580148 581432
rect 574344 581210 574746 581270
rect 574532 509262 574850 509302
rect 560374 509174 560758 509234
rect 560374 507764 560434 509174
rect 565840 507854 566212 507914
rect 574532 507800 574572 509262
rect 579986 507882 580388 507942
rect 560450 507686 560782 507746
rect 574586 507720 575030 507780
rect 560378 446468 560626 446528
rect 560378 445062 560438 446468
rect 574374 446282 574604 446322
rect 565696 445148 566062 445208
rect 560452 444982 560734 445042
rect 573711 444745 574124 444805
rect 574374 444800 574414 446282
rect 579724 444902 580092 444962
rect 574316 444740 574696 444800
rect 574344 403298 574614 403338
rect 560630 403208 560980 403268
rect 560630 402538 560690 403208
rect 560630 401782 560690 402420
rect 566060 401888 566434 401948
rect 574344 401818 574384 403298
rect 579736 401918 580130 401978
rect 560630 401722 561082 401782
rect 574406 401756 574774 401816
rect 574282 356856 574488 356896
rect 560358 356638 560718 356698
rect 560358 355218 560418 356638
rect 565735 355318 566208 355378
rect 574282 355382 574322 356856
rect 579640 355476 580084 355536
rect 574328 355314 574606 355374
rect 560426 355152 560732 355212
rect 560342 311618 560602 311678
rect 574280 311644 574638 311684
rect 560342 310204 560402 311618
rect 565689 310298 566178 310358
rect 560408 310132 560698 310192
rect 574280 310164 574320 311644
rect 579661 310264 580256 310324
rect 574334 310104 574676 310162
rect 574276 310102 574676 310104
<< viali >>
rect 566340 581520 566460 581634
rect 560334 581362 560406 581428
rect 580148 581372 580208 581432
rect 574284 581210 574344 581270
rect 566212 507840 566310 507940
rect 580388 507856 580498 507968
rect 560362 507684 560450 507764
rect 574502 507710 574586 507800
rect 566062 445132 566148 445220
rect 560354 444972 560452 445062
rect 574238 444730 574316 444806
rect 580092 444888 580182 444984
rect 560606 402420 560708 402538
rect 566434 401878 566514 401956
rect 580130 401904 580236 401996
rect 574330 401744 574406 401818
rect 566208 355300 566294 355406
rect 580084 355456 580174 355556
rect 574264 355304 574328 355382
rect 560348 355134 560426 355218
rect 566178 310286 566266 310370
rect 560334 310124 560408 310204
rect 580256 310246 580346 310344
rect 574274 310104 574334 310164
<< metal1 >>
rect 565961 583972 574678 584092
rect 565961 582986 566081 583972
rect 566334 583690 566510 583696
rect 566330 583578 566340 583690
rect 566492 583578 566510 583690
rect 566334 581640 566510 583578
rect 574558 583286 574678 583972
rect 580122 583568 580132 583676
rect 580222 583568 580232 583676
rect 566328 581634 566510 581640
rect 559778 581318 559788 581528
rect 560010 581442 560020 581528
rect 566328 581520 566340 581634
rect 566460 581520 566510 581634
rect 566328 581514 566510 581520
rect 573650 583166 574678 583286
rect 560010 581428 560420 581442
rect 573650 581438 573770 583166
rect 574558 582918 574678 583166
rect 580132 581438 580216 583568
rect 560010 581362 560334 581428
rect 560406 581362 560420 581428
rect 560010 581360 560420 581362
rect 560010 581318 560020 581360
rect 560322 581356 560418 581360
rect 559852 581226 559972 581318
rect 559852 581106 560887 581226
rect 565822 581106 572612 581226
rect 573618 581122 573628 581438
rect 573910 581278 573920 581438
rect 580132 581432 580220 581438
rect 580132 581372 580148 581432
rect 580208 581372 580220 581432
rect 580132 581366 580220 581372
rect 573910 581276 574352 581278
rect 573910 581270 574356 581276
rect 573910 581210 574284 581270
rect 574344 581210 574356 581270
rect 573910 581204 574356 581210
rect 573910 581186 574352 581204
rect 573910 581122 573920 581186
rect 572492 580962 572612 581106
rect 574882 580962 575002 581072
rect 572492 580842 575002 580962
rect 574066 509470 574886 509590
rect 574066 509424 574186 509470
rect 565728 509304 574186 509424
rect 566200 507830 566210 507952
rect 566316 507830 566326 507952
rect 573642 507912 573762 509304
rect 580382 507968 580504 507980
rect 566206 507828 566316 507830
rect 559794 507792 559914 507796
rect 559784 507678 559794 507792
rect 559918 507788 559928 507792
rect 559918 507770 560458 507788
rect 559918 507764 560462 507770
rect 559918 507684 560362 507764
rect 560450 507684 560462 507764
rect 559918 507678 560462 507684
rect 559794 507544 559914 507678
rect 573606 507620 573616 507912
rect 573914 507822 573924 507912
rect 580378 507856 580388 507968
rect 580498 507856 580508 507968
rect 580382 507844 580504 507856
rect 573914 507800 574594 507822
rect 573914 507710 574502 507800
rect 574586 507710 574594 507800
rect 573914 507698 574594 507710
rect 573914 507620 573924 507698
rect 559794 507424 560894 507544
rect 565574 507424 573414 507544
rect 573294 507384 573414 507424
rect 574796 507384 574916 507608
rect 573294 507264 574916 507384
rect 567252 446718 567262 446796
rect 565759 446598 567262 446718
rect 567252 446548 567262 446598
rect 567506 446548 567516 446796
rect 573564 446348 573574 446592
rect 573832 446532 573842 446592
rect 573832 446412 574956 446532
rect 573832 446348 573842 446412
rect 566056 445220 566154 445232
rect 566052 445132 566062 445220
rect 566148 445132 566158 445220
rect 566056 445120 566154 445132
rect 560342 445062 560464 445068
rect 560342 444972 560354 445062
rect 560452 444972 560464 445062
rect 580086 444984 580188 444996
rect 560342 444966 560464 444972
rect 580082 444888 580092 444984
rect 580182 444888 580192 444984
rect 580086 444876 580188 444888
rect 559844 444700 559854 444846
rect 559988 444838 559998 444846
rect 566810 444838 567030 444842
rect 559988 444718 560685 444838
rect 565398 444718 567030 444838
rect 574226 444806 574328 444812
rect 574226 444730 574238 444806
rect 574316 444730 574328 444806
rect 574226 444724 574328 444730
rect 559988 444700 559998 444718
rect 566810 444362 567030 444718
rect 574344 444532 575540 444652
rect 574344 444362 574464 444532
rect 566810 444142 574470 444362
rect 567264 403458 567274 403520
rect 565948 403338 567274 403458
rect 567264 403278 567274 403338
rect 567518 403278 567528 403520
rect 573582 403352 573592 403624
rect 573842 403548 573852 403624
rect 573842 403428 574742 403548
rect 573842 403352 573852 403428
rect 560600 402538 560714 402550
rect 560596 402420 560606 402538
rect 560708 402420 560718 402538
rect 560600 402408 560714 402420
rect 580118 401996 580248 402002
rect 566422 401956 566526 401962
rect 566422 401878 566434 401956
rect 566514 401878 566526 401956
rect 580118 401904 580130 401996
rect 580236 401904 580248 401996
rect 580118 401898 580248 401904
rect 566422 401872 566526 401878
rect 574318 401818 574418 401824
rect 574318 401744 574330 401818
rect 574406 401744 574418 401818
rect 574318 401738 574418 401744
rect 559760 401458 559844 401578
rect 559834 401456 559844 401458
rect 559968 401458 561112 401578
rect 565774 401458 566944 401578
rect 559968 401456 559978 401458
rect 566722 401409 566944 401458
rect 574514 401409 574666 401670
rect 566722 401187 574666 401409
rect 574514 401186 574666 401187
rect 567232 356888 567242 356952
rect 565616 356768 567242 356888
rect 567232 356694 567242 356768
rect 567508 356694 567518 356952
rect 573596 356914 573606 357166
rect 573850 357106 573860 357166
rect 573850 356986 574638 357106
rect 573850 356914 573860 356986
rect 580078 355556 580180 355568
rect 580074 355456 580084 355556
rect 580174 355456 580184 355556
rect 580078 355444 580180 355456
rect 566202 355406 566300 355418
rect 566198 355300 566208 355406
rect 566294 355300 566304 355406
rect 574258 355382 574334 355394
rect 574254 355304 574264 355382
rect 574328 355304 574338 355382
rect 566202 355288 566300 355300
rect 574258 355292 574334 355304
rect 560342 355218 560432 355230
rect 560338 355134 560348 355218
rect 560426 355134 560436 355218
rect 560342 355122 560432 355134
rect 559742 354888 559752 355008
rect 559872 354888 560764 355008
rect 565744 354888 566876 355008
rect 566756 354876 566876 354888
rect 574380 354876 574500 355218
rect 566756 354700 574500 354876
rect 567196 311868 567206 311944
rect 565566 311748 567206 311868
rect 567196 311670 567206 311748
rect 567462 311670 567472 311944
rect 573592 311692 573602 311954
rect 573864 311894 573874 311954
rect 573864 311774 574658 311894
rect 573864 311692 573874 311774
rect 566166 310370 566278 310376
rect 566166 310286 566178 310370
rect 566266 310286 566278 310370
rect 580250 310344 580352 310356
rect 566166 310280 566278 310286
rect 580246 310246 580256 310344
rect 580346 310246 580356 310344
rect 580250 310234 580352 310246
rect 560328 310204 560414 310216
rect 560324 310124 560334 310204
rect 560408 310124 560418 310204
rect 574262 310164 574346 310170
rect 560328 310112 560414 310124
rect 574262 310104 574274 310164
rect 574334 310104 574346 310164
rect 574262 310098 574346 310104
rect 559754 309868 559764 309988
rect 559884 309868 560724 309988
rect 565566 309868 566842 309988
rect 566722 309758 566842 309868
rect 574434 309758 574626 309974
rect 566722 309566 574626 309758
<< via1 >>
rect 566340 583578 566492 583690
rect 580132 583568 580222 583676
rect 559788 581318 560010 581528
rect 573628 581122 573910 581438
rect 566210 507940 566316 507952
rect 566210 507840 566212 507940
rect 566212 507840 566310 507940
rect 566310 507840 566316 507940
rect 566210 507830 566316 507840
rect 559794 507678 559918 507792
rect 573616 507620 573914 507912
rect 580388 507856 580498 507968
rect 567262 446548 567506 446796
rect 573574 446348 573832 446592
rect 566062 445132 566148 445220
rect 560354 444972 560452 445062
rect 580092 444888 580182 444984
rect 559854 444700 559988 444846
rect 574238 444730 574316 444806
rect 567274 403278 567518 403520
rect 573592 403352 573842 403624
rect 560606 402420 560708 402538
rect 566434 401878 566514 401956
rect 580130 401904 580236 401996
rect 574330 401744 574406 401818
rect 559844 401456 559968 401578
rect 567242 356694 567508 356952
rect 573606 356914 573850 357166
rect 580084 355456 580174 355556
rect 566208 355300 566294 355406
rect 574264 355304 574328 355382
rect 560348 355134 560426 355218
rect 559752 354888 559872 355008
rect 567206 311670 567462 311944
rect 573602 311692 573864 311954
rect 566178 310286 566266 310370
rect 580256 310246 580346 310344
rect 560334 310124 560408 310204
rect 574274 310104 574334 310164
rect 559764 309868 559884 309988
<< metal2 >>
rect 566340 583690 566492 583700
rect 566340 583568 566492 583578
rect 580132 583676 580222 583686
rect 580132 583558 580222 583568
rect 559788 581528 560010 581538
rect 559788 581308 560010 581318
rect 573628 581438 573910 581448
rect 573628 581112 573910 581122
rect 580388 507968 580498 507978
rect 566210 507956 566316 507962
rect 566204 507952 566316 507956
rect 566204 507946 566210 507952
rect 566204 507830 566210 507838
rect 566204 507828 566316 507830
rect 566210 507820 566316 507828
rect 573616 507912 573914 507922
rect 559794 507792 559918 507802
rect 559794 507668 559918 507678
rect 580388 507846 580498 507856
rect 573616 507610 573914 507620
rect 567262 446796 567506 446806
rect 567262 446538 567506 446548
rect 573574 446592 573832 446602
rect 573574 446338 573832 446348
rect 566062 445220 566148 445230
rect 566062 445122 566148 445132
rect 560354 445062 560452 445072
rect 560354 444962 560452 444972
rect 580092 444984 580182 444994
rect 580092 444878 580182 444888
rect 559854 444846 559988 444856
rect 574238 444806 574316 444816
rect 574238 444720 574316 444730
rect 559854 444690 559988 444700
rect 540316 435368 540422 435378
rect 540316 435296 540422 435306
rect 540304 419924 540448 419934
rect 540304 419834 540448 419844
rect 573592 403624 573842 403634
rect 567274 403520 567518 403530
rect 573592 403342 573842 403352
rect 567274 403268 567518 403278
rect 560606 402538 560708 402548
rect 560606 402410 560708 402420
rect 580130 401996 580236 402006
rect 566434 401956 566514 401966
rect 580130 401894 580236 401904
rect 566434 401868 566514 401878
rect 574330 401818 574406 401828
rect 574330 401734 574406 401744
rect 559844 401578 559968 401588
rect 559844 401446 559968 401456
rect 573606 357166 573850 357176
rect 567242 356952 567508 356962
rect 573606 356904 573850 356914
rect 567242 356684 567508 356694
rect 580084 355556 580174 355566
rect 580084 355446 580174 355456
rect 566208 355406 566294 355416
rect 566208 355290 566294 355300
rect 574264 355382 574328 355392
rect 574264 355294 574328 355304
rect 560348 355218 560426 355228
rect 560348 355124 560426 355134
rect 559752 355008 559872 355018
rect 559752 354878 559872 354888
rect 573602 311954 573864 311964
rect 567206 311944 567462 311954
rect 573602 311682 573864 311692
rect 567206 311660 567462 311670
rect 566178 310370 566266 310380
rect 566178 310276 566266 310286
rect 580256 310344 580346 310354
rect 580256 310236 580346 310246
rect 560334 310204 560408 310214
rect 560334 310114 560408 310124
rect 574274 310164 574334 310174
rect 574274 310094 574334 310104
rect 559764 309988 559884 309998
rect 559764 309858 559884 309868
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 566340 583578 566492 583690
rect 580132 583568 580222 583676
rect 559788 581318 560010 581528
rect 573628 581122 573910 581438
rect 566204 507838 566210 507946
rect 566210 507838 566316 507946
rect 559794 507678 559918 507792
rect 573616 507620 573914 507912
rect 580388 507856 580498 507968
rect 567262 446548 567506 446796
rect 573574 446348 573832 446592
rect 566062 445132 566148 445220
rect 560354 444972 560452 445062
rect 580092 444888 580182 444984
rect 559854 444700 559988 444846
rect 574238 444730 574316 444806
rect 540316 435306 540422 435368
rect 540304 419844 540448 419924
rect 567274 403278 567518 403520
rect 573592 403352 573842 403624
rect 560606 402420 560708 402538
rect 566434 401878 566514 401956
rect 580130 401904 580236 401996
rect 574330 401744 574406 401818
rect 559844 401456 559968 401578
rect 567242 356694 567508 356952
rect 573606 356914 573850 357166
rect 580084 355456 580174 355556
rect 566208 355300 566294 355406
rect 574264 355304 574328 355382
rect 560348 355134 560426 355218
rect 559752 354888 559872 355008
rect 567206 311670 567462 311944
rect 573602 311692 573864 311954
rect 566178 310286 566266 310370
rect 580256 310246 580346 310344
rect 560334 310124 560408 310204
rect 574274 310104 574334 310164
rect 559764 309868 559884 309988
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 703482 418394 704800
rect 413128 701890 418426 703482
rect 465394 702876 470394 704800
rect 510594 703613 515394 704800
rect 465042 702008 470794 702876
rect 510574 701285 515408 703613
rect 520594 703131 525394 704800
rect 510566 701189 515408 701285
rect 510566 700101 515400 701189
rect 520568 700588 525402 703131
rect 566594 702300 571594 704800
rect 510566 699600 515406 700101
rect 510550 698548 515406 699600
rect 520566 698548 525402 700588
rect 510550 687360 515248 698548
rect 520566 687360 525388 698548
rect 510550 687048 515408 687360
rect 520566 687048 525404 687360
rect 510554 686489 515408 687048
rect 510554 686163 515388 686489
rect 510554 685661 510737 686163
rect -800 680242 1700 685242
rect 510576 678739 510737 685661
rect 515201 678739 515388 686163
rect 510576 678487 515388 678739
rect 520570 686139 525404 687048
rect 520570 678715 520737 686139
rect 525201 678715 525404 686139
rect 520570 678548 525404 678715
rect 582300 677984 584800 682984
rect -800 643842 1660 648642
rect 567119 644605 581246 644615
rect 567119 644584 582932 644605
rect 567119 644323 584800 644584
rect 567119 640099 567336 644323
rect 573720 640099 584800 644323
rect 567119 639784 584800 640099
rect 567119 639769 582932 639784
rect -800 633842 1660 638642
rect 567322 634584 583190 634597
rect 567322 634265 584800 634584
rect 567310 634255 584800 634265
rect 567310 630031 567336 634255
rect 573720 630031 584800 634255
rect 567310 630021 584800 630031
rect 567322 629784 584800 630021
rect 567322 629761 583190 629784
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 507976 583288 507986 583852
rect 508658 583674 508668 583852
rect 566330 583690 566502 583695
rect 566330 583674 566340 583690
rect 508658 583578 566340 583674
rect 566492 583674 566502 583690
rect 580122 583676 580232 583681
rect 580122 583674 580132 583676
rect 566492 583578 580132 583674
rect 508658 583568 580132 583578
rect 580222 583674 580232 583676
rect 580222 583568 584800 583674
rect 508658 583562 584800 583568
rect 508658 583288 508668 583562
rect 559778 581528 560020 581533
rect 559778 581318 559788 581528
rect 560010 581318 560020 581528
rect 559778 581313 560020 581318
rect 573618 581438 573920 581443
rect 573618 581122 573628 581438
rect 573910 581122 573920 581438
rect 573618 581117 573920 581122
rect 457252 565074 457262 571686
rect 463874 571176 574176 571686
rect 463874 565074 566918 571176
rect 458534 564368 566918 565074
rect 574066 564368 574176 571176
rect -800 559442 1660 564242
rect 458534 564226 574176 564368
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 552438 543310 552448 543448
rect 533090 536792 552448 543310
rect 559104 543310 559114 543448
rect 559104 536792 559862 543310
rect 582340 540562 584800 545362
rect 533090 536654 559862 536792
rect 457490 515352 457500 515868
rect -800 511530 480 511642
rect -800 510348 480 510460
rect 457142 509644 457500 515352
rect 463724 515352 463734 515868
rect 463724 509644 493426 515352
rect -800 509166 480 509278
rect -800 507984 480 508096
rect 457142 507742 493426 509644
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 457142 501632 457846 507742
rect 457836 501518 457846 501632
rect 464070 501632 493426 507742
rect 524200 513300 543128 513312
rect 524200 506708 554094 513300
rect 580380 507973 580582 507980
rect 580378 507968 580582 507973
rect 566200 507951 566210 507952
rect 566194 507946 566210 507951
rect 566194 507838 566204 507946
rect 566316 507944 566326 507952
rect 566194 507833 566210 507838
rect 566200 507830 566210 507833
rect 566316 507830 566412 507944
rect 559784 507792 559928 507797
rect 559784 507678 559794 507792
rect 559918 507678 559928 507792
rect 559784 507673 559928 507678
rect 566208 506708 566412 507830
rect 573606 507912 573924 507917
rect 573606 507620 573616 507912
rect 573914 507620 573924 507912
rect 580378 507856 580388 507968
rect 580498 507856 580582 507968
rect 580378 507851 580582 507856
rect 573606 507615 573924 507620
rect 580380 506708 580582 507851
rect 464070 501518 464080 501632
rect 524200 497912 581748 506708
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 544502 494257 581748 497912
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 544502 494252 583876 494257
rect 544502 494140 584800 494252
rect 544502 494133 583876 494140
rect 544502 492988 581748 494133
rect 533090 479346 553036 486002
rect 559692 479346 559702 486002
rect 457120 472368 574088 472534
rect 457120 472012 566954 472368
rect 457120 471992 535652 472012
rect -800 468308 480 468420
rect -800 467126 480 467238
rect 457120 466286 457230 471992
rect 463886 471814 535652 471992
rect 463886 471788 488088 471814
rect 463886 471134 487194 471788
rect 487810 471160 488088 471788
rect 488704 471358 535652 471814
rect 536268 471358 536478 472012
rect 537094 471358 566954 472012
rect 488704 471160 566954 471358
rect 487810 471134 566954 471160
rect 463886 470812 566954 471134
rect 463886 470614 535652 470812
rect 463886 470588 488088 470614
rect 463886 469934 487194 470588
rect 487810 469960 488088 470588
rect 488704 470158 535652 470614
rect 536268 470158 536478 470812
rect 537094 470158 566954 470812
rect 488704 469960 566954 470158
rect 487810 469934 566954 469960
rect 463886 469612 566954 469934
rect 463886 469414 535652 469612
rect 463886 469388 488088 469414
rect 463886 468734 487194 469388
rect 487810 468760 488088 469388
rect 488704 468958 535652 469414
rect 536268 468958 536478 469612
rect 537094 468958 566954 469612
rect 488704 468760 566954 468958
rect 487810 468734 566954 468760
rect 463886 468412 566954 468734
rect 463886 468214 535652 468412
rect 463886 468188 488088 468214
rect 463886 467534 487194 468188
rect 487810 467560 488088 468188
rect 488704 467758 535652 468214
rect 536268 467758 536478 468412
rect 537094 467758 566954 468412
rect 488704 467560 566954 467758
rect 487810 467534 566954 467560
rect 463886 467212 566954 467534
rect 463886 467014 535652 467212
rect 463886 466988 488088 467014
rect 463886 466334 487194 466988
rect 487810 466360 488088 466988
rect 488704 466558 535652 467014
rect 536268 466558 536478 467212
rect 537094 466558 566954 467212
rect 488704 466360 566954 466558
rect 487810 466334 566954 466360
rect 463886 466286 566954 466334
rect -800 465944 480 466056
rect 457120 465896 566954 466286
rect 574254 465896 574264 472368
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 542181 449830 582982 450926
rect 583520 450900 584800 451012
rect 542181 449718 584800 449830
rect 542181 447208 582982 449718
rect 542181 435432 545899 447208
rect 566266 445252 566394 447208
rect 567252 446796 567516 446801
rect 567252 446548 567262 446796
rect 567506 446548 567516 446796
rect 567252 446543 567516 446548
rect 573564 446592 573842 446597
rect 573564 446348 573574 446592
rect 573832 446348 573842 446592
rect 573564 446343 573842 446348
rect 566048 445220 566394 445252
rect 566048 445132 566062 445220
rect 566148 445132 566394 445220
rect 566048 445114 566394 445132
rect 559850 445082 560466 445084
rect 559838 444942 559848 445082
rect 559996 445062 560466 445082
rect 559996 444972 560354 445062
rect 560452 444972 560466 445062
rect 580262 445010 580402 447208
rect 559996 444948 560466 444972
rect 580080 444984 580402 445010
rect 559996 444942 560006 444948
rect 559824 444700 559834 444854
rect 560008 444700 560018 444854
rect 559844 444695 559998 444700
rect 573582 444642 573592 444908
rect 573890 444834 573900 444908
rect 580080 444888 580092 444984
rect 580182 444888 580402 444984
rect 580080 444870 580402 444888
rect 580080 444860 580322 444870
rect 573890 444806 574330 444834
rect 573890 444730 574238 444806
rect 574316 444730 574330 444806
rect 573890 444712 574330 444730
rect 573890 444642 573900 444712
rect 540288 435368 545899 435432
rect 540288 435306 540316 435368
rect 540422 435306 545899 435368
rect 540288 435222 545899 435306
rect 542181 434678 545899 435222
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect 541532 419980 544951 420358
rect 540284 419924 544951 419980
rect 540284 419844 540304 419924
rect 540448 419844 544951 419924
rect 540284 419812 544951 419844
rect -800 419176 480 419288
rect 541532 419247 544951 419812
rect 541537 407656 544951 419247
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 541537 405409 582845 407656
rect 583520 406478 584800 406590
rect 541537 405408 583886 405409
rect 541537 405297 584800 405408
rect 541537 404242 582845 405297
rect 583520 405296 584800 405297
rect 559743 402374 559804 402584
rect 559794 402372 559804 402374
rect 559994 402538 560730 402584
rect 559994 402420 560606 402538
rect 560708 402420 560730 402538
rect 559994 402374 560730 402420
rect 559994 402372 560004 402374
rect 566412 401956 566548 404242
rect 573582 403624 573852 403629
rect 567264 403520 567528 403525
rect 567264 403278 567274 403520
rect 567518 403278 567528 403520
rect 573582 403352 573592 403624
rect 573842 403352 573852 403624
rect 573582 403347 573852 403352
rect 567264 403273 567528 403278
rect 580264 402040 580440 404242
rect 566412 401878 566434 401956
rect 566514 401878 566548 401956
rect 580090 401996 580440 402040
rect 566412 401864 566548 401878
rect 573638 401658 573648 401912
rect 573884 401852 573894 401912
rect 580090 401904 580130 401996
rect 580236 401904 580440 401996
rect 580090 401864 580440 401904
rect 573884 401818 574422 401852
rect 573884 401744 574330 401818
rect 574406 401744 574422 401818
rect 573884 401730 574422 401744
rect 573884 401658 573894 401730
rect 559834 401578 559978 401583
rect 559834 401456 559844 401578
rect 559968 401456 559978 401578
rect 559834 401451 559978 401456
rect 484398 394112 573636 394226
rect 484398 394104 488026 394112
rect 484398 393598 487244 394104
rect 487754 393606 488026 394104
rect 488536 394060 573636 394112
rect 488536 394020 536458 394060
rect 488536 393688 535658 394020
rect 536176 393728 536458 394020
rect 536976 394012 573636 394060
rect 536976 393998 571960 394012
rect 536976 393986 570844 393998
rect 536976 393728 567458 393986
rect 536176 393688 567458 393728
rect 488536 393606 567458 393688
rect 487754 393598 567458 393606
rect 484398 393560 567458 393598
rect 484398 393520 536458 393560
rect 484398 393512 535658 393520
rect 484398 393504 488026 393512
rect 484398 392998 487244 393504
rect 487754 393006 488026 393504
rect 488536 393188 535658 393512
rect 536176 393228 536458 393520
rect 536976 393494 567458 393560
rect 568134 393494 568626 393986
rect 569302 393494 569754 393986
rect 570430 393506 570844 393986
rect 571520 393520 571960 393998
rect 572636 393520 573636 394012
rect 571520 393506 573636 393520
rect 570430 393494 573636 393506
rect 536976 393284 573636 393494
rect 536976 393272 571960 393284
rect 536976 393258 570856 393272
rect 536976 393246 569742 393258
rect 536976 393228 568612 393246
rect 536176 393220 568612 393228
rect 536176 393188 567484 393220
rect 488536 393060 567484 393188
rect 488536 393020 536458 393060
rect 488536 393006 535658 393020
rect 487754 392998 535658 393006
rect 484398 392912 535658 392998
rect 484398 392904 488026 392912
rect 484398 392398 487244 392904
rect 487754 392406 488026 392904
rect 488536 392688 535658 392912
rect 536176 392728 536458 393020
rect 536976 392728 567484 393060
rect 568160 392754 568612 393220
rect 569288 392766 569742 393246
rect 570418 392780 570856 393258
rect 571532 392792 571960 393272
rect 572636 392792 573636 393284
rect 571532 392780 573636 392792
rect 570418 392766 573636 392780
rect 569288 392754 573636 392766
rect 568160 392728 573636 392754
rect 536176 392688 573636 392728
rect 488536 392560 573636 392688
rect 488536 392520 536458 392560
rect 488536 392406 535658 392520
rect 487754 392398 535658 392406
rect 484398 392312 535658 392398
rect 484398 392304 488026 392312
rect 484398 391798 487244 392304
rect 487754 391806 488026 392304
rect 488536 392188 535658 392312
rect 536176 392228 536458 392520
rect 536976 392520 573636 392560
rect 536976 392494 570870 392520
rect 536976 392468 569768 392494
rect 536976 392454 568612 392468
rect 536976 392228 567498 392454
rect 536176 392188 567498 392228
rect 488536 392060 567498 392188
rect 488536 392020 536458 392060
rect 488536 391806 535658 392020
rect 487754 391798 535658 391806
rect 484398 391714 535658 391798
rect 535648 391688 535658 391714
rect 536176 391728 536458 392020
rect 536976 391962 567498 392060
rect 568174 391976 568612 392454
rect 569288 392002 569768 392468
rect 570444 392028 570870 392494
rect 571546 392506 573636 392520
rect 571546 392028 571934 392506
rect 570444 392014 571934 392028
rect 572610 392014 573636 392506
rect 570444 392002 573636 392014
rect 569288 391976 573636 392002
rect 568174 391962 573636 391976
rect 536976 391728 573636 391962
rect 536176 391714 573636 391728
rect 536176 391688 536186 391714
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 481374 371880 577042 372170
rect 481374 371614 491672 371880
rect 492902 371822 577042 371880
rect 492902 371614 537048 371822
rect 481374 371556 537048 371614
rect 538278 371804 577042 371822
rect 538278 371778 569548 371804
rect 538278 371556 567382 371778
rect 481374 371388 567382 371556
rect 481374 371122 491672 371388
rect 492902 371360 567382 371388
rect 492902 371122 537066 371360
rect 481374 371094 537066 371122
rect 538296 371094 567382 371360
rect 481374 370886 567382 371094
rect 481374 370620 491682 370886
rect 492912 370810 567382 370886
rect 492912 370620 537076 370810
rect 481374 370544 537076 370620
rect 538306 370544 567382 370810
rect 481374 370412 567382 370544
rect 481374 370146 491690 370412
rect 492920 370318 567382 370412
rect 492920 370146 537076 370318
rect 481374 370052 537076 370146
rect 538306 370316 567382 370318
rect 569210 370342 569548 371778
rect 571376 370342 571674 371804
rect 573502 370342 577042 371804
rect 569210 370316 577042 370342
rect 538306 370052 577042 370316
rect 481374 370042 577042 370052
rect 481374 370028 571688 370042
rect 481374 369976 569548 370028
rect 481374 369882 567396 369976
rect 481374 369616 491672 369882
rect 492902 369788 567396 369882
rect 492902 369616 537086 369788
rect 481374 369522 537086 369616
rect 538316 369522 567396 369788
rect 481374 369362 567396 369522
rect 481374 369096 491672 369362
rect 492902 369286 567396 369362
rect 492902 369096 537066 369286
rect 481374 369020 537066 369096
rect 538296 369246 567396 369286
rect 569170 369298 569548 369976
rect 571322 369312 571688 370028
rect 573462 369312 577042 370042
rect 571322 369298 577042 369312
rect 569170 369246 577042 369298
rect 538296 369020 577042 369246
rect 481374 368832 577042 369020
rect 481374 368566 491682 368832
rect 492912 368804 577042 368832
rect 492912 368566 537076 368804
rect 481374 368538 537076 368566
rect 538306 368778 577042 368804
rect 538306 368752 571714 368778
rect 538306 368700 569536 368752
rect 538306 368538 567396 368700
rect 481374 368340 567396 368538
rect 481374 368074 491690 368340
rect 492920 368236 567396 368340
rect 492920 368074 537094 368236
rect 481374 367970 537094 368074
rect 538324 367970 567396 368236
rect 481374 367914 567396 367970
rect 481374 367648 491682 367914
rect 492912 367810 567396 367914
rect 492912 367648 537086 367810
rect 481374 367544 537086 367648
rect 538316 367544 567396 367810
rect 481374 367450 567396 367544
rect 481374 367184 491690 367450
rect 492920 367394 567396 367450
rect 492920 367184 537086 367394
rect 481374 367128 537086 367184
rect 538316 367290 567396 367394
rect 569118 367342 569536 368700
rect 571258 367368 571714 368752
rect 573436 367368 577042 368778
rect 571258 367342 577042 367368
rect 569118 367290 577042 367342
rect 538316 367128 577042 367290
rect 481374 367048 577042 367128
rect 583520 364784 584800 364896
rect 542526 364026 550666 364416
rect 541204 363514 550666 364026
rect 583520 363602 584800 363714
rect 542526 361160 550666 363514
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 547410 360812 550666 361160
rect 547410 358993 582986 360812
rect 583520 360056 584800 360168
rect 547410 358986 583854 358993
rect 547410 358875 584800 358986
rect 547410 357556 582986 358875
rect 583520 358874 584800 358875
rect 566176 355406 566328 357556
rect 573596 357166 573860 357171
rect 567232 356952 567518 356957
rect 567232 356694 567242 356952
rect 567508 356694 567518 356952
rect 573596 356914 573606 357166
rect 573850 356914 573860 357166
rect 573596 356909 573860 356914
rect 567232 356689 567518 356694
rect 580062 355556 580192 357556
rect 566176 355300 566208 355406
rect 566294 355300 566328 355406
rect 566176 355282 566328 355300
rect 559942 355244 560446 355246
rect 559890 355116 559900 355244
rect 560014 355218 560446 355244
rect 573650 355236 573660 355486
rect 573898 355412 573908 355486
rect 580062 355456 580084 355556
rect 580174 355456 580192 355556
rect 580062 355434 580192 355456
rect 573898 355382 574346 355412
rect 573898 355304 574264 355382
rect 574328 355304 574346 355382
rect 573898 355290 574346 355304
rect 573898 355236 573908 355290
rect 560014 355134 560348 355218
rect 560426 355134 560446 355218
rect 560014 355120 560446 355134
rect 560014 355116 560024 355120
rect 559742 355008 559882 355013
rect 559742 354888 559752 355008
rect 559872 354888 559882 355008
rect 559742 354883 559882 354888
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 544592 313779 583148 314974
rect 583520 314834 584800 314946
rect 544592 313764 583752 313779
rect 544592 313652 584800 313764
rect 544592 313602 583887 313652
rect 544592 312682 583148 313602
rect 544592 309524 546884 312682
rect 566201 310382 566368 312682
rect 573592 311954 573874 311959
rect 567196 311944 567472 311949
rect 567196 311670 567206 311944
rect 567462 311670 567472 311944
rect 573592 311692 573602 311954
rect 573864 311692 573874 311954
rect 573592 311687 573874 311692
rect 567196 311665 567472 311670
rect 566146 310370 566368 310382
rect 566146 310286 566178 310370
rect 566266 310286 566368 310370
rect 566146 310272 566368 310286
rect 580240 310344 580384 312682
rect 559962 310208 560424 310220
rect 559952 310118 559962 310208
rect 560026 310204 560424 310208
rect 560026 310124 560334 310204
rect 560408 310124 560424 310204
rect 560026 310118 560424 310124
rect 559962 310108 560424 310118
rect 573640 310034 573650 310278
rect 573894 310190 573904 310278
rect 580240 310246 580256 310344
rect 580346 310246 580384 310344
rect 580240 310228 580384 310246
rect 573894 310164 574348 310190
rect 573894 310104 574274 310164
rect 574334 310104 574348 310164
rect 573894 310084 574348 310104
rect 573894 310034 573904 310084
rect 559754 309988 559894 309993
rect 559754 309868 559764 309988
rect 559884 309868 559894 309988
rect 559754 309863 559894 309868
rect 541204 309040 546884 309524
rect 544592 308556 546884 309040
rect 482880 305824 578548 306030
rect 482880 305792 567402 305824
rect 482880 305288 491614 305792
rect 492938 305756 567402 305792
rect 492938 305288 536988 305756
rect 482880 305252 536988 305288
rect 538312 305252 567402 305756
rect 482880 304982 567402 305252
rect 482880 304478 491634 304982
rect 492958 304934 567402 304982
rect 492958 304478 536988 304934
rect 482880 304430 536988 304478
rect 538312 304430 567402 304934
rect 482880 304414 567402 304430
rect 569124 304414 569488 305824
rect 571210 304414 571510 305824
rect 573232 304414 578548 305824
rect 482880 304200 578548 304414
rect 482880 303696 491634 304200
rect 492958 304184 578548 304200
rect 492958 304132 571484 304184
rect 492958 303696 537026 304132
rect 482880 303628 537026 303696
rect 538350 304092 569488 304132
rect 538350 303628 567414 304092
rect 482880 303408 567414 303628
rect 482880 302904 491652 303408
rect 492976 303350 567414 303408
rect 492976 302904 537026 303350
rect 482880 302846 537026 302904
rect 538350 302846 567414 303350
rect 482880 302682 567414 302846
rect 569136 302722 569488 304092
rect 571210 302774 571484 304132
rect 573206 302774 578548 304184
rect 571210 302722 578548 302774
rect 569136 302682 578548 302722
rect 482880 302646 578548 302682
rect 482880 302142 491652 302646
rect 492976 302566 578548 302646
rect 492976 302142 537026 302566
rect 482880 302062 537026 302142
rect 538350 302452 578548 302566
rect 538350 302412 571536 302452
rect 538350 302400 569462 302412
rect 538350 302062 567440 302400
rect 482880 301846 567440 302062
rect 482880 301342 491662 301846
rect 492986 301708 567440 301846
rect 492986 301342 537026 301708
rect 482880 301204 537026 301342
rect 538350 301204 567440 301708
rect 482880 300990 567440 301204
rect 569162 301002 569462 302400
rect 571184 301042 571536 302412
rect 573258 301042 578548 302452
rect 571184 301002 578548 301042
rect 569162 300990 578548 301002
rect 482880 300908 578548 300990
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 510737 678739 515201 686163
rect 520737 678715 525201 686139
rect 567336 640099 573720 644323
rect 567336 630031 573720 634255
rect 507986 583288 508658 583852
rect 559788 581318 560010 581528
rect 573628 581122 573910 581438
rect 457262 565074 463874 571686
rect 566918 564368 574066 571176
rect 552448 536792 559104 543448
rect 457500 509644 463724 515868
rect 457846 501518 464070 507742
rect 566210 507946 566316 507952
rect 566210 507838 566316 507946
rect 566210 507830 566316 507838
rect 559794 507678 559918 507792
rect 573616 507620 573914 507912
rect 553036 479346 559692 486002
rect 457230 466286 463886 471992
rect 487194 471134 487810 471788
rect 488088 471160 488704 471814
rect 535652 471358 536268 472012
rect 536478 471358 537094 472012
rect 487194 469934 487810 470588
rect 488088 469960 488704 470614
rect 535652 470158 536268 470812
rect 536478 470158 537094 470812
rect 487194 468734 487810 469388
rect 488088 468760 488704 469414
rect 535652 468958 536268 469612
rect 536478 468958 537094 469612
rect 487194 467534 487810 468188
rect 488088 467560 488704 468214
rect 535652 467758 536268 468412
rect 536478 467758 537094 468412
rect 487194 466334 487810 466988
rect 488088 466360 488704 467014
rect 535652 466558 536268 467212
rect 536478 466558 537094 467212
rect 566954 465896 574254 472368
rect 567262 446548 567506 446796
rect 573574 446348 573832 446592
rect 559848 444942 559996 445082
rect 559834 444846 560008 444854
rect 559834 444700 559854 444846
rect 559854 444700 559988 444846
rect 559988 444700 560008 444846
rect 573592 444642 573890 444908
rect 559804 402372 559994 402584
rect 567274 403278 567518 403520
rect 573592 403352 573842 403624
rect 573648 401658 573884 401912
rect 559844 401456 559968 401578
rect 487244 393598 487754 394104
rect 488026 393606 488536 394112
rect 535658 393688 536176 394020
rect 536458 393728 536976 394060
rect 487244 392998 487754 393504
rect 488026 393006 488536 393512
rect 535658 393188 536176 393520
rect 536458 393228 536976 393560
rect 567458 393494 568134 393986
rect 568626 393494 569302 393986
rect 569754 393494 570430 393986
rect 570844 393506 571520 393998
rect 571960 393520 572636 394012
rect 487244 392398 487754 392904
rect 488026 392406 488536 392912
rect 535658 392688 536176 393020
rect 536458 392728 536976 393060
rect 567484 392728 568160 393220
rect 568612 392754 569288 393246
rect 569742 392766 570418 393258
rect 570856 392780 571532 393272
rect 571960 392792 572636 393284
rect 487244 391798 487754 392304
rect 488026 391806 488536 392312
rect 535658 392188 536176 392520
rect 536458 392228 536976 392560
rect 535658 391688 536176 392020
rect 536458 391728 536976 392060
rect 567498 391962 568174 392454
rect 568612 391976 569288 392468
rect 569768 392002 570444 392494
rect 570870 392028 571546 392520
rect 571934 392014 572610 392506
rect 491672 371614 492902 371880
rect 537048 371556 538278 371822
rect 491672 371122 492902 371388
rect 537066 371094 538296 371360
rect 491682 370620 492912 370886
rect 537076 370544 538306 370810
rect 491690 370146 492920 370412
rect 537076 370052 538306 370318
rect 567382 370316 569210 371778
rect 569548 370342 571376 371804
rect 571674 370342 573502 371804
rect 491672 369616 492902 369882
rect 537086 369522 538316 369788
rect 491672 369096 492902 369362
rect 537066 369020 538296 369286
rect 567396 369246 569170 369976
rect 569548 369298 571322 370028
rect 571688 369312 573462 370042
rect 491682 368566 492912 368832
rect 537076 368538 538306 368804
rect 491690 368074 492920 368340
rect 537094 367970 538324 368236
rect 491682 367648 492912 367914
rect 537086 367544 538316 367810
rect 491690 367184 492920 367450
rect 537086 367128 538316 367394
rect 567396 367290 569118 368700
rect 569536 367342 571258 368752
rect 571714 367368 573436 368778
rect 567242 356694 567508 356952
rect 573606 356914 573850 357166
rect 559900 355116 560014 355244
rect 573660 355236 573898 355486
rect 559752 354888 559872 355008
rect 567206 311670 567462 311944
rect 573602 311692 573864 311954
rect 559962 310118 560026 310208
rect 573650 310034 573894 310278
rect 559764 309868 559884 309988
rect 491614 305288 492938 305792
rect 536988 305252 538312 305756
rect 491634 304478 492958 304982
rect 536988 304430 538312 304934
rect 567402 304414 569124 305824
rect 569488 304414 571210 305824
rect 571510 304414 573232 305824
rect 491634 303696 492958 304200
rect 537026 303628 538350 304132
rect 491652 302904 492976 303408
rect 537026 302846 538350 303350
rect 567414 302682 569136 304092
rect 569488 302722 571210 304132
rect 571484 302774 573206 304184
rect 491652 302142 492976 302646
rect 537026 302062 538350 302566
rect 491662 301342 492986 301846
rect 537026 301204 538350 301708
rect 567440 300990 569162 302400
rect 569462 301002 571184 302412
rect 571536 301042 573258 302452
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 395244 686163 560048 686611
rect 395244 678739 510737 686163
rect 515201 686139 560048 686163
rect 515201 678739 520737 686139
rect 395244 678715 520737 678739
rect 525201 678715 560048 686139
rect 395244 678563 560048 678715
rect 507985 583852 508659 583853
rect 507985 583288 507986 583852
rect 508658 583288 508659 583852
rect 507985 583287 508659 583288
rect 457261 571686 463875 571687
rect 457261 565074 457262 571686
rect 463874 565074 463875 571686
rect 457261 565073 463875 565074
rect 457262 515868 463874 565073
rect 508046 547268 508622 583287
rect 551988 581528 560036 678563
rect 567319 644323 573737 644334
rect 567319 640099 567336 644323
rect 573720 640099 573737 644323
rect 567319 640088 573737 640099
rect 567319 634255 573737 634266
rect 567319 630031 567336 634255
rect 573720 630031 573737 634255
rect 567319 630020 573737 630031
rect 551988 581318 559788 581528
rect 560010 581318 560036 581528
rect 457262 509644 457500 515868
rect 463724 509644 463874 515868
rect 457262 507743 463874 509644
rect 551988 543448 560036 581318
rect 573627 581438 573911 581439
rect 573627 581122 573628 581438
rect 573910 581122 573911 581438
rect 573627 581121 573911 581122
rect 566917 571176 574067 571177
rect 566917 564368 566918 571176
rect 574066 564368 574067 571176
rect 566917 564367 574067 564368
rect 551988 536792 552448 543448
rect 559104 536792 560036 543448
rect 551988 507792 560036 536792
rect 566209 507952 566317 507953
rect 566209 507830 566210 507952
rect 566316 507830 566317 507952
rect 566209 507829 566317 507830
rect 573615 507912 573915 507913
rect 457262 507742 464071 507743
rect 457262 501518 457846 507742
rect 464070 501518 464071 507742
rect 457262 501517 464071 501518
rect 551988 507678 559794 507792
rect 559918 507678 560036 507792
rect 457262 471993 463874 501517
rect 551988 486002 560036 507678
rect 573615 507620 573616 507912
rect 573914 507620 573915 507912
rect 573615 507619 573915 507620
rect 551988 479346 553036 486002
rect 559692 479346 560036 486002
rect 535651 472012 536269 472013
rect 457229 471992 463887 471993
rect 457229 466286 457230 471992
rect 463886 466286 463887 471992
rect 488087 471814 488705 471815
rect 487193 471788 487811 471789
rect 487193 471134 487194 471788
rect 487810 471134 487811 471788
rect 488087 471160 488088 471814
rect 488704 471160 488705 471814
rect 535651 471358 535652 472012
rect 536268 471358 536269 472012
rect 535651 471357 536269 471358
rect 536477 472012 537095 472013
rect 536477 471358 536478 472012
rect 537094 471358 537095 472012
rect 536477 471357 537095 471358
rect 488087 471159 488705 471160
rect 487193 471133 487811 471134
rect 535651 470812 536269 470813
rect 488087 470614 488705 470615
rect 487193 470588 487811 470589
rect 487193 469934 487194 470588
rect 487810 469934 487811 470588
rect 488087 469960 488088 470614
rect 488704 469960 488705 470614
rect 535651 470158 535652 470812
rect 536268 470158 536269 470812
rect 535651 470157 536269 470158
rect 536477 470812 537095 470813
rect 536477 470158 536478 470812
rect 537094 470158 537095 470812
rect 536477 470157 537095 470158
rect 488087 469959 488705 469960
rect 487193 469933 487811 469934
rect 535651 469612 536269 469613
rect 488087 469414 488705 469415
rect 487193 469388 487811 469389
rect 487193 468734 487194 469388
rect 487810 468734 487811 469388
rect 488087 468760 488088 469414
rect 488704 468760 488705 469414
rect 535651 468958 535652 469612
rect 536268 468958 536269 469612
rect 535651 468957 536269 468958
rect 536477 469612 537095 469613
rect 536477 468958 536478 469612
rect 537094 468958 537095 469612
rect 536477 468957 537095 468958
rect 488087 468759 488705 468760
rect 487193 468733 487811 468734
rect 535651 468412 536269 468413
rect 488087 468214 488705 468215
rect 487193 468188 487811 468189
rect 487193 467534 487194 468188
rect 487810 467534 487811 468188
rect 488087 467560 488088 468214
rect 488704 467560 488705 468214
rect 535651 467758 535652 468412
rect 536268 467758 536269 468412
rect 535651 467757 536269 467758
rect 536477 468412 537095 468413
rect 536477 467758 536478 468412
rect 537094 467758 537095 468412
rect 536477 467757 537095 467758
rect 488087 467559 488705 467560
rect 487193 467533 487811 467534
rect 535651 467212 536269 467213
rect 488087 467014 488705 467015
rect 487193 466988 487811 466989
rect 487193 466334 487194 466988
rect 487810 466334 487811 466988
rect 488087 466360 488088 467014
rect 488704 466360 488705 467014
rect 535651 466558 535652 467212
rect 536268 466558 536269 467212
rect 535651 466557 536269 466558
rect 536477 467212 537095 467213
rect 536477 466558 536478 467212
rect 537094 466558 537095 467212
rect 536477 466557 537095 466558
rect 488087 466359 488705 466360
rect 487193 466333 487811 466334
rect 457229 466285 463887 466286
rect 551988 454814 560036 479346
rect 566953 472368 574255 472369
rect 566953 465896 566954 472368
rect 574254 465896 574255 472368
rect 566953 465895 574255 465896
rect 533228 453182 560036 454814
rect 551988 445694 560036 453182
rect 567261 446796 567507 446797
rect 567261 446548 567262 446796
rect 567506 446548 567507 446796
rect 567261 446547 567507 446548
rect 573573 446592 573833 446593
rect 573573 446348 573574 446592
rect 573832 446348 573833 446592
rect 573573 446347 573833 446348
rect 551964 445082 560036 445694
rect 551964 444942 559848 445082
rect 559996 444942 560036 445082
rect 551964 444854 560036 444942
rect 551964 444700 559834 444854
rect 560008 444700 560036 444854
rect 551964 444696 560036 444700
rect 551988 402584 560036 444696
rect 573591 444908 573891 444909
rect 573591 444642 573592 444908
rect 573890 444642 573891 444908
rect 573591 444641 573891 444642
rect 573591 403624 573843 403625
rect 567273 403520 567519 403521
rect 567273 403278 567274 403520
rect 567518 403278 567519 403520
rect 573591 403352 573592 403624
rect 573842 403352 573843 403624
rect 573591 403351 573843 403352
rect 567273 403277 567519 403278
rect 551988 402372 559804 402584
rect 559994 402372 560036 402584
rect 551988 401578 560036 402372
rect 573647 401912 573885 401913
rect 573647 401658 573648 401912
rect 573884 401658 573885 401912
rect 573647 401657 573885 401658
rect 551988 401456 559844 401578
rect 559968 401456 560036 401578
rect 551988 399810 560036 401456
rect 528746 398178 560036 399810
rect 488025 394112 488537 394113
rect 487243 394104 487755 394105
rect 487243 393598 487244 394104
rect 487754 393598 487755 394104
rect 488025 393606 488026 394112
rect 488536 393606 488537 394112
rect 536457 394060 536977 394061
rect 535657 394020 536177 394021
rect 535657 393688 535658 394020
rect 536176 393688 536177 394020
rect 536457 393728 536458 394060
rect 536976 393728 536977 394060
rect 536457 393727 536977 393728
rect 535657 393687 536177 393688
rect 488025 393605 488537 393606
rect 487243 393597 487755 393598
rect 536457 393560 536977 393561
rect 535657 393520 536177 393521
rect 488025 393512 488537 393513
rect 487243 393504 487755 393505
rect 487243 392998 487244 393504
rect 487754 392998 487755 393504
rect 488025 393006 488026 393512
rect 488536 393006 488537 393512
rect 535657 393188 535658 393520
rect 536176 393188 536177 393520
rect 536457 393228 536458 393560
rect 536976 393228 536977 393560
rect 536457 393227 536977 393228
rect 535657 393187 536177 393188
rect 536457 393060 536977 393061
rect 488025 393005 488537 393006
rect 535657 393020 536177 393021
rect 487243 392997 487755 392998
rect 488025 392912 488537 392913
rect 487243 392904 487755 392905
rect 487243 392398 487244 392904
rect 487754 392398 487755 392904
rect 488025 392406 488026 392912
rect 488536 392406 488537 392912
rect 535657 392688 535658 393020
rect 536176 392688 536177 393020
rect 536457 392728 536458 393060
rect 536976 392728 536977 393060
rect 536457 392727 536977 392728
rect 535657 392687 536177 392688
rect 536457 392560 536977 392561
rect 488025 392405 488537 392406
rect 535657 392520 536177 392521
rect 487243 392397 487755 392398
rect 488025 392312 488537 392313
rect 487243 392304 487755 392305
rect 487243 391798 487244 392304
rect 487754 391798 487755 392304
rect 488025 391806 488026 392312
rect 488536 391806 488537 392312
rect 535657 392188 535658 392520
rect 536176 392188 536177 392520
rect 536457 392228 536458 392560
rect 536976 392228 536977 392560
rect 536457 392227 536977 392228
rect 535657 392187 536177 392188
rect 536457 392060 536977 392061
rect 488025 391805 488537 391806
rect 535657 392020 536177 392021
rect 487243 391797 487755 391798
rect 535657 391688 535658 392020
rect 536176 391688 536177 392020
rect 536457 391728 536458 392060
rect 536976 391728 536977 392060
rect 536457 391727 536977 391728
rect 535657 391687 536177 391688
rect 551988 377437 560036 398178
rect 571959 394012 572637 394013
rect 570843 393998 571521 393999
rect 567457 393986 568135 393987
rect 567457 393494 567458 393986
rect 568134 393494 568135 393986
rect 567457 393493 568135 393494
rect 568625 393986 569303 393987
rect 568625 393494 568626 393986
rect 569302 393494 569303 393986
rect 568625 393493 569303 393494
rect 569753 393986 570431 393987
rect 569753 393494 569754 393986
rect 570430 393494 570431 393986
rect 570843 393506 570844 393998
rect 571520 393506 571521 393998
rect 571959 393520 571960 394012
rect 572636 393520 572637 394012
rect 571959 393519 572637 393520
rect 570843 393505 571521 393506
rect 569753 393493 570431 393494
rect 571959 393284 572637 393285
rect 570855 393272 571533 393273
rect 569741 393258 570419 393259
rect 568611 393246 569289 393247
rect 567483 393220 568161 393221
rect 567483 392728 567484 393220
rect 568160 392728 568161 393220
rect 568611 392754 568612 393246
rect 569288 392754 569289 393246
rect 569741 392766 569742 393258
rect 570418 392766 570419 393258
rect 570855 392780 570856 393272
rect 571532 392780 571533 393272
rect 571959 392792 571960 393284
rect 572636 392792 572637 393284
rect 571959 392791 572637 392792
rect 570855 392779 571533 392780
rect 569741 392765 570419 392766
rect 568611 392753 569289 392754
rect 567483 392727 568161 392728
rect 570869 392520 571547 392521
rect 569767 392494 570445 392495
rect 568611 392468 569289 392469
rect 567497 392454 568175 392455
rect 567497 391962 567498 392454
rect 568174 391962 568175 392454
rect 568611 391976 568612 392468
rect 569288 391976 569289 392468
rect 569767 392002 569768 392494
rect 570444 392002 570445 392494
rect 570869 392028 570870 392520
rect 571546 392028 571547 392520
rect 570869 392027 571547 392028
rect 571933 392506 572611 392507
rect 571933 392014 571934 392506
rect 572610 392014 572611 392506
rect 571933 392013 572611 392014
rect 569767 392001 570445 392002
rect 568611 391975 569289 391976
rect 567497 391961 568175 391962
rect 513017 374435 560036 377437
rect 491671 371880 492903 371881
rect 491671 371614 491672 371880
rect 492902 371614 492903 371880
rect 491671 371613 492903 371614
rect 491671 371388 492903 371389
rect 491671 371122 491672 371388
rect 492902 371122 492903 371388
rect 491671 371121 492903 371122
rect 491681 370886 492913 370887
rect 491681 370620 491682 370886
rect 492912 370620 492913 370886
rect 491681 370619 492913 370620
rect 491689 370412 492921 370413
rect 491689 370146 491690 370412
rect 492920 370146 492921 370412
rect 491689 370145 492921 370146
rect 491671 369882 492903 369883
rect 491671 369616 491672 369882
rect 492902 369616 492903 369882
rect 491671 369615 492903 369616
rect 491671 369362 492903 369363
rect 491671 369096 491672 369362
rect 492902 369096 492903 369362
rect 491671 369095 492903 369096
rect 491681 368832 492913 368833
rect 491681 368566 491682 368832
rect 492912 368566 492913 368832
rect 491681 368565 492913 368566
rect 491689 368340 492921 368341
rect 491689 368074 491690 368340
rect 492920 368074 492921 368340
rect 491689 368073 492921 368074
rect 491681 367914 492913 367915
rect 491681 367648 491682 367914
rect 491681 367647 492913 367648
rect 491689 367450 492921 367451
rect 491689 367184 491690 367450
rect 492920 367184 492921 367450
rect 491689 367183 492921 367184
rect 513017 362231 515493 374435
rect 537047 371822 538279 371823
rect 537047 371556 537048 371822
rect 538278 371556 538279 371822
rect 537047 371555 538279 371556
rect 537065 371360 538297 371361
rect 537065 371094 537066 371360
rect 538296 371094 538297 371360
rect 537065 371093 538297 371094
rect 537075 370810 538307 370811
rect 537075 370544 537076 370810
rect 538306 370544 538307 370810
rect 537075 370543 538307 370544
rect 537075 370318 538307 370319
rect 537075 370052 537076 370318
rect 538306 370052 538307 370318
rect 537075 370051 538307 370052
rect 537085 369788 538317 369789
rect 537085 369522 537086 369788
rect 538316 369522 538317 369788
rect 537085 369521 538317 369522
rect 537065 369286 538297 369287
rect 537065 369020 537066 369286
rect 538296 369020 538297 369286
rect 537065 369019 538297 369020
rect 537075 368804 538307 368805
rect 537075 368538 537076 368804
rect 538306 368538 538307 368804
rect 537075 368537 538307 368538
rect 537093 368236 538325 368237
rect 537093 367970 537094 368236
rect 538324 367970 538325 368236
rect 537093 367969 538325 367970
rect 537085 367810 538317 367811
rect 537085 367544 537086 367810
rect 538316 367544 538317 367810
rect 537085 367543 538317 367544
rect 537085 367394 538317 367395
rect 537085 367128 537086 367394
rect 538316 367128 538317 367394
rect 537085 367127 538317 367128
rect 513847 361665 515493 362231
rect 551988 355244 560036 374435
rect 569547 371804 571377 371805
rect 567381 371778 569211 371779
rect 567381 370316 567382 371778
rect 569210 370316 569211 371778
rect 569547 370342 569548 371804
rect 571376 370342 571377 371804
rect 569547 370341 571377 370342
rect 571673 371804 573503 371805
rect 571673 370342 571674 371804
rect 573502 370342 573503 371804
rect 571673 370341 573503 370342
rect 567381 370315 569211 370316
rect 571687 370042 573463 370043
rect 569547 370028 571323 370029
rect 567395 369976 569171 369977
rect 567395 369246 567396 369976
rect 569170 369246 569171 369976
rect 569547 369298 569548 370028
rect 571322 369298 571323 370028
rect 571687 369312 571688 370042
rect 573462 369312 573463 370042
rect 571687 369311 573463 369312
rect 569547 369297 571323 369298
rect 567395 369245 569171 369246
rect 571713 368778 573437 368779
rect 569535 368752 571259 368753
rect 567395 368700 569119 368701
rect 567395 367290 567396 368700
rect 569118 367290 569119 368700
rect 569535 367342 569536 368752
rect 571258 367342 571259 368752
rect 571713 367368 571714 368778
rect 573436 367368 573437 368778
rect 571713 367367 573437 367368
rect 569535 367341 571259 367342
rect 567395 367289 569119 367290
rect 573605 357166 573851 357167
rect 567241 356952 567509 356953
rect 567241 356694 567242 356952
rect 567508 356694 567509 356952
rect 573605 356914 573606 357166
rect 573850 356914 573851 357166
rect 573605 356913 573851 356914
rect 567241 356693 567509 356694
rect 551988 355116 559900 355244
rect 560014 355116 560036 355244
rect 573659 355486 573899 355487
rect 573659 355236 573660 355486
rect 573898 355236 573899 355486
rect 573659 355235 573899 355236
rect 551988 355008 560036 355116
rect 551988 354888 559752 355008
rect 559872 354888 560036 355008
rect 521455 311449 523101 311573
rect 491613 305792 492939 305793
rect 491613 305288 491614 305792
rect 492938 305288 492939 305792
rect 491613 305287 492939 305288
rect 491633 304982 492959 304983
rect 491633 304478 491634 304982
rect 492958 304478 492959 304982
rect 491633 304477 492959 304478
rect 491633 304200 492959 304201
rect 491633 303696 491634 304200
rect 492958 303696 492959 304200
rect 491633 303695 492959 303696
rect 491651 303408 492977 303409
rect 491651 302904 491652 303408
rect 492976 302904 492977 303408
rect 491651 302903 492977 302904
rect 491651 302646 492977 302647
rect 491651 302142 491652 302646
rect 492976 302142 492977 302646
rect 491651 302141 492977 302142
rect 491661 301846 492987 301847
rect 491661 301342 491662 301846
rect 492986 301342 492987 301846
rect 491661 301341 492987 301342
rect 521455 297663 523853 311449
rect 551988 310208 560036 354888
rect 573601 311954 573865 311955
rect 567205 311944 567463 311945
rect 567205 311670 567206 311944
rect 567462 311670 567463 311944
rect 573601 311692 573602 311954
rect 573864 311692 573865 311954
rect 573601 311691 573865 311692
rect 567205 311669 567463 311670
rect 551988 310118 559962 310208
rect 560026 310118 560036 310208
rect 551988 309988 560036 310118
rect 573649 310278 573895 310279
rect 573649 310034 573650 310278
rect 573894 310034 573895 310278
rect 573649 310033 573895 310034
rect 551988 309868 559764 309988
rect 559884 309868 560036 309988
rect 536987 305756 538313 305757
rect 536987 305252 536988 305756
rect 538312 305252 538313 305756
rect 536987 305251 538313 305252
rect 536987 304934 538313 304935
rect 536987 304430 536988 304934
rect 538312 304430 538313 304934
rect 536987 304429 538313 304430
rect 537025 304132 538351 304133
rect 537025 303628 537026 304132
rect 538350 303628 538351 304132
rect 537025 303627 538351 303628
rect 537025 303350 538351 303351
rect 537025 302846 537026 303350
rect 538350 302846 538351 303350
rect 537025 302845 538351 302846
rect 537025 302566 538351 302567
rect 537025 302062 537026 302566
rect 538350 302062 538351 302566
rect 537025 302061 538351 302062
rect 537025 301708 538351 301709
rect 537025 301204 537026 301708
rect 538350 301204 538351 301708
rect 537025 301203 538351 301204
rect 551988 297663 560036 309868
rect 567401 305824 569125 305825
rect 567401 304414 567402 305824
rect 569124 304414 569125 305824
rect 567401 304413 569125 304414
rect 569487 305824 571211 305825
rect 569487 304414 569488 305824
rect 571210 304414 571211 305824
rect 569487 304413 571211 304414
rect 571509 305824 573233 305825
rect 571509 304414 571510 305824
rect 573232 304414 573233 305824
rect 571509 304413 573233 304414
rect 571483 304184 573207 304185
rect 569487 304132 571211 304133
rect 567413 304092 569137 304093
rect 567413 302682 567414 304092
rect 569136 302682 569137 304092
rect 569487 302722 569488 304132
rect 571210 302722 571211 304132
rect 571483 302774 571484 304184
rect 573206 302774 573207 304184
rect 571483 302773 573207 302774
rect 569487 302721 571211 302722
rect 567413 302681 569137 302682
rect 571535 302452 573259 302453
rect 569461 302412 571185 302413
rect 567439 302400 569163 302401
rect 567439 300990 567440 302400
rect 569162 300990 569163 302400
rect 569461 301002 569462 302412
rect 571184 301002 571185 302412
rect 571535 301042 571536 302452
rect 573258 301042 573259 302452
rect 571535 301041 573259 301042
rect 569461 301001 571185 301002
rect 567439 300989 569163 300990
rect 521455 296157 560036 297663
rect 521379 294511 560036 296157
rect 551988 154943 560036 294511
<< via4 >>
rect 567370 640173 573686 644249
rect 567370 630105 573686 634181
rect 573628 581122 573910 581438
rect 566918 564368 574066 571176
rect 573616 507620 573914 507912
rect 487194 471134 487810 471788
rect 488088 471160 488704 471814
rect 535652 471358 536268 472012
rect 536478 471358 537094 472012
rect 487194 469934 487810 470588
rect 488088 469960 488704 470614
rect 535652 470158 536268 470812
rect 536478 470158 537094 470812
rect 487194 468734 487810 469388
rect 488088 468760 488704 469414
rect 535652 468958 536268 469612
rect 536478 468958 537094 469612
rect 487194 467534 487810 468188
rect 488088 467560 488704 468214
rect 535652 467758 536268 468412
rect 536478 467758 537094 468412
rect 487194 466334 487810 466988
rect 488088 466360 488704 467014
rect 535652 466558 536268 467212
rect 536478 466558 537094 467212
rect 566954 465896 574254 472368
rect 567262 446548 567506 446796
rect 573574 446348 573832 446592
rect 573592 444642 573890 444908
rect 567274 403278 567518 403520
rect 573592 403352 573842 403624
rect 573648 401658 573884 401912
rect 487244 393598 487754 394104
rect 488026 393606 488536 394112
rect 535658 393688 536176 394020
rect 536458 393728 536976 394060
rect 487244 392998 487754 393504
rect 488026 393006 488536 393512
rect 535658 393188 536176 393520
rect 536458 393228 536976 393560
rect 487244 392398 487754 392904
rect 488026 392406 488536 392912
rect 535658 392688 536176 393020
rect 536458 392728 536976 393060
rect 487244 391798 487754 392304
rect 488026 391806 488536 392312
rect 535658 392188 536176 392520
rect 536458 392228 536976 392560
rect 535658 391688 536176 392020
rect 536458 391728 536976 392060
rect 567458 393494 568134 393986
rect 568626 393494 569302 393986
rect 569754 393494 570430 393986
rect 570844 393506 571520 393998
rect 571960 393520 572636 394012
rect 567484 392728 568160 393220
rect 568612 392754 569288 393246
rect 569742 392766 570418 393258
rect 570856 392780 571532 393272
rect 571960 392792 572636 393284
rect 567498 391962 568174 392454
rect 568612 391976 569288 392468
rect 569768 392002 570444 392494
rect 570870 392028 571546 392520
rect 571934 392014 572610 392506
rect 491672 371614 492902 371880
rect 491672 371122 492902 371388
rect 491682 370620 492912 370886
rect 491690 370146 492920 370412
rect 491672 369616 492902 369882
rect 491672 369096 492902 369362
rect 491682 368566 492912 368832
rect 491690 368074 492920 368340
rect 491690 367648 492912 367914
rect 492912 367648 492920 367914
rect 491690 367184 492920 367450
rect 537048 371556 538278 371822
rect 537066 371094 538296 371360
rect 537076 370544 538306 370810
rect 537076 370052 538306 370318
rect 537086 369522 538316 369788
rect 537066 369020 538296 369286
rect 537076 368538 538306 368804
rect 537094 367970 538324 368236
rect 537086 367544 538316 367810
rect 537086 367128 538316 367394
rect 567382 370316 569210 371778
rect 569548 370342 571376 371804
rect 571674 370342 573502 371804
rect 567396 369246 569170 369976
rect 569548 369298 571322 370028
rect 571688 369312 573462 370042
rect 567396 367290 569118 368700
rect 569536 367342 571258 368752
rect 571714 367368 573436 368778
rect 567242 356694 567508 356952
rect 573606 356914 573850 357166
rect 573660 355236 573898 355486
rect 491614 305288 492938 305792
rect 491634 304478 492958 304982
rect 491634 303696 492958 304200
rect 491652 302904 492976 303408
rect 491652 302142 492976 302646
rect 491662 301342 492986 301846
rect 567206 311670 567462 311944
rect 573602 311692 573864 311954
rect 573650 310034 573894 310278
rect 536988 305252 538312 305756
rect 536988 304430 538312 304934
rect 537026 303628 538350 304132
rect 537026 302846 538350 303350
rect 537026 302062 538350 302566
rect 537026 301204 538350 301708
rect 567402 304414 569124 305824
rect 569488 304414 571210 305824
rect 571510 304414 573232 305824
rect 567414 302682 569136 304092
rect 569488 302722 571210 304132
rect 571484 302774 573206 304184
rect 567440 300990 569162 302400
rect 569462 301002 571184 302412
rect 571536 301042 573258 302452
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 395311 691057 573934 697819
rect 567172 644249 573934 691057
rect 567172 640173 567370 644249
rect 573686 640173 573934 644249
rect 567172 634181 573934 640173
rect 567172 630105 567370 634181
rect 573686 630105 573934 634181
rect 567172 627323 573934 630105
rect 567170 621961 573956 627323
rect 567172 581438 573934 621961
rect 567172 581122 573628 581438
rect 573910 581122 573934 581438
rect 567172 571200 573934 581122
rect 566894 571176 574090 571200
rect 566894 564368 566918 571176
rect 574066 564368 574090 571176
rect 566894 564344 574090 564368
rect 567172 507936 573934 564344
rect 567172 507912 573938 507936
rect 567172 507620 573616 507912
rect 573914 507620 573938 507912
rect 567172 507596 573938 507620
rect 567172 472392 573934 507596
rect 566930 472368 574278 472392
rect 487136 471814 488768 472104
rect 487136 471788 488088 471814
rect 487136 471134 487194 471788
rect 487810 471160 488088 471788
rect 488704 471160 488768 471814
rect 487810 471134 488768 471160
rect 487136 470614 488768 471134
rect 487136 470588 488088 470614
rect 487136 469934 487194 470588
rect 487810 469960 488088 470588
rect 488704 469960 488768 470614
rect 487810 469934 488768 469960
rect 487136 469414 488768 469934
rect 487136 469388 488088 469414
rect 487136 468734 487194 469388
rect 487810 468760 488088 469388
rect 488704 468760 488768 469414
rect 487810 468734 488768 468760
rect 487136 468214 488768 468734
rect 487136 468188 488088 468214
rect 487136 467534 487194 468188
rect 487810 467560 488088 468188
rect 488704 467560 488768 468214
rect 487810 467534 488768 467560
rect 487136 467014 488768 467534
rect 487136 466988 488088 467014
rect 487136 466334 487194 466988
rect 487810 466360 488088 466988
rect 488704 466360 488768 467014
rect 487810 466334 488768 466360
rect 487136 452232 488768 466334
rect 535520 472012 537152 472260
rect 535520 471358 535652 472012
rect 536268 471358 536478 472012
rect 537094 471358 537152 472012
rect 535520 470812 537152 471358
rect 535520 470158 535652 470812
rect 536268 470158 536478 470812
rect 537094 470158 537152 470812
rect 535520 469612 537152 470158
rect 535520 468958 535652 469612
rect 536268 468958 536478 469612
rect 537094 468958 537152 469612
rect 535520 468412 537152 468958
rect 535520 467758 535652 468412
rect 536268 467758 536478 468412
rect 537094 467758 537152 468412
rect 535520 467212 537152 467758
rect 535520 466558 535652 467212
rect 536268 466558 536478 467212
rect 537094 466558 537152 467212
rect 535520 454082 537152 466558
rect 566930 465896 566954 472368
rect 574254 465896 574278 472368
rect 566930 465872 574278 465896
rect 567172 446796 573934 465872
rect 567172 446548 567262 446796
rect 567506 446592 573934 446796
rect 567506 446548 573574 446592
rect 567172 446348 573574 446548
rect 573832 446348 573934 446592
rect 567172 445694 573934 446348
rect 567148 444908 573934 445694
rect 567148 444696 573592 444908
rect 567172 444642 573592 444696
rect 573890 444642 573934 444908
rect 567172 403624 573934 444642
rect 567172 403520 573592 403624
rect 567172 403278 567274 403520
rect 567518 403352 573592 403520
rect 573842 403352 573934 403624
rect 567518 403278 573934 403352
rect 567172 401912 573934 403278
rect 567172 401658 573648 401912
rect 573884 401658 573934 401912
rect 487136 394112 488768 398834
rect 487136 394104 488026 394112
rect 487136 393598 487244 394104
rect 487754 393606 488026 394104
rect 488536 393606 488768 394112
rect 487754 393598 488768 393606
rect 487136 393512 488768 393598
rect 487136 393504 488026 393512
rect 487136 392998 487244 393504
rect 487754 393006 488026 393504
rect 488536 393006 488768 393512
rect 487754 392998 488768 393006
rect 487136 392912 488768 392998
rect 487136 392904 488026 392912
rect 487136 392398 487244 392904
rect 487754 392406 488026 392904
rect 488536 392406 488768 392912
rect 487754 392398 488768 392406
rect 487136 392312 488768 392398
rect 487136 392304 488026 392312
rect 487136 391798 487244 392304
rect 487754 391806 488026 392304
rect 488536 391806 488768 392312
rect 487754 391798 488768 391806
rect 487136 390586 488768 391798
rect 535520 394060 537152 398834
rect 535520 394020 536458 394060
rect 535520 393688 535658 394020
rect 536176 393728 536458 394020
rect 536976 393728 537152 394060
rect 536176 393688 537152 393728
rect 535520 393560 537152 393688
rect 535520 393520 536458 393560
rect 535520 393188 535658 393520
rect 536176 393228 536458 393520
rect 536976 393228 537152 393560
rect 536176 393188 537152 393228
rect 535520 393060 537152 393188
rect 535520 393020 536458 393060
rect 535520 392688 535658 393020
rect 536176 392728 536458 393020
rect 536976 392728 537152 393060
rect 536176 392688 537152 392728
rect 535520 392560 537152 392688
rect 535520 392520 536458 392560
rect 535520 392188 535658 392520
rect 536176 392228 536458 392520
rect 536976 392228 537152 392560
rect 536176 392188 537152 392228
rect 535520 392060 537152 392188
rect 535520 392020 536458 392060
rect 535520 391688 535658 392020
rect 536176 391728 536458 392020
rect 536976 391728 537152 392060
rect 536176 391688 537152 391728
rect 535520 390820 537152 391688
rect 567172 394012 573934 401658
rect 567172 393998 571960 394012
rect 567172 393986 570844 393998
rect 567172 393494 567458 393986
rect 568134 393494 568626 393986
rect 569302 393494 569754 393986
rect 570430 393506 570844 393986
rect 571520 393520 571960 393998
rect 572636 393520 573934 394012
rect 571520 393506 573934 393520
rect 570430 393494 573934 393506
rect 567172 393284 573934 393494
rect 567172 393272 571960 393284
rect 567172 393258 570856 393272
rect 567172 393246 569742 393258
rect 567172 393220 568612 393246
rect 567172 392728 567484 393220
rect 568160 392754 568612 393220
rect 569288 392766 569742 393246
rect 570418 392780 570856 393258
rect 571532 392792 571960 393272
rect 572636 392792 573934 393284
rect 571532 392780 573934 392792
rect 570418 392766 573934 392780
rect 569288 392754 573934 392766
rect 568160 392728 573934 392754
rect 567172 392520 573934 392728
rect 567172 392494 570870 392520
rect 567172 392468 569768 392494
rect 567172 392454 568612 392468
rect 567172 391962 567498 392454
rect 568174 391976 568612 392454
rect 569288 392002 569768 392468
rect 570444 392028 570870 392494
rect 571546 392506 573934 392520
rect 571546 392028 571934 392506
rect 570444 392014 571934 392028
rect 572610 392014 573934 392506
rect 570444 392002 573934 392014
rect 569288 391976 573934 392002
rect 568174 391962 573934 391976
rect 491505 371880 493151 372089
rect 491505 371614 491672 371880
rect 492902 371614 493151 371880
rect 491505 371388 493151 371614
rect 491505 371122 491672 371388
rect 492902 371122 493151 371388
rect 491505 370886 493151 371122
rect 491505 370620 491682 370886
rect 492912 370620 493151 370886
rect 491505 370412 493151 370620
rect 491505 370146 491690 370412
rect 492920 370146 493151 370412
rect 491505 369882 493151 370146
rect 491505 369616 491672 369882
rect 492902 369616 493151 369882
rect 491505 369362 493151 369616
rect 491505 369096 491672 369362
rect 492902 369096 493151 369362
rect 491505 368832 493151 369096
rect 491505 368566 491682 368832
rect 492912 368566 493151 368832
rect 491505 368340 493151 368566
rect 491505 368074 491690 368340
rect 492920 368074 493151 368340
rect 491505 367914 493151 368074
rect 491505 367648 491690 367914
rect 492920 367648 493151 367914
rect 491505 367450 493151 367648
rect 491505 367184 491690 367450
rect 492920 367184 493151 367450
rect 491505 354925 493151 367184
rect 536869 371822 538515 372013
rect 536869 371556 537048 371822
rect 538278 371556 538515 371822
rect 536869 371360 538515 371556
rect 536869 371094 537066 371360
rect 538296 371094 538515 371360
rect 536869 370810 538515 371094
rect 536869 370544 537076 370810
rect 538306 370544 538515 370810
rect 536869 370318 538515 370544
rect 536869 370052 537076 370318
rect 538306 370052 538515 370318
rect 536869 369788 538515 370052
rect 536869 369522 537086 369788
rect 538316 369522 538515 369788
rect 536869 369286 538515 369522
rect 536869 369020 537066 369286
rect 538296 369020 538515 369286
rect 536869 368804 538515 369020
rect 536869 368538 537076 368804
rect 538306 368538 538515 368804
rect 536869 368236 538515 368538
rect 536869 367970 537094 368236
rect 538324 367970 538515 368236
rect 536869 367810 538515 367970
rect 536869 367544 537086 367810
rect 538316 367544 538515 367810
rect 536869 367394 538515 367544
rect 536869 367128 537086 367394
rect 538316 367128 538515 367394
rect 536869 355301 538515 367128
rect 567172 371804 573934 391962
rect 567172 371778 569548 371804
rect 567172 370316 567382 371778
rect 569210 370342 569548 371778
rect 571376 370342 571674 371804
rect 573502 370342 573934 371804
rect 569210 370316 573934 370342
rect 567172 370042 573934 370316
rect 567172 370028 571688 370042
rect 567172 369976 569548 370028
rect 567172 369246 567396 369976
rect 569170 369298 569548 369976
rect 571322 369312 571688 370028
rect 573462 369312 573934 370042
rect 571322 369298 573934 369312
rect 569170 369246 573934 369298
rect 567172 368778 573934 369246
rect 567172 368752 571714 368778
rect 567172 368700 569536 368752
rect 567172 367290 567396 368700
rect 569118 367342 569536 368700
rect 571258 367368 571714 368752
rect 573436 367368 573934 368778
rect 571258 367342 573934 367368
rect 569118 367290 573934 367342
rect 567172 357166 573934 367290
rect 567172 356952 573606 357166
rect 567172 356694 567242 356952
rect 567508 356914 573606 356952
rect 573850 356914 573934 357166
rect 567508 356694 573934 356914
rect 567172 355486 573934 356694
rect 567172 355236 573660 355486
rect 573898 355236 573934 355486
rect 491505 305792 493151 317777
rect 491505 305288 491614 305792
rect 492938 305288 493151 305792
rect 491505 304982 493151 305288
rect 491505 304478 491634 304982
rect 492958 304478 493151 304982
rect 491505 304200 493151 304478
rect 491505 303696 491634 304200
rect 492958 303696 493151 304200
rect 491505 303408 493151 303696
rect 491505 302904 491652 303408
rect 492976 302904 493151 303408
rect 491505 302646 493151 302904
rect 491505 302142 491652 302646
rect 492976 302142 493151 302646
rect 491505 301846 493151 302142
rect 491505 301342 491662 301846
rect 492986 301342 493151 301846
rect 491505 300799 493151 301342
rect 536869 305756 538515 317173
rect 536869 305252 536988 305756
rect 538312 305252 538515 305756
rect 536869 304934 538515 305252
rect 536869 304430 536988 304934
rect 538312 304430 538515 304934
rect 536869 304132 538515 304430
rect 536869 303628 537026 304132
rect 538350 303628 538515 304132
rect 536869 303350 538515 303628
rect 536869 302846 537026 303350
rect 538350 302846 538515 303350
rect 536869 302566 538515 302846
rect 536869 302062 537026 302566
rect 538350 302062 538515 302566
rect 536869 301708 538515 302062
rect 536869 301204 537026 301708
rect 538350 301204 538515 301708
rect 536869 300571 538515 301204
rect 567172 311954 573934 355236
rect 567172 311944 573602 311954
rect 567172 311670 567206 311944
rect 567462 311692 573602 311944
rect 573864 311692 573934 311954
rect 567462 311670 573934 311692
rect 567172 310278 573934 311670
rect 567172 310034 573650 310278
rect 573894 310034 573934 310278
rect 567172 305824 573934 310034
rect 567172 304414 567402 305824
rect 569124 304414 569488 305824
rect 571210 304414 571510 305824
rect 573232 304414 573934 305824
rect 567172 304184 573934 304414
rect 567172 304132 571484 304184
rect 567172 304092 569488 304132
rect 567172 302682 567414 304092
rect 569136 302722 569488 304092
rect 571210 302774 571484 304132
rect 573206 302774 573934 304184
rect 571210 302722 573934 302774
rect 569136 302682 573934 302722
rect 567172 302452 573934 302682
rect 567172 302412 571536 302452
rect 567172 302400 569462 302412
rect 567172 300990 567440 302400
rect 569162 301002 569462 302400
rect 571184 301042 571536 302412
rect 573258 301042 573934 302452
rect 571184 301002 573934 301042
rect 569162 300990 573934 301002
rect 567172 147394 573934 300990
use bandgaptop_flat_io  bandgaptop_flat_io_0
timestamp 1656304949
transform 0 1 -129800 -1 0 972356
box 422960 603262 497922 669400
use bgr_gen7  bgr_gen7_0
timestamp 1656306043
transform 0 -1 541413 -1 0 363861
box -205 -1505 55275 53897
use bgr_top  bgr_top_0
timestamp 1656306043
transform 0 1 483840 -1 0 455714
box 0 0 58512 56576
use nmos_flat  nmos_flat_0
timestamp 1655700407
transform -1 0 563187 0 1 355948
box -2706 -1060 2635 940
use nmos_flat  nmos_flat_1
timestamp 1655700407
transform -1 0 563141 0 1 310928
box -2706 -1060 2635 940
use nmos_flat  nmos_flat_2
timestamp 1655700407
transform -1 0 563523 0 1 402518
box -2706 -1060 2635 940
use nmos_flat  nmos_flat_3
timestamp 1655700407
transform -1 0 563173 0 1 445778
box -2706 -1060 2635 940
use nmos_flat  nmos_flat_4
timestamp 1655700407
transform -1 0 563375 0 1 582166
box -2706 -1060 2635 940
use nmos_flat  nmos_flat_5
timestamp 1655700407
transform -1 0 563303 0 1 508484
box -2706 -1060 2635 940
use pmos_flat  pmos_flat_0
timestamp 1655503347
transform -1 0 577157 0 1 445592
box -2742 -1060 2645 940
use pmos_flat  pmos_flat_1
timestamp 1655503347
transform -1 0 577161 0 1 402608
box -2742 -1060 2645 940
use pmos_flat  pmos_flat_2
timestamp 1655503347
transform -1 0 577057 0 1 356166
box -2742 -1060 2645 940
use pmos_flat  pmos_flat_3
timestamp 1655503347
transform -1 0 577077 0 1 310954
box -2742 -1060 2645 940
use pmos_flat  pmos_flat_4
timestamp 1655503347
transform -1 0 577171 0 1 582062
box -2742 -1060 2645 940
use pmos_flat  pmos_flat_5
timestamp 1655503347
transform -1 0 577403 0 1 508572
box -2742 -1060 2645 940
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 41 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 42 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 43 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 44 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 45 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 46 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 47 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 48 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 49 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 50 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 51 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 52 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 53 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 54 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 55 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 56 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 57 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 58 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 59 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 60 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 61 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 62 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 63 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 64 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 65 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 66 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 67 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 68 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 69 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 70 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 71 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 72 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 73 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 74 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 75 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 76 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 77 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 78 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 79 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 80 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 81 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 85 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 86 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 87 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 88 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 89 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 90 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 91 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 92 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 93 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 94 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 95 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 96 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 97 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 98 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 99 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 100 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 101 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 102 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 103 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 104 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 105 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 106 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 107 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 108 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 109 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 110 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 111 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 112 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 113 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 114 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 115 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 116 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 117 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 118 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 119 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 120 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 121 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 122 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 123 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 124 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 125 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 126 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 127 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 128 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 129 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 130 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 131 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 132 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 133 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 134 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 135 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 136 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 137 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 138 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 139 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 140 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 141 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 142 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 143 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 144 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 145 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 146 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 147 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 148 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 149 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 150 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 151 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 152 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 153 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 154 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 155 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 156 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 157 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 158 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 159 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 160 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 161 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 162 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 163 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 164 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 165 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 166 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 167 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 168 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 169 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 170 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 171 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 172 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 173 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 174 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 175 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 176 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 177 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 178 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 179 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 180 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 181 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 182 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 183 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 184 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 185 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 186 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 187 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 188 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 189 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 190 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 191 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 192 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 193 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 194 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 195 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 196 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 197 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 198 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 199 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 200 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 201 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 202 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 203 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 204 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 205 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 206 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 207 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 208 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 209 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 210 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 211 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 212 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 213 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 214 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 215 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 216 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 217 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 218 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 219 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 220 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 221 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 222 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 223 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 224 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 225 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 226 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 227 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 228 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 229 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 230 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 231 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 232 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 233 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 234 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 235 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 236 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 237 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 238 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 239 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 240 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 241 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 242 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 243 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 244 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 245 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 246 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 247 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 248 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 249 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 250 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 251 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 252 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 253 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 254 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 255 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 256 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 257 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 258 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 259 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 260 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 261 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 262 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 263 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 264 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 265 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 266 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 267 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 268 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 269 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 270 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 271 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 272 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 273 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 274 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 275 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 276 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 277 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 278 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 279 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 280 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 281 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 282 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 283 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 284 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 285 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 286 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 287 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 288 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 289 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 290 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 291 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 292 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 293 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 294 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 295 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 296 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 297 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 298 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 299 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 300 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 301 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 302 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 303 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 304 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 305 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 306 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 307 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 308 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 309 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 310 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 311 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 312 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 313 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 314 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 315 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 316 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 317 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 318 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 319 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 320 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 321 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 322 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 323 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 324 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 325 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 326 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 327 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 328 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 329 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 330 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 331 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 332 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 333 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 334 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 335 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 336 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 337 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 338 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 339 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 340 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 341 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 342 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 343 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 344 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 345 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 346 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 347 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 348 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 349 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 350 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 351 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 352 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 353 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 354 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 355 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 356 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 357 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 358 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 359 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 360 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 361 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 362 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 363 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 364 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 365 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 366 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 367 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 368 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 369 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 370 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 371 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 372 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 373 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 374 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 375 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 376 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 377 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 378 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 379 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 380 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 381 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 382 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 383 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 384 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 385 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 386 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 387 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 388 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 389 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 390 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 391 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 392 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 393 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 394 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 395 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 396 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 397 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 398 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 399 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 400 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 401 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 402 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 403 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 404 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 405 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 406 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 407 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 408 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 409 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 410 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 411 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 412 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 413 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 414 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 415 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 416 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 417 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 418 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 419 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 420 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 421 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 422 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 423 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 424 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 425 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 426 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 427 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 428 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 429 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 430 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 431 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 432 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 433 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 434 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 435 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 436 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 437 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 438 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 439 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 440 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 441 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 442 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 443 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 444 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 445 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 446 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 447 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 448 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 449 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 450 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 451 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 452 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 453 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 454 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 455 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 456 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 457 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 458 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 459 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 460 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 461 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 462 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 463 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 464 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 465 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 466 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 467 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 468 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 469 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 470 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 471 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 472 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 473 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 474 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 475 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 476 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 477 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 478 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 479 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 480 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 481 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 482 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 483 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 484 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 485 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 486 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 487 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 488 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 489 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 490 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 491 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 492 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 493 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 494 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 495 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 496 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 497 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 498 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 499 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 500 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 501 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 502 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 503 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 504 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 505 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 506 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 507 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 508 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 509 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 510 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 511 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 512 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 513 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 514 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 515 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 516 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 517 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 518 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 519 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 520 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 521 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 522 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 523 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 524 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 525 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 526 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 527 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 528 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 529 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 530 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 531 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 532 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 533 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 534 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 535 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 536 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 537 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 538 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 539 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 540 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 541 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 542 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 543 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 544 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 545 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 546 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 547 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 548 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 549 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 550 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 551 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 552 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 553 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 554 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 555 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 556 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 557 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 558 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 559 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 560 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 561 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 562 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 563 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 564 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 565 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 566 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 567 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 568 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 569 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 570 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 571 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 572 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 573 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 574 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 575 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 576 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 577 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 578 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 579 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 580 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 581 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 582 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 583 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 584 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 585 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 586 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 587 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 588 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 589 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 590 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 590 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 591 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 591 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 592 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 592 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 592 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 592 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 593 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 593 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 594 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 594 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 594 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 594 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 595 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 595 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 596 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 596 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 597 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 597 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 598 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 599 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 600 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 601 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 602 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 603 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 604 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 605 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 606 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 607 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 608 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 609 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 610 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 611 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 612 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 613 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 614 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 615 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 616 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 617 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 618 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 619 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 620 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 621 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 622 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 623 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 624 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 625 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 626 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 627 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 628 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 629 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 630 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 631 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 632 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 633 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 634 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 635 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 636 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 637 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 638 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 639 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 640 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 641 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 642 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 643 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 644 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 645 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 646 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 647 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 648 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 649 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 650 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 651 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 652 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 653 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 654 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 655 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 656 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 657 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 658 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 659 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 660 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 661 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 662 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 663 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 664 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 665 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 666 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 667 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 668 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 669 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 670 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 671 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 672 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 673 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 674 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 675 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 676 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 677 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 678 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 679 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 680 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 681 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 682 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 683 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 684 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 685 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 686 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 687 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 688 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 689 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 690 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 691 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 692 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 693 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 694 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 695 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 696 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 697 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 698 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 699 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 700 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 701 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 702 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 703 nsew
<< end >>
