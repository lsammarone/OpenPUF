magic
tech sky130A
timestamp 1656729169
<< metal2 >>
rect -90 74 90 90
rect -90 -74 -74 74
rect 74 -74 90 74
rect -90 -90 90 -74
<< via2 >>
rect -74 -74 74 74
<< metal3 >>
rect -90 74 90 90
rect -90 -74 -74 74
rect 74 -74 90 74
rect -90 -90 90 -74
<< properties >>
string GDS_END 9349174
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/merge/design_merged.gds
string GDS_START 9348018
<< end >>
