magic
tech sky130A
timestamp 1655322987
<< metal4 >>
rect -500 379 500 455
rect -500 -379 -459 379
rect 459 -379 500 379
rect -500 -455 500 -379
<< via4 >>
rect -459 -379 459 379
<< metal5 >>
rect -500 379 500 455
rect -500 -379 -459 379
rect 459 -379 500 379
rect -500 -455 500 -379
<< end >>
