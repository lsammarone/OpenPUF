magic
tech sky130A
magscale 1 2
timestamp 1655322987
<< nwell >>
rect 33027 4847 33405 5966
rect 32760 4818 33405 4847
rect 32760 4526 33296 4818
rect 17040 4150 17422 4471
rect 47182 4310 47564 4631
<< nsubdiff >>
rect 47307 4483 47441 4502
rect 47307 4449 47379 4483
rect 47413 4449 47441 4483
rect 47307 4432 47441 4449
rect 17165 4323 17299 4342
rect 17165 4289 17237 4323
rect 17271 4289 17299 4323
rect 17165 4272 17299 4289
<< nsubdiffcont >>
rect 47379 4449 47413 4483
rect 17237 4289 17271 4323
<< locali >>
rect 32002 4524 32358 4530
rect 32002 4490 32049 4524
rect 32083 4490 32137 4524
rect 32171 4490 32358 4524
rect 32002 4480 32358 4490
rect 47104 4483 47647 4503
rect 47104 4449 47379 4483
rect 47413 4449 47647 4483
rect 47104 4431 47647 4449
rect 45973 4409 46007 4415
rect 45805 4402 45839 4408
rect 46309 4411 46343 4417
rect 45973 4370 46007 4375
rect 46141 4399 46175 4405
rect 45805 4363 45839 4368
rect 46309 4372 46343 4377
rect 46475 4409 46509 4415
rect 46475 4370 46509 4375
rect 46641 4411 46675 4417
rect 46641 4372 46675 4377
rect 46809 4411 46843 4417
rect 46809 4372 46843 4377
rect 46983 4409 47017 4415
rect 46983 4370 47017 4375
rect 47739 4403 47773 4409
rect 46141 4360 46175 4365
rect 47739 4364 47773 4369
rect 47901 4407 47935 4413
rect 47901 4368 47935 4373
rect 48071 4411 48105 4417
rect 48071 4372 48105 4377
rect 48235 4407 48269 4413
rect 48235 4368 48269 4373
rect 48405 4407 48439 4413
rect 48405 4368 48439 4373
rect 48573 4403 48607 4409
rect 48573 4364 48607 4369
rect 48741 4407 48775 4413
rect 48741 4368 48775 4373
rect 48915 4403 48949 4409
rect 48915 4364 48949 4369
rect 16962 4323 17505 4343
rect 16962 4289 17237 4323
rect 17271 4289 17505 4323
rect 16962 4271 17505 4289
rect 15831 4249 15865 4255
rect 15663 4242 15697 4248
rect 16167 4251 16201 4257
rect 15831 4210 15865 4215
rect 15999 4239 16033 4245
rect 15663 4203 15697 4208
rect 16167 4212 16201 4217
rect 16333 4249 16367 4255
rect 16333 4210 16367 4215
rect 16499 4251 16533 4257
rect 16499 4212 16533 4217
rect 16667 4251 16701 4257
rect 16667 4212 16701 4217
rect 16841 4249 16875 4255
rect 16841 4210 16875 4215
rect 17597 4243 17631 4249
rect 15999 4200 16033 4205
rect 17597 4204 17631 4209
rect 17759 4247 17793 4253
rect 17759 4208 17793 4213
rect 17929 4251 17963 4257
rect 17929 4212 17963 4217
rect 18093 4247 18127 4253
rect 18093 4208 18127 4213
rect 18263 4247 18297 4253
rect 18263 4208 18297 4213
rect 18431 4243 18465 4249
rect 18431 4204 18465 4209
rect 18599 4247 18633 4253
rect 18599 4208 18633 4213
rect 18773 4243 18807 4249
rect 18773 4204 18807 4209
<< viali >>
rect 32049 4490 32083 4524
rect 32137 4490 32171 4524
rect 32714 4522 32748 4556
rect 32985 4486 33019 4520
rect 33073 4486 33107 4520
rect 33161 4486 33195 4520
rect 33249 4486 33283 4520
rect 33337 4486 33371 4520
rect 33425 4486 33459 4520
rect 33513 4486 33547 4520
rect 33601 4486 33635 4520
rect 32714 4442 32748 4476
rect 33339 4384 33373 4418
rect 33505 4380 33539 4414
rect 33673 4386 33707 4420
rect 33840 4384 33874 4418
rect 34010 4385 34044 4419
rect 34174 4386 34208 4420
rect 45805 4368 45839 4402
rect 45973 4375 46007 4409
rect 46141 4365 46175 4399
rect 46309 4377 46343 4411
rect 46475 4375 46509 4409
rect 46641 4377 46675 4411
rect 46809 4377 46843 4411
rect 46983 4375 47017 4409
rect 47739 4369 47773 4403
rect 47901 4373 47935 4407
rect 48071 4377 48105 4411
rect 48235 4373 48269 4407
rect 48405 4373 48439 4407
rect 48573 4369 48607 4403
rect 48741 4373 48775 4407
rect 48915 4369 48949 4403
rect 46005 4272 46039 4306
rect 46105 4272 46139 4306
rect 46205 4272 46239 4306
rect 46305 4272 46339 4306
rect 46405 4272 46439 4306
rect 46505 4272 46539 4306
rect 46605 4272 46639 4306
rect 46705 4272 46739 4306
rect 47665 4272 47699 4306
rect 47765 4272 47799 4306
rect 47865 4272 47899 4306
rect 47965 4272 47999 4306
rect 48065 4272 48099 4306
rect 48165 4272 48199 4306
rect 48265 4272 48299 4306
rect 48365 4272 48399 4306
rect 15663 4208 15697 4242
rect 15831 4215 15865 4249
rect 15999 4205 16033 4239
rect 16167 4217 16201 4251
rect 16333 4215 16367 4249
rect 16499 4217 16533 4251
rect 16667 4217 16701 4251
rect 16841 4215 16875 4249
rect 17597 4209 17631 4243
rect 17759 4213 17793 4247
rect 17929 4217 17963 4251
rect 18093 4213 18127 4247
rect 18263 4213 18297 4247
rect 18431 4209 18465 4243
rect 18599 4213 18633 4247
rect 18773 4209 18807 4243
rect 15863 4112 15897 4146
rect 15963 4112 15997 4146
rect 16063 4112 16097 4146
rect 16163 4112 16197 4146
rect 16263 4112 16297 4146
rect 16363 4112 16397 4146
rect 16463 4112 16497 4146
rect 16563 4112 16597 4146
rect 17523 4112 17557 4146
rect 17623 4112 17657 4146
rect 17723 4112 17757 4146
rect 17823 4112 17857 4146
rect 17923 4112 17957 4146
rect 18023 4112 18057 4146
rect 18123 4112 18157 4146
rect 18223 4112 18257 4146
<< metal1 >>
rect 16714 5441 16969 5797
rect 32650 5464 32984 5788
rect 16714 5389 16734 5441
rect 16786 5389 16812 5441
rect 16864 5389 16905 5441
rect 16957 5389 16969 5441
rect 16714 5359 16969 5389
rect 32650 5412 32693 5464
rect 32745 5412 32806 5464
rect 32858 5412 32907 5464
rect 32959 5412 32984 5464
rect 32650 5368 32984 5412
rect 46854 5441 47081 5809
rect 46854 5389 46885 5441
rect 46937 5389 46968 5441
rect 47020 5389 47081 5441
rect 46854 5355 47081 5389
rect 9370 5224 9906 5308
rect 24404 5233 25012 5291
rect 39508 5241 40132 5299
rect 54514 5247 55247 5305
rect 32778 4844 32886 4857
rect 32778 4792 32808 4844
rect 32860 4792 32886 4844
rect 32778 4761 32886 4792
rect 34318 4761 34353 4857
rect 1 4690 19384 4691
rect 0 4626 19384 4690
rect 1 4625 19384 4626
rect 19318 4539 19384 4625
rect 47023 4617 47690 4626
rect 32699 4556 32778 4584
rect 47033 4568 47690 4617
rect 19318 4524 32265 4539
rect 19318 4490 32049 4524
rect 32083 4490 32137 4524
rect 32171 4490 32265 4524
rect 19318 4473 32265 4490
rect 32699 4522 32714 4556
rect 32748 4528 32778 4556
rect 32748 4522 33697 4528
rect 32699 4520 33697 4522
rect 32699 4486 32985 4520
rect 33019 4486 33073 4520
rect 33107 4486 33161 4520
rect 33195 4486 33249 4520
rect 33283 4486 33337 4520
rect 33371 4486 33425 4520
rect 33459 4486 33513 4520
rect 33547 4486 33601 4520
rect 33635 4486 33697 4520
rect 32699 4480 33697 4486
rect 32699 4476 32781 4480
rect 16933 4412 17582 4462
rect 32699 4442 32714 4476
rect 32748 4442 32781 4476
rect 32699 4424 32781 4442
rect 33270 4435 34215 4448
rect 16881 4404 17582 4412
rect 33270 4418 33486 4435
rect 33270 4384 33339 4418
rect 33373 4384 33486 4418
rect 33538 4414 33646 4435
rect 33698 4420 33779 4435
rect 33270 4383 33486 4384
rect 33539 4383 33646 4414
rect 33707 4386 33779 4420
rect 33698 4383 33779 4386
rect 33831 4418 33892 4435
rect 33831 4384 33840 4418
rect 33874 4384 33892 4418
rect 33831 4383 33892 4384
rect 33944 4420 34215 4435
rect 33944 4419 34174 4420
rect 33944 4385 34010 4419
rect 34044 4386 34174 4419
rect 34208 4386 34215 4420
rect 34044 4385 34215 4386
rect 33944 4383 34215 4385
rect 33270 4380 33505 4383
rect 33539 4380 34215 4383
rect 33270 4365 34215 4380
rect 39672 4411 55107 4427
rect 39672 4409 46309 4411
rect 39672 4408 45973 4409
rect 39672 4407 39854 4408
rect 39672 4355 39751 4407
rect 39803 4356 39854 4407
rect 39906 4402 45973 4408
rect 39906 4368 45805 4402
rect 45839 4375 45973 4402
rect 46007 4399 46309 4409
rect 46007 4375 46141 4399
rect 45839 4368 46141 4375
rect 39906 4365 46141 4368
rect 46175 4377 46309 4399
rect 46343 4409 46641 4411
rect 46343 4377 46475 4409
rect 46175 4375 46475 4377
rect 46509 4377 46641 4409
rect 46675 4377 46809 4411
rect 46843 4409 48071 4411
rect 46843 4377 46983 4409
rect 46509 4375 46983 4377
rect 47017 4407 48071 4409
rect 47017 4403 47901 4407
rect 47017 4375 47739 4403
rect 46175 4369 47739 4375
rect 47773 4373 47901 4403
rect 47935 4377 48071 4407
rect 48105 4408 55107 4411
rect 48105 4407 54955 4408
rect 48105 4377 48235 4407
rect 47935 4373 48235 4377
rect 48269 4373 48405 4407
rect 48439 4403 48741 4407
rect 48439 4373 48573 4403
rect 47773 4369 48573 4373
rect 48607 4373 48741 4403
rect 48775 4403 54955 4407
rect 48775 4373 48915 4403
rect 48607 4369 48915 4373
rect 48949 4369 54864 4403
rect 46175 4365 54864 4369
rect 39906 4356 54864 4365
rect 39803 4355 54864 4356
rect 39672 4351 54864 4355
rect 54916 4356 54955 4403
rect 55007 4356 55107 4408
rect 54916 4351 55107 4356
rect 39672 4346 55107 4351
rect 32778 4294 32881 4313
rect 32778 4291 32868 4294
rect 9515 4252 24881 4267
rect 9515 4200 9556 4252
rect 9608 4200 9652 4252
rect 9704 4251 24881 4252
rect 9704 4249 16167 4251
rect 9704 4242 15831 4249
rect 9704 4208 15663 4242
rect 15697 4215 15831 4242
rect 15865 4239 16167 4249
rect 15865 4215 15999 4239
rect 15697 4208 15999 4215
rect 9704 4205 15999 4208
rect 16033 4217 16167 4239
rect 16201 4249 16499 4251
rect 16201 4217 16333 4249
rect 16033 4215 16333 4217
rect 16367 4217 16499 4249
rect 16533 4217 16667 4251
rect 16701 4249 17929 4251
rect 16701 4217 16841 4249
rect 16367 4215 16841 4217
rect 16875 4247 17929 4249
rect 16875 4243 17759 4247
rect 16875 4215 17597 4243
rect 16033 4209 17597 4215
rect 17631 4213 17759 4243
rect 17793 4217 17929 4247
rect 17963 4250 24881 4251
rect 17963 4247 24766 4250
rect 17963 4217 18093 4247
rect 17793 4213 18093 4217
rect 18127 4213 18263 4247
rect 18297 4243 18599 4247
rect 18297 4213 18431 4243
rect 17631 4209 18431 4213
rect 18465 4213 18599 4243
rect 18633 4243 24766 4247
rect 18633 4213 18773 4243
rect 18465 4209 18773 4213
rect 18807 4209 24667 4243
rect 16033 4205 24667 4209
rect 9704 4200 24667 4205
rect 9515 4191 24667 4200
rect 24719 4198 24766 4243
rect 24818 4198 24881 4250
rect 32809 4242 32868 4291
rect 32809 4239 32881 4242
rect 32778 4217 32881 4239
rect 34318 4217 34353 4313
rect 45973 4306 48576 4312
rect 45973 4272 46005 4306
rect 46039 4272 46105 4306
rect 46139 4272 46205 4306
rect 46239 4272 46305 4306
rect 46339 4272 46405 4306
rect 46439 4272 46505 4306
rect 46539 4272 46605 4306
rect 46639 4272 46705 4306
rect 46739 4272 47665 4306
rect 47699 4272 47765 4306
rect 47799 4272 47865 4306
rect 47899 4272 47965 4306
rect 47999 4272 48065 4306
rect 48099 4272 48165 4306
rect 48199 4272 48265 4306
rect 48299 4272 48365 4306
rect 48399 4272 48576 4306
rect 45973 4267 48576 4272
rect 45973 4264 47419 4267
rect 47269 4263 47419 4264
rect 24719 4191 24881 4198
rect 9515 4186 24881 4191
rect 47269 4211 47314 4263
rect 47366 4215 47419 4263
rect 47471 4264 48576 4267
rect 47471 4215 47497 4264
rect 47366 4211 47497 4215
rect 47269 4172 47497 4211
rect 15831 4146 18434 4152
rect 15831 4112 15863 4146
rect 15897 4112 15963 4146
rect 15997 4112 16063 4146
rect 16097 4112 16163 4146
rect 16197 4112 16263 4146
rect 16297 4112 16363 4146
rect 16397 4112 16463 4146
rect 16497 4112 16563 4146
rect 16597 4112 17523 4146
rect 17557 4112 17623 4146
rect 17657 4112 17723 4146
rect 17757 4112 17823 4146
rect 17857 4112 17923 4146
rect 17957 4112 18023 4146
rect 18057 4112 18123 4146
rect 18157 4112 18223 4146
rect 18257 4112 18434 4146
rect 15831 4107 18434 4112
rect 15831 4104 17277 4107
rect 17127 4103 17277 4104
rect 17127 4051 17172 4103
rect 17224 4055 17277 4103
rect 17329 4104 18434 4107
rect 17329 4055 17355 4104
rect 17224 4051 17355 4055
rect 17127 4012 17355 4051
rect 47023 4020 47775 4078
rect 15493 3842 15544 3938
rect 16881 3866 17562 3924
rect 22012 3869 47523 3913
rect 22012 3867 47411 3869
rect 15493 3841 15543 3842
rect 22012 3815 33475 3867
rect 33527 3815 33619 3867
rect 33671 3815 33763 3867
rect 33815 3866 47411 3867
rect 33815 3815 47322 3866
rect 22012 3814 47322 3815
rect 47374 3817 47411 3866
rect 47463 3817 47523 3869
rect 47374 3814 47523 3817
rect 22012 3790 47523 3814
rect 22012 3783 47322 3790
rect 22012 3731 33474 3783
rect 33526 3731 33618 3783
rect 33670 3731 33762 3783
rect 33814 3738 47322 3783
rect 47374 3738 47415 3790
rect 47467 3738 47523 3790
rect 33814 3731 47523 3738
rect 17139 3707 47523 3731
rect 17139 3686 22218 3707
rect 17139 3634 17176 3686
rect 17228 3681 22218 3686
rect 17228 3634 17270 3681
rect 17139 3629 17270 3634
rect 17322 3629 22218 3681
rect 17139 3608 22218 3629
rect 17139 3606 17270 3608
rect 9306 3532 9969 3590
rect 17139 3554 17176 3606
rect 17228 3556 17270 3606
rect 17322 3556 22218 3608
rect 17228 3554 22218 3556
rect 17139 3525 22218 3554
rect 24404 3544 25032 3602
rect 39416 3544 40179 3602
rect 54606 3535 55257 3593
rect 62673 1474 62895 1552
<< via1 >>
rect 9555 5455 9607 5507
rect 9636 5454 9688 5506
rect 24671 5452 24723 5504
rect 24766 5452 24818 5504
rect 16734 5389 16786 5441
rect 16812 5389 16864 5441
rect 16905 5389 16957 5441
rect 32693 5412 32745 5464
rect 32806 5412 32858 5464
rect 32907 5412 32959 5464
rect 39748 5454 39800 5506
rect 39850 5454 39902 5506
rect 46885 5389 46937 5441
rect 46968 5389 47020 5441
rect 54866 5427 54918 5479
rect 54961 5427 55013 5479
rect 8563 5233 8615 5285
rect 8670 5235 8722 5287
rect 8772 5235 8824 5287
rect 8872 5236 8924 5288
rect 23593 5239 23645 5291
rect 23696 5239 23748 5291
rect 23779 5239 23831 5291
rect 23880 5239 23932 5291
rect 23967 5239 24019 5291
rect 38725 5235 38777 5287
rect 38813 5235 38865 5287
rect 38898 5240 38950 5292
rect 55641 5232 55693 5284
rect 55735 5232 55787 5284
rect 55812 5232 55864 5284
rect 55892 5231 55944 5283
rect 55966 5232 56018 5284
rect 32705 4789 32757 4841
rect 32808 4792 32860 4844
rect 32909 4792 32961 4844
rect 46891 4564 46943 4616
rect 46981 4565 47033 4617
rect 16758 4412 16810 4464
rect 16881 4412 16933 4464
rect 33486 4414 33538 4435
rect 33646 4420 33698 4435
rect 33486 4383 33505 4414
rect 33505 4383 33538 4414
rect 33646 4386 33673 4420
rect 33673 4386 33698 4420
rect 33646 4383 33698 4386
rect 33779 4383 33831 4435
rect 33892 4383 33944 4435
rect 39751 4355 39803 4407
rect 39854 4356 39906 4408
rect 54864 4351 54916 4403
rect 54955 4356 55007 4408
rect 9556 4200 9608 4252
rect 9652 4200 9704 4252
rect 24667 4191 24719 4243
rect 24766 4198 24818 4250
rect 32661 4237 32713 4289
rect 32757 4239 32809 4291
rect 32868 4242 32920 4294
rect 32960 4239 33012 4291
rect 47314 4211 47366 4263
rect 47419 4215 47471 4267
rect 17172 4051 17224 4103
rect 17277 4055 17329 4107
rect 48326 4024 48378 4076
rect 48418 4025 48470 4077
rect 48508 4024 48560 4076
rect 48596 4023 48648 4075
rect 15971 3863 16023 3915
rect 16055 3863 16107 3915
rect 16148 3864 16200 3916
rect 33475 3815 33527 3867
rect 33619 3815 33671 3867
rect 33763 3815 33815 3867
rect 47322 3814 47374 3866
rect 47411 3817 47463 3869
rect 33474 3731 33526 3783
rect 33618 3731 33670 3783
rect 33762 3731 33814 3783
rect 47322 3738 47374 3790
rect 47415 3738 47467 3790
rect 17176 3634 17228 3686
rect 17270 3629 17322 3681
rect 8557 3535 8609 3587
rect 8655 3535 8707 3587
rect 8750 3535 8802 3587
rect 8855 3535 8907 3587
rect 17176 3554 17228 3606
rect 17270 3556 17322 3608
rect 23607 3540 23659 3592
rect 23707 3540 23759 3592
rect 23806 3540 23858 3592
rect 23909 3540 23961 3592
rect 38715 3534 38767 3586
rect 38803 3534 38855 3586
rect 38901 3530 38953 3582
rect 55637 3531 55689 3583
rect 55725 3531 55777 3583
rect 55808 3531 55860 3583
rect 55895 3531 55947 3583
rect 9556 3317 9608 3369
rect 9636 3315 9688 3367
rect 24672 3332 24724 3384
rect 24755 3332 24807 3384
rect 39750 3322 39802 3374
rect 39841 3322 39893 3374
rect 54867 3307 54919 3359
rect 54950 3307 55002 3359
<< metal2 >>
rect 5569 7342 5613 8498
rect 7457 7342 7501 8498
rect 9345 7342 9389 8498
rect 11233 7342 11277 8498
rect 13121 7342 13165 8498
rect 15009 7342 15053 8498
rect 16897 7342 16941 8498
rect 18785 7342 18829 8498
rect 20673 7342 20717 8498
rect 22561 7342 22605 8498
rect 24449 7342 24493 8498
rect 26337 7342 26381 8498
rect 28225 7342 28269 8498
rect 30113 7342 30157 8498
rect 32001 7342 32045 8498
rect 33889 7342 33933 8498
rect 35777 7342 35821 8498
rect 37665 7342 37709 8498
rect 39553 7342 39597 8498
rect 41441 7342 41485 8498
rect 43329 7342 43373 8498
rect 45217 7342 45261 8498
rect 47105 7342 47149 8498
rect 48993 7342 49037 8498
rect 50881 7342 50925 8498
rect 52769 7342 52813 8498
rect 54657 7342 54701 8498
rect 56545 7342 56589 8498
rect 58433 7342 58477 8498
rect 60321 7342 60365 8498
rect 62209 7342 62253 8498
rect 208 6660 322 6695
rect 64230 6660 64344 6699
rect 208 6624 4285 6660
rect 62229 6624 64344 6660
rect 208 2204 322 6624
rect 9531 5507 9720 5537
rect 9531 5455 9555 5507
rect 9607 5506 9720 5507
rect 9607 5455 9636 5506
rect 9531 5454 9636 5455
rect 9688 5454 9720 5506
rect 8499 5288 8983 5413
rect 8499 5287 8872 5288
rect 8499 5285 8670 5287
rect 8499 5233 8563 5285
rect 8615 5235 8670 5285
rect 8722 5235 8772 5287
rect 8824 5236 8872 5287
rect 8924 5236 8983 5288
rect 8824 5235 8983 5236
rect 8615 5233 8983 5235
rect 8499 4066 8983 5233
rect 8499 4010 8566 4066
rect 8622 4010 8680 4066
rect 8736 4010 8794 4066
rect 8850 4010 8983 4066
rect 8499 3951 8983 4010
rect 8499 3895 8566 3951
rect 8622 3895 8680 3951
rect 8736 3895 8794 3951
rect 8850 3895 8983 3951
rect 8499 3836 8983 3895
rect 8499 3780 8566 3836
rect 8622 3780 8680 3836
rect 8736 3780 8794 3836
rect 8850 3780 8983 3836
rect 8499 3587 8983 3780
rect 8499 3535 8557 3587
rect 8609 3535 8655 3587
rect 8707 3535 8750 3587
rect 8802 3535 8855 3587
rect 8907 3535 8983 3587
rect 8499 3423 8983 3535
rect 9531 4252 9720 5454
rect 16714 5441 16974 5512
rect 16714 5389 16734 5441
rect 16786 5389 16812 5441
rect 16864 5389 16905 5441
rect 16957 5389 16974 5441
rect 24642 5504 24831 5527
rect 24642 5452 24671 5504
rect 24723 5452 24766 5504
rect 24818 5452 24831 5504
rect 16714 4464 16974 5389
rect 16714 4412 16758 4464
rect 16810 4412 16881 4464
rect 16933 4412 16974 4464
rect 16714 4368 16974 4412
rect 23555 5291 24022 5391
rect 23555 5239 23593 5291
rect 23645 5239 23696 5291
rect 23748 5239 23779 5291
rect 23831 5239 23880 5291
rect 23932 5239 23967 5291
rect 24019 5239 24022 5291
rect 9531 4200 9556 4252
rect 9608 4200 9652 4252
rect 9704 4200 9720 4252
rect 9531 3369 9720 4200
rect 17139 4107 17345 4152
rect 17139 4103 17277 4107
rect 17139 4051 17172 4103
rect 17224 4055 17277 4103
rect 17329 4055 17345 4107
rect 17224 4051 17345 4055
rect 9531 3317 9556 3369
rect 9608 3367 9720 3369
rect 9608 3317 9636 3367
rect 9531 3315 9636 3317
rect 9688 3315 9720 3367
rect 15920 3916 16273 3962
rect 15920 3915 16148 3916
rect 15920 3863 15971 3915
rect 16023 3863 16055 3915
rect 16107 3864 16148 3915
rect 16200 3864 16273 3916
rect 16107 3863 16273 3864
rect 15920 3505 16273 3863
rect 17139 3686 17345 4051
rect 17139 3634 17176 3686
rect 17228 3681 17345 3686
rect 17228 3634 17270 3681
rect 17139 3629 17270 3634
rect 17322 3629 17345 3681
rect 17139 3608 17345 3629
rect 17139 3606 17270 3608
rect 17139 3554 17176 3606
rect 17228 3556 17270 3606
rect 17322 3556 17345 3608
rect 17228 3554 17345 3556
rect 17139 3525 17345 3554
rect 23555 3976 24022 5239
rect 23555 3920 23605 3976
rect 23661 3920 23709 3976
rect 23765 3920 23813 3976
rect 23869 3920 23917 3976
rect 23973 3920 24022 3976
rect 23555 3860 24022 3920
rect 23555 3804 23605 3860
rect 23661 3804 23709 3860
rect 23765 3804 23813 3860
rect 23869 3804 23917 3860
rect 23973 3804 24022 3860
rect 23555 3744 24022 3804
rect 23555 3688 23605 3744
rect 23661 3688 23709 3744
rect 23765 3688 23813 3744
rect 23869 3688 23917 3744
rect 23973 3688 24022 3744
rect 23555 3592 24022 3688
rect 23555 3540 23607 3592
rect 23659 3540 23707 3592
rect 23759 3540 23806 3592
rect 23858 3540 23909 3592
rect 23961 3540 24022 3592
rect 15920 3449 15960 3505
rect 16016 3449 16068 3505
rect 16124 3449 16176 3505
rect 16232 3449 16273 3505
rect 15920 3411 16273 3449
rect 23555 3440 24022 3540
rect 24642 4250 24831 5452
rect 32647 5464 32982 5507
rect 32647 5412 32693 5464
rect 32745 5412 32806 5464
rect 32858 5412 32907 5464
rect 32959 5412 32982 5464
rect 32647 4844 32982 5412
rect 39733 5506 39920 5525
rect 39733 5454 39748 5506
rect 39800 5454 39850 5506
rect 39902 5454 39920 5506
rect 32647 4841 32808 4844
rect 32647 4789 32705 4841
rect 32757 4792 32808 4841
rect 32860 4792 32909 4844
rect 32961 4792 32982 4844
rect 32757 4789 32982 4792
rect 32647 4757 32982 4789
rect 38671 5292 38971 5389
rect 38671 5287 38898 5292
rect 38671 5235 38725 5287
rect 38777 5235 38813 5287
rect 38865 5240 38898 5287
rect 38950 5240 38971 5292
rect 38865 5235 38971 5240
rect 33418 4435 33957 4458
rect 33418 4383 33486 4435
rect 33538 4383 33646 4435
rect 33698 4383 33779 4435
rect 33831 4383 33892 4435
rect 33944 4383 33957 4435
rect 24642 4243 24766 4250
rect 24642 4191 24667 4243
rect 24719 4198 24766 4243
rect 24818 4198 24831 4250
rect 24719 4191 24831 4198
rect 15920 3355 15960 3411
rect 16016 3355 16068 3411
rect 16124 3355 16176 3411
rect 16232 3355 16273 3411
rect 15920 3329 16273 3355
rect 24642 3384 24831 4191
rect 32609 4294 33034 4312
rect 32609 4291 32868 4294
rect 32609 4289 32757 4291
rect 32609 4237 32661 4289
rect 32713 4239 32757 4289
rect 32809 4242 32868 4291
rect 32920 4291 33034 4294
rect 32920 4242 32960 4291
rect 32809 4239 32960 4242
rect 33012 4239 33034 4291
rect 32713 4237 33034 4239
rect 32609 3625 33034 4237
rect 33418 3867 33957 4383
rect 33418 3815 33475 3867
rect 33527 3815 33619 3867
rect 33671 3815 33763 3867
rect 33815 3815 33957 3867
rect 33418 3783 33957 3815
rect 33418 3731 33474 3783
rect 33526 3731 33618 3783
rect 33670 3731 33762 3783
rect 33814 3731 33957 3783
rect 33418 3657 33957 3731
rect 38671 4325 38971 5235
rect 38671 4269 38692 4325
rect 38748 4269 38786 4325
rect 38842 4269 38880 4325
rect 38936 4269 38971 4325
rect 38671 4237 38971 4269
rect 38671 4181 38692 4237
rect 38748 4181 38786 4237
rect 38842 4181 38880 4237
rect 38936 4181 38971 4237
rect 38671 4149 38971 4181
rect 38671 4093 38692 4149
rect 38748 4093 38786 4149
rect 38842 4093 38880 4149
rect 38936 4093 38971 4149
rect 32609 3569 32655 3625
rect 32711 3569 32780 3625
rect 32836 3569 32905 3625
rect 32961 3569 33034 3625
rect 32609 3529 33034 3569
rect 32609 3473 32655 3529
rect 32711 3473 32780 3529
rect 32836 3473 32905 3529
rect 32961 3473 33034 3529
rect 32609 3441 33034 3473
rect 38671 3586 38971 4093
rect 38671 3534 38715 3586
rect 38767 3534 38803 3586
rect 38855 3582 38971 3586
rect 38855 3534 38901 3582
rect 38671 3530 38901 3534
rect 38953 3530 38971 3582
rect 38671 3437 38971 3530
rect 39733 4408 39920 5454
rect 46862 5441 47081 5494
rect 46862 5389 46885 5441
rect 46937 5389 46968 5441
rect 47020 5389 47081 5441
rect 46862 4617 47081 5389
rect 46862 4616 46981 4617
rect 46862 4564 46891 4616
rect 46943 4565 46981 4616
rect 47033 4565 47081 4617
rect 46943 4564 47081 4565
rect 46862 4529 47081 4564
rect 54837 5479 55026 5502
rect 54837 5427 54866 5479
rect 54918 5427 54961 5479
rect 55013 5427 55026 5479
rect 39733 4407 39854 4408
rect 39733 4355 39751 4407
rect 39803 4356 39854 4407
rect 39906 4356 39920 4408
rect 39803 4355 39920 4356
rect 24642 3332 24672 3384
rect 24724 3332 24755 3384
rect 24807 3332 24831 3384
rect 24642 3319 24831 3332
rect 39733 3374 39920 4355
rect 54837 4408 55026 5427
rect 54837 4403 54955 4408
rect 54837 4351 54864 4403
rect 54916 4356 54955 4403
rect 55007 4356 55026 4408
rect 54916 4351 55026 4356
rect 47281 4267 47487 4312
rect 47281 4263 47419 4267
rect 47281 4211 47314 4263
rect 47366 4215 47419 4263
rect 47471 4215 47487 4267
rect 47366 4211 47487 4215
rect 47281 3869 47487 4211
rect 47281 3866 47411 3869
rect 47281 3814 47322 3866
rect 47374 3817 47411 3866
rect 47463 3817 47487 3869
rect 47374 3814 47487 3817
rect 47281 3790 47487 3814
rect 47281 3738 47322 3790
rect 47374 3738 47415 3790
rect 47467 3738 47487 3790
rect 47281 3695 47487 3738
rect 48289 4077 48703 4099
rect 48289 4076 48418 4077
rect 48289 4024 48326 4076
rect 48378 4025 48418 4076
rect 48470 4076 48703 4077
rect 48470 4025 48508 4076
rect 48378 4024 48508 4025
rect 48560 4075 48703 4076
rect 48560 4024 48596 4075
rect 48289 4023 48596 4024
rect 48648 4023 48703 4075
rect 39733 3322 39750 3374
rect 39802 3322 39841 3374
rect 39893 3322 39920 3374
rect 9531 3297 9720 3315
rect 39733 3314 39920 3322
rect 48289 3478 48703 4023
rect 48289 3422 48326 3478
rect 48382 3422 48419 3478
rect 48475 3422 48512 3478
rect 48568 3422 48605 3478
rect 48661 3422 48703 3478
rect 48289 3396 48703 3422
rect 48289 3340 48326 3396
rect 48382 3340 48419 3396
rect 48475 3340 48512 3396
rect 48568 3340 48605 3396
rect 48661 3340 48703 3396
rect 48289 3303 48703 3340
rect 54837 3359 55026 4351
rect 55602 5284 56023 5389
rect 55602 5232 55641 5284
rect 55693 5232 55735 5284
rect 55787 5232 55812 5284
rect 55864 5283 55966 5284
rect 55864 5232 55892 5283
rect 55602 5231 55892 5232
rect 55944 5232 55966 5283
rect 56018 5232 56023 5284
rect 55944 5231 56023 5232
rect 55602 3870 56023 5231
rect 55602 3814 55639 3870
rect 55695 3814 55743 3870
rect 55799 3814 55847 3870
rect 55903 3814 55951 3870
rect 56007 3814 56023 3870
rect 55602 3780 56023 3814
rect 55602 3724 55639 3780
rect 55695 3724 55743 3780
rect 55799 3724 55847 3780
rect 55903 3724 55951 3780
rect 56007 3724 56023 3780
rect 55602 3583 56023 3724
rect 55602 3531 55637 3583
rect 55689 3531 55725 3583
rect 55777 3531 55808 3583
rect 55860 3531 55895 3583
rect 55947 3531 56023 3583
rect 55602 3439 56023 3531
rect 54837 3307 54867 3359
rect 54919 3307 54950 3359
rect 55002 3307 55026 3359
rect 54837 3294 55026 3307
rect 932 3058 2360 3248
rect 932 2804 1818 3058
rect 932 2718 2340 2804
rect 932 2710 1818 2718
rect 64230 2204 64344 6624
rect 208 2168 603 2204
rect 1752 2168 2342 2204
rect 62578 2168 64344 2204
rect 208 2156 322 2168
rect 64230 2160 64344 2168
rect 2311 1168 2355 1486
rect 4199 1168 4243 1486
rect 6087 1168 6131 1486
rect 7975 1168 8019 1486
rect 9863 1168 9907 1486
rect 11751 1168 11795 1486
rect 13639 1168 13683 1486
rect 15527 1168 15571 1486
rect 17415 1168 17459 1486
rect 19303 1168 19347 1486
rect 21191 1168 21235 1486
rect 23079 1168 23123 1486
rect 24967 1168 25011 1486
rect 26855 1168 26899 1486
rect 28743 1168 28787 1486
rect 30631 1168 30675 1486
rect 32519 1168 32563 1486
rect 34407 1168 34451 1486
rect 36295 1168 36339 1486
rect 38183 1168 38227 1486
rect 40071 1168 40115 1486
rect 41959 1168 42003 1486
rect 43847 1168 43891 1486
rect 45735 1168 45779 1486
rect 47623 1168 47667 1486
rect 49511 1168 49555 1486
rect 51399 1168 51443 1486
rect 53287 1168 53331 1486
rect 55175 1168 55219 1486
rect 57063 1168 57107 1486
rect 58951 1366 58995 1486
rect 58951 1168 58997 1366
rect 422 22 467 1168
rect 2310 22 2355 1168
rect 4198 22 4243 1168
rect 6086 22 6131 1168
rect 7974 22 8019 1168
rect 9862 22 9907 1168
rect 11750 22 11795 1168
rect 13638 22 13683 1168
rect 15526 22 15571 1168
rect 17414 22 17459 1168
rect 19302 22 19347 1168
rect 21190 22 21235 1168
rect 23078 22 23123 1168
rect 24966 22 25011 1168
rect 26854 22 26899 1168
rect 28742 22 28787 1168
rect 30630 22 30675 1168
rect 32518 22 32563 1168
rect 34406 22 34451 1168
rect 36294 22 36339 1168
rect 38182 22 38227 1168
rect 40070 22 40115 1168
rect 41958 22 42003 1168
rect 43846 22 43891 1168
rect 45734 22 45779 1168
rect 47622 22 47667 1168
rect 49510 22 49555 1168
rect 51398 22 51443 1168
rect 53286 22 53331 1168
rect 55174 22 55219 1168
rect 57062 22 57107 1168
rect 58950 468 58997 1168
rect 58950 22 58995 468
rect 60827 0 60883 1486
<< via2 >>
rect 8566 4010 8622 4066
rect 8680 4010 8736 4066
rect 8794 4010 8850 4066
rect 8566 3895 8622 3951
rect 8680 3895 8736 3951
rect 8794 3895 8850 3951
rect 8566 3780 8622 3836
rect 8680 3780 8736 3836
rect 8794 3780 8850 3836
rect 23605 3920 23661 3976
rect 23709 3920 23765 3976
rect 23813 3920 23869 3976
rect 23917 3920 23973 3976
rect 23605 3804 23661 3860
rect 23709 3804 23765 3860
rect 23813 3804 23869 3860
rect 23917 3804 23973 3860
rect 23605 3688 23661 3744
rect 23709 3688 23765 3744
rect 23813 3688 23869 3744
rect 23917 3688 23973 3744
rect 15960 3449 16016 3505
rect 16068 3449 16124 3505
rect 16176 3449 16232 3505
rect 15960 3355 16016 3411
rect 16068 3355 16124 3411
rect 16176 3355 16232 3411
rect 38692 4269 38748 4325
rect 38786 4269 38842 4325
rect 38880 4269 38936 4325
rect 38692 4181 38748 4237
rect 38786 4181 38842 4237
rect 38880 4181 38936 4237
rect 38692 4093 38748 4149
rect 38786 4093 38842 4149
rect 38880 4093 38936 4149
rect 32655 3569 32711 3625
rect 32780 3569 32836 3625
rect 32905 3569 32961 3625
rect 32655 3473 32711 3529
rect 32780 3473 32836 3529
rect 32905 3473 32961 3529
rect 48326 3422 48382 3478
rect 48419 3422 48475 3478
rect 48512 3422 48568 3478
rect 48605 3422 48661 3478
rect 48326 3340 48382 3396
rect 48419 3340 48475 3396
rect 48512 3340 48568 3396
rect 48605 3340 48661 3396
rect 55639 3814 55695 3870
rect 55743 3814 55799 3870
rect 55847 3814 55903 3870
rect 55951 3814 56007 3870
rect 55639 3724 55695 3780
rect 55743 3724 55799 3780
rect 55847 3724 55903 3780
rect 55951 3724 56007 3780
<< metal3 >>
rect 4809 8066 4915 8083
rect 4809 8002 4830 8066
rect 4894 8002 4915 8066
rect 4809 7986 4915 8002
rect 4809 7922 4830 7986
rect 4894 7922 4915 7986
rect 4809 7905 4915 7922
rect 5018 8065 5124 8082
rect 5018 8001 5039 8065
rect 5103 8001 5124 8065
rect 5018 7985 5124 8001
rect 5018 7921 5039 7985
rect 5103 7921 5124 7985
rect 5018 7904 5124 7921
rect 5184 8065 5290 8082
rect 5184 8001 5205 8065
rect 5269 8001 5290 8065
rect 5184 7985 5290 8001
rect 5184 7921 5205 7985
rect 5269 7921 5290 7985
rect 5184 7904 5290 7921
rect 5364 8067 5470 8084
rect 5364 8003 5385 8067
rect 5449 8003 5470 8067
rect 5364 7987 5470 8003
rect 5364 7923 5385 7987
rect 5449 7923 5470 7987
rect 5364 7906 5470 7923
rect 21438 8083 21544 8100
rect 21438 8019 21459 8083
rect 21523 8019 21544 8083
rect 21438 8003 21544 8019
rect 21438 7939 21459 8003
rect 21523 7939 21544 8003
rect 21438 7922 21544 7939
rect 21654 8083 21760 8100
rect 21654 8019 21675 8083
rect 21739 8019 21760 8083
rect 21654 8003 21760 8019
rect 21654 7939 21675 8003
rect 21739 7939 21760 8003
rect 21654 7922 21760 7939
rect 21870 8083 21976 8100
rect 21870 8019 21891 8083
rect 21955 8019 21976 8083
rect 21870 8003 21976 8019
rect 21870 7939 21891 8003
rect 21955 7939 21976 8003
rect 21870 7922 21976 7939
rect 29930 8082 30036 8099
rect 29930 8018 29951 8082
rect 30015 8018 30036 8082
rect 29930 8002 30036 8018
rect 29930 7938 29951 8002
rect 30015 7938 30036 8002
rect 29930 7921 30036 7938
rect 30146 8082 30252 8099
rect 30146 8018 30167 8082
rect 30231 8018 30252 8082
rect 30146 8002 30252 8018
rect 30146 7938 30167 8002
rect 30231 7938 30252 8002
rect 30146 7921 30252 7938
rect 30362 8082 30468 8099
rect 30362 8018 30383 8082
rect 30447 8018 30468 8082
rect 30362 8002 30468 8018
rect 30362 7938 30383 8002
rect 30447 7938 30468 8002
rect 30362 7921 30468 7938
rect 43458 8088 43564 8105
rect 43458 8024 43479 8088
rect 43543 8024 43564 8088
rect 43458 8008 43564 8024
rect 43458 7944 43479 8008
rect 43543 7944 43564 8008
rect 43458 7927 43564 7944
rect 43674 8088 43780 8105
rect 43674 8024 43695 8088
rect 43759 8024 43780 8088
rect 43674 8008 43780 8024
rect 43674 7944 43695 8008
rect 43759 7944 43780 8008
rect 43674 7927 43780 7944
rect 43890 8088 43996 8105
rect 43890 8024 43911 8088
rect 43975 8024 43996 8088
rect 43890 8008 43996 8024
rect 43890 7944 43911 8008
rect 43975 7944 43996 8008
rect 43890 7927 43996 7944
rect 59943 8081 60049 8098
rect 59943 8017 59964 8081
rect 60028 8017 60049 8081
rect 59943 8001 60049 8017
rect 59943 7937 59964 8001
rect 60028 7937 60049 8001
rect 59943 7920 60049 7937
rect 60159 8081 60265 8098
rect 60159 8017 60180 8081
rect 60244 8017 60265 8081
rect 60159 8001 60265 8017
rect 60159 7937 60180 8001
rect 60244 7937 60265 8001
rect 60159 7920 60265 7937
rect 60375 8081 60481 8098
rect 60375 8017 60396 8081
rect 60460 8017 60481 8081
rect 60375 8001 60481 8017
rect 60375 7937 60396 8001
rect 60460 7937 60481 8001
rect 60375 7920 60481 7937
rect 3463 5949 4358 6012
rect 3463 5948 3768 5949
rect 3463 5884 3596 5948
rect 3660 5885 3768 5948
rect 3832 5948 4358 5949
rect 3832 5885 3942 5948
rect 3660 5884 3942 5885
rect 4006 5884 4358 5948
rect 3463 5869 4358 5884
rect 3463 5868 3768 5869
rect 3463 5804 3596 5868
rect 3660 5805 3768 5868
rect 3832 5868 4358 5869
rect 3832 5805 3942 5868
rect 3660 5804 3942 5805
rect 4006 5804 4358 5868
rect 19903 5969 20009 5986
rect 19903 5905 19924 5969
rect 19988 5905 20009 5969
rect 19903 5889 20009 5905
rect 19903 5825 19924 5889
rect 19988 5825 20009 5889
rect 19903 5808 20009 5825
rect 20119 5969 20225 5986
rect 20119 5905 20140 5969
rect 20204 5905 20225 5969
rect 20119 5889 20225 5905
rect 20119 5825 20140 5889
rect 20204 5825 20225 5889
rect 20119 5808 20225 5825
rect 20335 5969 20441 5986
rect 20335 5905 20356 5969
rect 20420 5905 20441 5969
rect 20335 5889 20441 5905
rect 20335 5825 20356 5889
rect 20420 5825 20441 5889
rect 20335 5808 20441 5825
rect 28411 5961 28517 5978
rect 28411 5897 28432 5961
rect 28496 5897 28517 5961
rect 28411 5881 28517 5897
rect 28411 5817 28432 5881
rect 28496 5817 28517 5881
rect 3463 5758 4358 5804
rect 28411 5800 28517 5817
rect 28627 5961 28733 5978
rect 28627 5897 28648 5961
rect 28712 5897 28733 5961
rect 28627 5881 28733 5897
rect 28627 5817 28648 5881
rect 28712 5817 28733 5881
rect 28627 5800 28733 5817
rect 28843 5961 28949 5978
rect 28843 5897 28864 5961
rect 28928 5897 28949 5961
rect 28843 5881 28949 5897
rect 28843 5817 28864 5881
rect 28928 5817 28949 5881
rect 28843 5800 28949 5817
rect 41883 5956 41989 5973
rect 41883 5892 41904 5956
rect 41968 5892 41989 5956
rect 41883 5876 41989 5892
rect 41883 5812 41904 5876
rect 41968 5812 41989 5876
rect 41883 5795 41989 5812
rect 42099 5956 42205 5973
rect 42099 5892 42120 5956
rect 42184 5892 42205 5956
rect 42099 5876 42205 5892
rect 42099 5812 42120 5876
rect 42184 5812 42205 5876
rect 42099 5795 42205 5812
rect 42315 5956 42421 5973
rect 42315 5892 42336 5956
rect 42400 5892 42421 5956
rect 42315 5876 42421 5892
rect 42315 5812 42336 5876
rect 42400 5812 42421 5876
rect 42315 5795 42421 5812
rect 58434 5948 58540 5965
rect 58434 5884 58455 5948
rect 58519 5884 58540 5948
rect 58434 5868 58540 5884
rect 58434 5804 58455 5868
rect 58519 5804 58540 5868
rect 58434 5787 58540 5804
rect 58650 5948 58756 5965
rect 58650 5884 58671 5948
rect 58735 5884 58756 5948
rect 58650 5868 58756 5884
rect 58650 5804 58671 5868
rect 58735 5804 58756 5868
rect 58650 5787 58756 5804
rect 58866 5948 58972 5965
rect 58866 5884 58887 5948
rect 58951 5884 58972 5948
rect 58866 5868 58972 5884
rect 58866 5804 58887 5868
rect 58951 5804 58972 5868
rect 58866 5787 58972 5804
rect 38669 4325 38973 4339
rect 38669 4269 38692 4325
rect 38748 4269 38786 4325
rect 38842 4269 38880 4325
rect 38936 4269 38973 4325
rect 38669 4237 38973 4269
rect 38669 4181 38692 4237
rect 38748 4202 38786 4237
rect 38780 4181 38786 4202
rect 38842 4203 38880 4237
rect 38842 4181 38870 4203
rect 38936 4181 38973 4237
rect 38669 4149 38716 4181
rect 38780 4149 38870 4181
rect 38934 4149 38973 4181
rect 8565 4092 8907 4125
rect 38669 4093 38692 4149
rect 38780 4138 38786 4149
rect 38748 4093 38786 4138
rect 38842 4139 38870 4149
rect 38842 4093 38880 4139
rect 38936 4093 38973 4149
rect 8497 4066 8986 4092
rect 38669 4073 38973 4093
rect 8497 4010 8566 4066
rect 8622 4010 8680 4066
rect 8736 4010 8794 4066
rect 8850 4010 8986 4066
rect 8497 3951 8986 4010
rect 8497 3895 8566 3951
rect 8622 3909 8680 3951
rect 8736 3915 8794 3951
rect 8638 3895 8680 3909
rect 8789 3895 8794 3915
rect 8850 3915 8986 3951
rect 8850 3895 8870 3915
rect 8497 3845 8574 3895
rect 8638 3851 8725 3895
rect 8789 3851 8870 3895
rect 8934 3851 8986 3915
rect 8638 3845 8986 3851
rect 8497 3836 8986 3845
rect 8497 3780 8566 3836
rect 8622 3780 8680 3836
rect 8736 3780 8794 3836
rect 8850 3780 8986 3836
rect 8497 3725 8986 3780
rect 23555 3976 24022 4030
rect 23555 3920 23605 3976
rect 23661 3923 23709 3976
rect 23681 3920 23709 3923
rect 23765 3923 23813 3976
rect 23765 3920 23784 3923
rect 23869 3920 23917 3976
rect 23973 3920 24022 3976
rect 23555 3860 23617 3920
rect 23681 3860 23784 3920
rect 23848 3860 24022 3920
rect 23555 3804 23605 3860
rect 23681 3859 23709 3860
rect 23661 3804 23709 3859
rect 23765 3859 23784 3860
rect 23765 3804 23813 3859
rect 23869 3804 23917 3860
rect 23973 3804 24022 3860
rect 23555 3762 24022 3804
rect 23555 3744 23617 3762
rect 23681 3744 23784 3762
rect 23848 3744 24022 3762
rect 23555 3688 23605 3744
rect 23681 3698 23709 3744
rect 23661 3688 23709 3698
rect 23765 3698 23784 3744
rect 23765 3688 23813 3698
rect 23869 3688 23917 3744
rect 23973 3688 24022 3744
rect 55602 3870 56024 3898
rect 55602 3814 55639 3870
rect 55720 3814 55743 3870
rect 55841 3814 55847 3870
rect 55903 3814 55915 3870
rect 56007 3814 56024 3870
rect 55602 3806 55656 3814
rect 55720 3806 55777 3814
rect 55841 3806 55915 3814
rect 55979 3806 56024 3814
rect 55602 3790 56024 3806
rect 55602 3780 55656 3790
rect 55720 3780 55777 3790
rect 55841 3780 55915 3790
rect 55979 3780 56024 3790
rect 55602 3724 55639 3780
rect 55720 3726 55743 3780
rect 55841 3726 55847 3780
rect 55695 3724 55743 3726
rect 55799 3724 55847 3726
rect 55903 3726 55915 3780
rect 55903 3724 55951 3726
rect 56007 3724 56024 3780
rect 55602 3690 56024 3724
rect 23555 3644 24022 3688
rect 32607 3625 33032 3663
rect 32607 3569 32655 3625
rect 32711 3569 32780 3625
rect 32836 3569 32905 3625
rect 32961 3569 33032 3625
rect 32607 3562 33032 3569
rect 32607 3529 32664 3562
rect 32728 3529 32783 3562
rect 15920 3505 16273 3528
rect 15920 3454 15960 3505
rect 16016 3454 16068 3505
rect 16124 3454 16176 3505
rect 15920 3390 15950 3454
rect 16016 3449 16053 3454
rect 16124 3449 16156 3454
rect 16232 3449 16273 3505
rect 16014 3411 16053 3449
rect 16117 3411 16156 3449
rect 16220 3411 16273 3449
rect 32607 3473 32655 3529
rect 32728 3498 32780 3529
rect 32847 3498 32902 3562
rect 32966 3498 33032 3562
rect 32711 3473 32780 3498
rect 32836 3473 32905 3498
rect 32961 3473 33032 3498
rect 32607 3436 33032 3473
rect 48289 3495 48704 3545
rect 48289 3494 48477 3495
rect 48289 3478 48337 3494
rect 48401 3478 48477 3494
rect 48541 3478 48605 3495
rect 16016 3390 16053 3411
rect 16124 3390 16156 3411
rect 15920 3355 15960 3390
rect 16016 3355 16068 3390
rect 16124 3355 16176 3390
rect 16232 3355 16273 3411
rect 15920 3329 16273 3355
rect 48289 3422 48326 3478
rect 48401 3430 48419 3478
rect 48382 3422 48419 3430
rect 48475 3431 48477 3478
rect 48475 3422 48512 3431
rect 48568 3422 48605 3478
rect 48669 3431 48704 3495
rect 48661 3422 48704 3431
rect 48289 3415 48704 3422
rect 48289 3414 48477 3415
rect 48289 3396 48337 3414
rect 48401 3396 48477 3414
rect 48541 3396 48605 3415
rect 48289 3340 48326 3396
rect 48401 3350 48419 3396
rect 48382 3340 48419 3350
rect 48475 3351 48477 3396
rect 48475 3340 48512 3351
rect 48568 3340 48605 3396
rect 48669 3351 48704 3415
rect 48661 3340 48704 3351
rect 48289 3304 48704 3340
rect 3577 3000 3683 3017
rect 3577 2936 3598 3000
rect 3662 2936 3683 3000
rect 3577 2920 3683 2936
rect 3577 2856 3598 2920
rect 3662 2856 3683 2920
rect 3577 2839 3683 2856
rect 3782 3002 3888 3019
rect 3782 2938 3803 3002
rect 3867 2938 3888 3002
rect 3782 2922 3888 2938
rect 3782 2858 3803 2922
rect 3867 2858 3888 2922
rect 3782 2841 3888 2858
rect 3981 3002 4087 3019
rect 3981 2938 4002 3002
rect 4066 2938 4087 3002
rect 3981 2922 4087 2938
rect 3981 2858 4002 2922
rect 4066 2858 4087 2922
rect 3981 2841 4087 2858
rect 19894 3018 20000 3035
rect 19894 2954 19915 3018
rect 19979 2954 20000 3018
rect 19894 2938 20000 2954
rect 19894 2874 19915 2938
rect 19979 2874 20000 2938
rect 19894 2857 20000 2874
rect 20110 3018 20216 3035
rect 20110 2954 20131 3018
rect 20195 2954 20216 3018
rect 20110 2938 20216 2954
rect 20110 2874 20131 2938
rect 20195 2874 20216 2938
rect 20110 2857 20216 2874
rect 20326 3018 20432 3035
rect 20326 2954 20347 3018
rect 20411 2954 20432 3018
rect 20326 2938 20432 2954
rect 20326 2874 20347 2938
rect 20411 2874 20432 2938
rect 20326 2857 20432 2874
rect 28416 3013 28522 3030
rect 28416 2949 28437 3013
rect 28501 2949 28522 3013
rect 28416 2933 28522 2949
rect 28416 2869 28437 2933
rect 28501 2869 28522 2933
rect 28416 2852 28522 2869
rect 28632 3013 28738 3030
rect 28632 2949 28653 3013
rect 28717 2949 28738 3013
rect 28632 2933 28738 2949
rect 28632 2869 28653 2933
rect 28717 2869 28738 2933
rect 28632 2852 28738 2869
rect 28848 3013 28954 3030
rect 28848 2949 28869 3013
rect 28933 2949 28954 3013
rect 28848 2933 28954 2949
rect 28848 2869 28869 2933
rect 28933 2869 28954 2933
rect 28848 2852 28954 2869
rect 41919 3015 42025 3032
rect 41919 2951 41940 3015
rect 42004 2951 42025 3015
rect 41919 2935 42025 2951
rect 41919 2871 41940 2935
rect 42004 2871 42025 2935
rect 41919 2854 42025 2871
rect 42135 3015 42241 3032
rect 42135 2951 42156 3015
rect 42220 2951 42241 3015
rect 42135 2935 42241 2951
rect 42135 2871 42156 2935
rect 42220 2871 42241 2935
rect 42135 2854 42241 2871
rect 42351 3015 42457 3032
rect 42351 2951 42372 3015
rect 42436 2951 42457 3015
rect 42351 2935 42457 2951
rect 42351 2871 42372 2935
rect 42436 2871 42457 2935
rect 42351 2854 42457 2871
rect 58414 3026 58520 3043
rect 58414 2962 58435 3026
rect 58499 2962 58520 3026
rect 58414 2946 58520 2962
rect 58414 2882 58435 2946
rect 58499 2882 58520 2946
rect 58414 2865 58520 2882
rect 58630 3026 58736 3043
rect 58630 2962 58651 3026
rect 58715 2962 58736 3026
rect 58630 2946 58736 2962
rect 58630 2882 58651 2946
rect 58715 2882 58736 2946
rect 58630 2865 58736 2882
rect 58846 3026 58952 3043
rect 58846 2962 58867 3026
rect 58931 2962 58952 3026
rect 58846 2946 58952 2962
rect 58846 2882 58867 2946
rect 58931 2882 58952 2946
rect 58846 2865 58952 2882
rect 4823 889 4929 906
rect 4823 825 4844 889
rect 4908 825 4929 889
rect 4823 809 4929 825
rect 4823 745 4844 809
rect 4908 745 4929 809
rect 4823 728 4929 745
rect 5044 889 5150 906
rect 5044 825 5065 889
rect 5129 825 5150 889
rect 5044 809 5150 825
rect 5044 745 5065 809
rect 5129 745 5150 809
rect 5044 728 5150 745
rect 5253 889 5359 906
rect 5253 825 5274 889
rect 5338 825 5359 889
rect 5253 809 5359 825
rect 5253 745 5274 809
rect 5338 745 5359 809
rect 5253 728 5359 745
rect 5427 889 5533 906
rect 5427 825 5448 889
rect 5512 825 5533 889
rect 16070 900 16147 903
rect 5427 809 5533 825
rect 5427 745 5448 809
rect 5512 745 5533 809
rect 8551 837 8637 851
rect 8551 773 8562 837
rect 8626 773 8637 837
rect 8551 760 8637 773
rect 8699 837 8785 851
rect 8699 773 8710 837
rect 8774 773 8785 837
rect 8699 760 8785 773
rect 8847 837 8933 851
rect 8847 773 8858 837
rect 8922 773 8933 837
rect 16070 836 16076 900
rect 16140 836 16147 900
rect 16070 834 16147 836
rect 21456 888 21562 905
rect 21456 824 21477 888
rect 21541 824 21562 888
rect 21456 808 21562 824
rect 8847 760 8933 773
rect 16093 781 16170 784
rect 5427 728 5533 745
rect 16093 717 16099 781
rect 16163 717 16170 781
rect 21456 744 21477 808
rect 21541 744 21562 808
rect 21456 727 21562 744
rect 21672 888 21778 905
rect 21672 824 21693 888
rect 21757 824 21778 888
rect 21672 808 21778 824
rect 21672 744 21693 808
rect 21757 744 21778 808
rect 21672 727 21778 744
rect 21888 888 21994 905
rect 21888 824 21909 888
rect 21973 824 21994 888
rect 29885 893 29991 910
rect 21888 808 21994 824
rect 21888 744 21909 808
rect 21973 744 21994 808
rect 23608 841 23704 863
rect 23608 777 23624 841
rect 23688 777 23704 841
rect 23608 755 23704 777
rect 23741 841 23837 863
rect 23741 777 23757 841
rect 23821 777 23837 841
rect 23741 755 23837 777
rect 23874 841 23970 863
rect 23874 777 23890 841
rect 23954 777 23970 841
rect 23874 755 23970 777
rect 29885 829 29906 893
rect 29970 829 29991 893
rect 29885 813 29991 829
rect 21888 727 21994 744
rect 29885 749 29906 813
rect 29970 749 29991 813
rect 29885 732 29991 749
rect 30101 893 30207 910
rect 30101 829 30122 893
rect 30186 829 30207 893
rect 30101 813 30207 829
rect 30101 749 30122 813
rect 30186 749 30207 813
rect 30101 732 30207 749
rect 30317 893 30423 910
rect 30317 829 30338 893
rect 30402 829 30423 893
rect 43403 883 43509 900
rect 30317 813 30423 829
rect 30317 749 30338 813
rect 30402 749 30423 813
rect 30317 732 30423 749
rect 32674 830 32761 854
rect 32674 766 32685 830
rect 32749 766 32761 830
rect 32674 742 32761 766
rect 32797 830 32884 854
rect 32797 766 32808 830
rect 32872 766 32884 830
rect 32797 742 32884 766
rect 32929 830 33016 854
rect 32929 766 32940 830
rect 33004 766 33016 830
rect 32929 742 33016 766
rect 38703 827 38790 851
rect 38703 763 38714 827
rect 38778 763 38790 827
rect 38703 739 38790 763
rect 38872 827 38959 851
rect 38872 763 38883 827
rect 38947 763 38959 827
rect 38872 739 38959 763
rect 43403 819 43424 883
rect 43488 819 43509 883
rect 43403 803 43509 819
rect 43403 739 43424 803
rect 43488 739 43509 803
rect 43403 722 43509 739
rect 43619 883 43725 900
rect 43619 819 43640 883
rect 43704 819 43725 883
rect 43619 803 43725 819
rect 43619 739 43640 803
rect 43704 739 43725 803
rect 43619 722 43725 739
rect 43835 883 43941 900
rect 55652 887 55736 894
rect 43835 819 43856 883
rect 43920 819 43941 883
rect 43835 803 43941 819
rect 43835 739 43856 803
rect 43920 739 43941 803
rect 43835 722 43941 739
rect 48329 877 48413 884
rect 48329 813 48339 877
rect 48403 813 48413 877
rect 48329 797 48413 813
rect 48329 733 48339 797
rect 48403 733 48413 797
rect 48329 726 48413 733
rect 48442 877 48526 884
rect 48442 813 48452 877
rect 48516 813 48526 877
rect 48442 797 48526 813
rect 48442 733 48452 797
rect 48516 733 48526 797
rect 48442 726 48526 733
rect 48557 877 48641 884
rect 48557 813 48567 877
rect 48631 813 48641 877
rect 48557 797 48641 813
rect 48557 733 48567 797
rect 48631 733 48641 797
rect 55652 823 55662 887
rect 55726 823 55736 887
rect 55652 807 55736 823
rect 55652 743 55662 807
rect 55726 743 55736 807
rect 55652 736 55736 743
rect 55771 887 55855 894
rect 55771 823 55781 887
rect 55845 823 55855 887
rect 55771 807 55855 823
rect 55771 743 55781 807
rect 55845 743 55855 807
rect 55771 736 55855 743
rect 55900 887 55984 894
rect 55900 823 55910 887
rect 55974 823 55984 887
rect 55900 807 55984 823
rect 55900 743 55910 807
rect 55974 743 55984 807
rect 55900 736 55984 743
rect 59915 878 60021 895
rect 59915 814 59936 878
rect 60000 814 60021 878
rect 59915 798 60021 814
rect 48557 726 48641 733
rect 59915 734 59936 798
rect 60000 734 60021 798
rect 59915 717 60021 734
rect 60131 878 60237 895
rect 60131 814 60152 878
rect 60216 814 60237 878
rect 60131 798 60237 814
rect 60131 734 60152 798
rect 60216 734 60237 798
rect 60131 717 60237 734
rect 60347 878 60453 895
rect 60347 814 60368 878
rect 60432 814 60453 878
rect 60347 798 60453 814
rect 60347 734 60368 798
rect 60432 734 60453 798
rect 60347 717 60453 734
rect 16093 715 16170 717
<< via3 >>
rect 4830 8002 4894 8066
rect 4830 7922 4894 7986
rect 5039 8001 5103 8065
rect 5039 7921 5103 7985
rect 5205 8001 5269 8065
rect 5205 7921 5269 7985
rect 5385 8003 5449 8067
rect 5385 7923 5449 7987
rect 21459 8019 21523 8083
rect 21459 7939 21523 8003
rect 21675 8019 21739 8083
rect 21675 7939 21739 8003
rect 21891 8019 21955 8083
rect 21891 7939 21955 8003
rect 29951 8018 30015 8082
rect 29951 7938 30015 8002
rect 30167 8018 30231 8082
rect 30167 7938 30231 8002
rect 30383 8018 30447 8082
rect 30383 7938 30447 8002
rect 43479 8024 43543 8088
rect 43479 7944 43543 8008
rect 43695 8024 43759 8088
rect 43695 7944 43759 8008
rect 43911 8024 43975 8088
rect 43911 7944 43975 8008
rect 59964 8017 60028 8081
rect 59964 7937 60028 8001
rect 60180 8017 60244 8081
rect 60180 7937 60244 8001
rect 60396 8017 60460 8081
rect 60396 7937 60460 8001
rect 3596 5884 3660 5948
rect 3768 5885 3832 5949
rect 3942 5884 4006 5948
rect 3596 5804 3660 5868
rect 3768 5805 3832 5869
rect 3942 5804 4006 5868
rect 19924 5905 19988 5969
rect 19924 5825 19988 5889
rect 20140 5905 20204 5969
rect 20140 5825 20204 5889
rect 20356 5905 20420 5969
rect 20356 5825 20420 5889
rect 28432 5897 28496 5961
rect 28432 5817 28496 5881
rect 28648 5897 28712 5961
rect 28648 5817 28712 5881
rect 28864 5897 28928 5961
rect 28864 5817 28928 5881
rect 41904 5892 41968 5956
rect 41904 5812 41968 5876
rect 42120 5892 42184 5956
rect 42120 5812 42184 5876
rect 42336 5892 42400 5956
rect 42336 5812 42400 5876
rect 58455 5884 58519 5948
rect 58455 5804 58519 5868
rect 58671 5884 58735 5948
rect 58671 5804 58735 5868
rect 58887 5884 58951 5948
rect 58887 5804 58951 5868
rect 38716 4181 38748 4202
rect 38748 4181 38780 4202
rect 38870 4181 38880 4203
rect 38880 4181 38934 4203
rect 38716 4149 38780 4181
rect 38870 4149 38934 4181
rect 38716 4138 38748 4149
rect 38748 4138 38780 4149
rect 38870 4139 38880 4149
rect 38880 4139 38934 4149
rect 8574 3895 8622 3909
rect 8622 3895 8638 3909
rect 8725 3895 8736 3915
rect 8736 3895 8789 3915
rect 8574 3845 8638 3895
rect 8725 3851 8789 3895
rect 8870 3851 8934 3915
rect 23617 3920 23661 3923
rect 23661 3920 23681 3923
rect 23784 3920 23813 3923
rect 23813 3920 23848 3923
rect 23617 3860 23681 3920
rect 23784 3860 23848 3920
rect 23617 3859 23661 3860
rect 23661 3859 23681 3860
rect 23784 3859 23813 3860
rect 23813 3859 23848 3860
rect 23617 3744 23681 3762
rect 23784 3744 23848 3762
rect 23617 3698 23661 3744
rect 23661 3698 23681 3744
rect 23784 3698 23813 3744
rect 23813 3698 23848 3744
rect 55656 3814 55695 3870
rect 55695 3814 55720 3870
rect 55777 3814 55799 3870
rect 55799 3814 55841 3870
rect 55915 3814 55951 3870
rect 55951 3814 55979 3870
rect 55656 3806 55720 3814
rect 55777 3806 55841 3814
rect 55915 3806 55979 3814
rect 55656 3780 55720 3790
rect 55777 3780 55841 3790
rect 55915 3780 55979 3790
rect 55656 3726 55695 3780
rect 55695 3726 55720 3780
rect 55777 3726 55799 3780
rect 55799 3726 55841 3780
rect 55915 3726 55951 3780
rect 55951 3726 55979 3780
rect 32664 3529 32728 3562
rect 32783 3529 32847 3562
rect 15950 3449 15960 3454
rect 15960 3449 16014 3454
rect 16053 3449 16068 3454
rect 16068 3449 16117 3454
rect 16156 3449 16176 3454
rect 16176 3449 16220 3454
rect 15950 3411 16014 3449
rect 16053 3411 16117 3449
rect 16156 3411 16220 3449
rect 32664 3498 32711 3529
rect 32711 3498 32728 3529
rect 32783 3498 32836 3529
rect 32836 3498 32847 3529
rect 32902 3529 32966 3562
rect 32902 3498 32905 3529
rect 32905 3498 32961 3529
rect 32961 3498 32966 3529
rect 48337 3478 48401 3494
rect 48477 3478 48541 3495
rect 48605 3478 48669 3495
rect 15950 3390 15960 3411
rect 15960 3390 16014 3411
rect 16053 3390 16068 3411
rect 16068 3390 16117 3411
rect 16156 3390 16176 3411
rect 16176 3390 16220 3411
rect 48337 3430 48382 3478
rect 48382 3430 48401 3478
rect 48477 3431 48512 3478
rect 48512 3431 48541 3478
rect 48605 3431 48661 3478
rect 48661 3431 48669 3478
rect 48337 3396 48401 3414
rect 48477 3396 48541 3415
rect 48605 3396 48669 3415
rect 48337 3350 48382 3396
rect 48382 3350 48401 3396
rect 48477 3351 48512 3396
rect 48512 3351 48541 3396
rect 48605 3351 48661 3396
rect 48661 3351 48669 3396
rect 3598 2936 3662 3000
rect 3598 2856 3662 2920
rect 3803 2938 3867 3002
rect 3803 2858 3867 2922
rect 4002 2938 4066 3002
rect 4002 2858 4066 2922
rect 19915 2954 19979 3018
rect 19915 2874 19979 2938
rect 20131 2954 20195 3018
rect 20131 2874 20195 2938
rect 20347 2954 20411 3018
rect 20347 2874 20411 2938
rect 28437 2949 28501 3013
rect 28437 2869 28501 2933
rect 28653 2949 28717 3013
rect 28653 2869 28717 2933
rect 28869 2949 28933 3013
rect 28869 2869 28933 2933
rect 41940 2951 42004 3015
rect 41940 2871 42004 2935
rect 42156 2951 42220 3015
rect 42156 2871 42220 2935
rect 42372 2951 42436 3015
rect 42372 2871 42436 2935
rect 58435 2962 58499 3026
rect 58435 2882 58499 2946
rect 58651 2962 58715 3026
rect 58651 2882 58715 2946
rect 58867 2962 58931 3026
rect 58867 2882 58931 2946
rect 4844 825 4908 889
rect 4844 745 4908 809
rect 5065 825 5129 889
rect 5065 745 5129 809
rect 5274 825 5338 889
rect 5274 745 5338 809
rect 5448 825 5512 889
rect 5448 745 5512 809
rect 8562 773 8626 837
rect 8710 773 8774 837
rect 8858 773 8922 837
rect 16076 836 16140 900
rect 21477 824 21541 888
rect 16099 717 16163 781
rect 21477 744 21541 808
rect 21693 824 21757 888
rect 21693 744 21757 808
rect 21909 824 21973 888
rect 21909 744 21973 808
rect 23624 777 23688 841
rect 23757 777 23821 841
rect 23890 777 23954 841
rect 29906 829 29970 893
rect 29906 749 29970 813
rect 30122 829 30186 893
rect 30122 749 30186 813
rect 30338 829 30402 893
rect 30338 749 30402 813
rect 32685 766 32749 830
rect 32808 766 32872 830
rect 32940 766 33004 830
rect 38714 763 38778 827
rect 38883 763 38947 827
rect 43424 819 43488 883
rect 43424 739 43488 803
rect 43640 819 43704 883
rect 43640 739 43704 803
rect 43856 819 43920 883
rect 43856 739 43920 803
rect 48339 813 48403 877
rect 48339 733 48403 797
rect 48452 813 48516 877
rect 48452 733 48516 797
rect 48567 813 48631 877
rect 48567 733 48631 797
rect 55662 823 55726 887
rect 55662 743 55726 807
rect 55781 823 55845 887
rect 55781 743 55845 807
rect 55910 823 55974 887
rect 55910 743 55974 807
rect 59936 814 60000 878
rect 59936 734 60000 798
rect 60152 814 60216 878
rect 60152 734 60216 798
rect 60368 814 60432 878
rect 60368 734 60432 798
<< metal4 >>
rect 3431 5949 4237 8265
rect 3431 5948 3768 5949
rect 3431 5884 3596 5948
rect 3660 5885 3768 5948
rect 3832 5948 4237 5949
rect 3832 5885 3942 5948
rect 3660 5884 3942 5885
rect 4006 5884 4237 5948
rect 3431 5869 4237 5884
rect 3431 5868 3768 5869
rect 3431 5804 3596 5868
rect 3660 5805 3768 5868
rect 3832 5868 4237 5869
rect 3832 5805 3942 5868
rect 3660 5804 3942 5805
rect 4006 5804 4237 5868
rect 3431 3002 4237 5804
rect 3431 3000 3803 3002
rect 3431 2936 3598 3000
rect 3662 2938 3803 3000
rect 3867 2938 4002 3002
rect 4066 2938 4237 3002
rect 3662 2936 4237 2938
rect 3431 2922 4237 2936
rect 3431 2920 3803 2922
rect 3431 2856 3598 2920
rect 3662 2858 3803 2920
rect 3867 2858 4002 2922
rect 4066 2858 4237 2922
rect 3662 2856 4237 2858
rect 3431 559 4237 2856
rect 4774 8067 5580 8266
rect 4774 8066 5385 8067
rect 4774 8002 4830 8066
rect 4894 8065 5385 8066
rect 4894 8002 5039 8065
rect 4774 8001 5039 8002
rect 5103 8001 5205 8065
rect 5269 8003 5385 8065
rect 5449 8003 5580 8067
rect 5269 8001 5580 8003
rect 4774 7987 5580 8001
rect 4774 7986 5385 7987
rect 4774 7922 4830 7986
rect 4894 7985 5385 7986
rect 4894 7922 5039 7985
rect 4774 7921 5039 7922
rect 5103 7921 5205 7985
rect 5269 7923 5385 7985
rect 5449 7923 5580 7987
rect 5269 7921 5580 7923
rect 4774 889 5580 7921
rect 19774 5969 20580 8266
rect 19774 5905 19924 5969
rect 19988 5905 20140 5969
rect 20204 5905 20356 5969
rect 20420 5905 20580 5969
rect 19774 5889 20580 5905
rect 19774 5825 19924 5889
rect 19988 5825 20140 5889
rect 20204 5825 20356 5889
rect 20420 5825 20580 5889
rect 4774 825 4844 889
rect 4908 825 5065 889
rect 5129 825 5274 889
rect 5338 825 5448 889
rect 5512 825 5580 889
rect 4774 809 5580 825
rect 4774 745 4844 809
rect 4908 745 5065 809
rect 5129 745 5274 809
rect 5338 745 5448 809
rect 5512 745 5580 809
rect 4774 560 5580 745
rect 8505 3915 8974 4044
rect 8505 3909 8725 3915
rect 8505 3845 8574 3909
rect 8638 3851 8725 3909
rect 8789 3851 8870 3915
rect 8934 3851 8974 3915
rect 8638 3845 8974 3851
rect 8505 837 8974 3845
rect 15920 3454 16274 3529
rect 15920 3390 15950 3454
rect 16014 3390 16053 3454
rect 16117 3390 16156 3454
rect 16220 3390 16274 3454
rect 15920 3328 16274 3390
rect 8505 773 8562 837
rect 8626 773 8710 837
rect 8774 773 8858 837
rect 8922 773 8974 837
rect 8505 661 8974 773
rect 15996 900 16197 3328
rect 15996 836 16076 900
rect 16140 836 16197 900
rect 15996 781 16197 836
rect 15996 717 16099 781
rect 16163 717 16197 781
rect 15996 636 16197 717
rect 19774 3018 20580 5825
rect 19774 2954 19915 3018
rect 19979 2954 20131 3018
rect 20195 2954 20347 3018
rect 20411 2954 20580 3018
rect 19774 2938 20580 2954
rect 19774 2874 19915 2938
rect 19979 2874 20131 2938
rect 20195 2874 20347 2938
rect 20411 2874 20580 2938
rect 19774 560 20580 2874
rect 21274 8083 22080 8266
rect 21274 8019 21459 8083
rect 21523 8019 21675 8083
rect 21739 8019 21891 8083
rect 21955 8019 22080 8083
rect 21274 8003 22080 8019
rect 21274 7939 21459 8003
rect 21523 7939 21675 8003
rect 21739 7939 21891 8003
rect 21955 7939 22080 8003
rect 21274 888 22080 7939
rect 28274 5961 29080 8266
rect 28274 5897 28432 5961
rect 28496 5897 28648 5961
rect 28712 5897 28864 5961
rect 28928 5897 29080 5961
rect 28274 5881 29080 5897
rect 28274 5817 28432 5881
rect 28496 5817 28648 5881
rect 28712 5817 28864 5881
rect 28928 5817 29080 5881
rect 21274 824 21477 888
rect 21541 824 21693 888
rect 21757 824 21909 888
rect 21973 824 22080 888
rect 21274 808 22080 824
rect 21274 744 21477 808
rect 21541 744 21693 808
rect 21757 744 21909 808
rect 21973 744 22080 808
rect 21274 560 22080 744
rect 23555 3923 24022 4058
rect 23555 3859 23617 3923
rect 23681 3859 23784 3923
rect 23848 3859 24022 3923
rect 23555 3762 24022 3859
rect 23555 3698 23617 3762
rect 23681 3698 23784 3762
rect 23848 3698 24022 3762
rect 23555 841 24022 3698
rect 23555 777 23624 841
rect 23688 777 23757 841
rect 23821 777 23890 841
rect 23954 777 24022 841
rect 23555 686 24022 777
rect 28274 3013 29080 5817
rect 28274 2949 28437 3013
rect 28501 2949 28653 3013
rect 28717 2949 28869 3013
rect 28933 2949 29080 3013
rect 28274 2933 29080 2949
rect 28274 2869 28437 2933
rect 28501 2869 28653 2933
rect 28717 2869 28869 2933
rect 28933 2869 29080 2933
rect 28274 560 29080 2869
rect 29774 8082 30580 8266
rect 29774 8018 29951 8082
rect 30015 8018 30167 8082
rect 30231 8018 30383 8082
rect 30447 8018 30580 8082
rect 29774 8002 30580 8018
rect 29774 7938 29951 8002
rect 30015 7938 30167 8002
rect 30231 7938 30383 8002
rect 30447 7938 30580 8002
rect 29774 893 30580 7938
rect 41774 5956 42580 8266
rect 41774 5892 41904 5956
rect 41968 5892 42120 5956
rect 42184 5892 42336 5956
rect 42400 5892 42580 5956
rect 41774 5876 42580 5892
rect 41774 5812 41904 5876
rect 41968 5812 42120 5876
rect 42184 5812 42336 5876
rect 42400 5812 42580 5876
rect 38669 4203 38974 4384
rect 38669 4202 38870 4203
rect 38669 4138 38716 4202
rect 38780 4139 38870 4202
rect 38934 4139 38974 4203
rect 38780 4138 38974 4139
rect 29774 829 29906 893
rect 29970 829 30122 893
rect 30186 829 30338 893
rect 30402 829 30580 893
rect 29774 813 30580 829
rect 29774 749 29906 813
rect 29970 749 30122 813
rect 30186 749 30338 813
rect 30402 749 30580 813
rect 29774 560 30580 749
rect 32607 3562 33032 3665
rect 32607 3498 32664 3562
rect 32728 3498 32783 3562
rect 32847 3498 32902 3562
rect 32966 3498 33032 3562
rect 32607 830 33032 3498
rect 32607 766 32685 830
rect 32749 766 32808 830
rect 32872 766 32940 830
rect 33004 766 33032 830
rect 32607 700 33032 766
rect 38669 827 38974 4138
rect 38669 763 38714 827
rect 38778 763 38883 827
rect 38947 763 38974 827
rect 38669 691 38974 763
rect 41774 3015 42580 5812
rect 41774 2951 41940 3015
rect 42004 2951 42156 3015
rect 42220 2951 42372 3015
rect 42436 2951 42580 3015
rect 41774 2935 42580 2951
rect 41774 2871 41940 2935
rect 42004 2871 42156 2935
rect 42220 2871 42372 2935
rect 42436 2871 42580 2935
rect 41774 560 42580 2871
rect 43274 8088 44080 8266
rect 43274 8024 43479 8088
rect 43543 8024 43695 8088
rect 43759 8024 43911 8088
rect 43975 8024 44080 8088
rect 43274 8008 44080 8024
rect 43274 7944 43479 8008
rect 43543 7944 43695 8008
rect 43759 7944 43911 8008
rect 43975 7944 44080 8008
rect 43274 883 44080 7944
rect 58274 5948 59080 8266
rect 58274 5884 58455 5948
rect 58519 5884 58671 5948
rect 58735 5884 58887 5948
rect 58951 5884 59080 5948
rect 58274 5868 59080 5884
rect 58274 5804 58455 5868
rect 58519 5804 58671 5868
rect 58735 5804 58887 5868
rect 58951 5804 59080 5868
rect 55602 3870 56027 3900
rect 55602 3806 55656 3870
rect 55720 3806 55777 3870
rect 55841 3806 55915 3870
rect 55979 3806 56027 3870
rect 55602 3790 56027 3806
rect 55602 3726 55656 3790
rect 55720 3726 55777 3790
rect 55841 3726 55915 3790
rect 55979 3726 56027 3790
rect 43274 819 43424 883
rect 43488 819 43640 883
rect 43704 819 43856 883
rect 43920 819 44080 883
rect 43274 803 44080 819
rect 43274 739 43424 803
rect 43488 739 43640 803
rect 43704 739 43856 803
rect 43920 739 44080 803
rect 43274 560 44080 739
rect 48289 3495 48703 3591
rect 48289 3494 48477 3495
rect 48289 3430 48337 3494
rect 48401 3431 48477 3494
rect 48541 3431 48605 3495
rect 48669 3431 48703 3495
rect 48401 3430 48703 3431
rect 48289 3415 48703 3430
rect 48289 3414 48477 3415
rect 48289 3350 48337 3414
rect 48401 3351 48477 3414
rect 48541 3351 48605 3415
rect 48669 3351 48703 3415
rect 48401 3350 48703 3351
rect 48289 877 48703 3350
rect 48289 813 48339 877
rect 48403 813 48452 877
rect 48516 813 48567 877
rect 48631 813 48703 877
rect 48289 797 48703 813
rect 48289 733 48339 797
rect 48403 733 48452 797
rect 48516 733 48567 797
rect 48631 733 48703 797
rect 48289 638 48703 733
rect 55602 887 56027 3726
rect 55602 823 55662 887
rect 55726 823 55781 887
rect 55845 823 55910 887
rect 55974 823 56027 887
rect 55602 807 56027 823
rect 55602 743 55662 807
rect 55726 743 55781 807
rect 55845 743 55910 807
rect 55974 743 56027 807
rect 55602 650 56027 743
rect 58274 3026 59080 5804
rect 58274 2962 58435 3026
rect 58499 2962 58651 3026
rect 58715 2962 58867 3026
rect 58931 2962 59080 3026
rect 58274 2946 59080 2962
rect 58274 2882 58435 2946
rect 58499 2882 58651 2946
rect 58715 2882 58867 2946
rect 58931 2882 59080 2946
rect 58274 560 59080 2882
rect 59774 8081 60580 8266
rect 59774 8017 59964 8081
rect 60028 8017 60180 8081
rect 60244 8017 60396 8081
rect 60460 8017 60580 8081
rect 59774 8001 60580 8017
rect 59774 7937 59964 8001
rect 60028 7937 60180 8001
rect 60244 7937 60396 8001
rect 60460 7937 60580 8001
rect 59774 878 60580 7937
rect 59774 814 59936 878
rect 60000 814 60152 878
rect 60216 814 60368 878
rect 60432 814 60580 878
rect 59774 798 60580 814
rect 59774 734 59936 798
rect 60000 734 60152 798
rect 60216 734 60368 798
rect 60432 734 60580 798
rect 59774 560 60580 734
use brbufhalf  brbufhalf_0
timestamp 1655322987
transform -1 0 58721 0 -1 10662
box -3552 2527 26658 5446
use brbufhalf  brbufhalf_1
timestamp 1655322987
transform 1 0 36045 0 1 -1834
box -3552 2527 26658 5446
use brbufhalf  brbufhalf_2
timestamp 1655322987
transform 1 0 5843 0 1 -1834
box -3552 2527 26658 5446
use brbufhalf_64  brbufhalf_64_0
timestamp 1655322987
transform -1 0 28519 0 -1 10662
box -3552 2527 26308 5446
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0
timestamp 1655322987
transform 1 0 32318 0 1 4265
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0
timestamp 1655322987
transform 1 0 45672 0 1 4049
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1655322987
transform 1 0 47602 0 1 4049
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_2
timestamp 1655322987
transform 1 0 32866 0 1 4265
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_3
timestamp 1655322987
transform 1 0 15530 0 1 3889
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_4
timestamp 1655322987
transform 1 0 17460 0 1 3889
box -38 -48 1510 592
use unitcell2buf  unitcell2buf_0
timestamp 1655322987
transform 1 0 977 0 1 1878
box -574 -1185 1322 1192
<< labels >>
flabel metal1 s 62673 1474 62895 1552 1 FreeSans 2000 0 0 0 OUT
port 1 nsew
flabel metal4 s 3431 559 4237 8265 1 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal4 s 19774 560 20580 8266 1 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal4 s 28274 560 29080 8266 1 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal4 s 41774 560 42580 8266 1 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal4 s 58274 560 59080 8266 1 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal4 s 4774 560 5580 8266 1 FreeSans 2000 0 0 0 VSS
port 3 nsew
flabel metal4 s 21274 560 22080 8266 1 FreeSans 2000 0 0 0 VSS
port 3 nsew
flabel metal4 s 29774 560 30580 8266 1 FreeSans 2000 0 0 0 VSS
port 3 nsew
flabel metal4 s 43274 560 44080 8266 1 FreeSans 2000 0 0 0 VSS
port 3 nsew
flabel metal4 s 59774 560 60580 8266 1 FreeSans 2000 0 0 0 VSS
port 3 nsew
flabel metal1 s 0 4626 534 4690 1 FreeSans 2000 0 0 0 RESET
port 4 nsew
flabel metal2 s 62209 7342 62253 8498 1 FreeSans 2000 0 0 0 C[0]
port 5 nsew
flabel metal2 s 60321 7342 60365 8498 1 FreeSans 2000 0 0 0 C[1]
port 6 nsew
flabel metal2 s 58433 7342 58477 8498 1 FreeSans 2000 0 0 0 C[2]
port 7 nsew
flabel metal2 s 56545 7342 56589 8498 1 FreeSans 2000 0 0 0 C[3]
port 8 nsew
flabel metal2 s 54657 7342 54701 8498 1 FreeSans 2000 0 0 0 C[4]
port 9 nsew
flabel metal2 s 52769 7342 52813 8498 1 FreeSans 2000 0 0 0 C[5]
port 10 nsew
flabel metal2 s 50881 7342 50925 8498 1 FreeSans 2000 0 0 0 C[6]
port 11 nsew
flabel metal2 s 48993 7342 49037 8498 1 FreeSans 2000 0 0 0 C[7]
port 12 nsew
flabel metal2 s 47105 7342 47149 8498 1 FreeSans 2000 0 0 0 C[8]
port 13 nsew
flabel metal2 s 45217 7342 45261 8498 1 FreeSans 2000 0 0 0 C[9]
port 14 nsew
flabel metal2 s 43329 7342 43373 8498 1 FreeSans 2000 0 0 0 C[10]
port 15 nsew
flabel metal2 s 41441 7342 41485 8498 1 FreeSans 2000 0 0 0 C[11]
port 16 nsew
flabel metal2 s 39553 7342 39597 8498 1 FreeSans 2000 0 0 0 C[12]
port 17 nsew
flabel metal2 s 37665 7342 37709 8498 1 FreeSans 2000 0 0 0 C[13]
port 18 nsew
flabel metal2 s 35777 7342 35821 8498 1 FreeSans 2000 0 0 0 C[14]
port 19 nsew
flabel metal2 s 33889 7342 33933 8498 1 FreeSans 2000 0 0 0 C[15]
port 20 nsew
flabel metal2 s 32001 7342 32045 8498 1 FreeSans 2000 0 0 0 C[16]
port 21 nsew
flabel metal2 s 30113 7342 30157 8498 1 FreeSans 2000 0 0 0 C[17]
port 22 nsew
flabel metal2 s 28225 7342 28269 8498 1 FreeSans 2000 0 0 0 C[18]
port 23 nsew
flabel metal2 s 26337 7342 26381 8498 1 FreeSans 2000 0 0 0 C[19]
port 24 nsew
flabel metal2 s 24449 7342 24493 8498 1 FreeSans 2000 0 0 0 C[20]
port 25 nsew
flabel metal2 s 22561 7342 22605 8498 1 FreeSans 2000 0 0 0 C[21]
port 26 nsew
flabel metal2 s 20673 7342 20717 8498 1 FreeSans 2000 0 0 0 C[22]
port 27 nsew
flabel metal2 s 18785 7342 18829 8498 1 FreeSans 2000 0 0 0 C[23]
port 28 nsew
flabel metal2 s 16897 7342 16941 8498 1 FreeSans 2000 0 0 0 C[24]
port 29 nsew
flabel metal2 s 15009 7342 15053 8498 1 FreeSans 2000 0 0 0 C[25]
port 30 nsew
flabel metal2 s 13121 7342 13165 8498 1 FreeSans 2000 0 0 0 C[26]
port 31 nsew
flabel metal2 s 11233 7342 11277 8498 1 FreeSans 2000 0 0 0 C[27]
port 32 nsew
flabel metal2 s 9345 7342 9389 8498 1 FreeSans 2000 0 0 0 C[28]
port 33 nsew
flabel metal2 s 7457 7342 7501 8498 1 FreeSans 2000 0 0 0 C[29]
port 34 nsew
flabel metal2 s 5569 7342 5613 8498 1 FreeSans 2000 0 0 0 C[30]
port 35 nsew
flabel metal2 s 422 22 467 1168 1 FreeSans 2000 0 0 0 C[31]
port 36 nsew
flabel metal2 s 2310 22 2355 1168 1 FreeSans 2000 0 0 0 C[32]
port 37 nsew
flabel metal2 s 4198 22 4243 1168 1 FreeSans 2000 0 0 0 C[33]
port 38 nsew
flabel metal2 s 6086 22 6131 1168 1 FreeSans 2000 0 0 0 C[34]
port 39 nsew
flabel metal2 s 7974 22 8019 1168 1 FreeSans 2000 0 0 0 C[35]
port 40 nsew
flabel metal2 s 9862 22 9907 1168 1 FreeSans 2000 0 0 0 C[36]
port 41 nsew
flabel metal2 s 11750 22 11795 1168 1 FreeSans 2000 0 0 0 C[37]
port 42 nsew
flabel metal2 s 13638 22 13683 1168 1 FreeSans 2000 0 0 0 C[38]
port 43 nsew
flabel metal2 s 15526 22 15571 1168 1 FreeSans 2000 0 0 0 C[39]
port 44 nsew
flabel metal2 s 17414 22 17459 1168 1 FreeSans 2000 0 0 0 C[40]
port 45 nsew
flabel metal2 s 19302 22 19347 1168 1 FreeSans 2000 0 0 0 C[41]
port 46 nsew
flabel metal2 s 21190 22 21235 1168 1 FreeSans 2000 0 0 0 C[42]
port 47 nsew
flabel metal2 s 23078 22 23123 1168 1 FreeSans 2000 0 0 0 C[43]
port 48 nsew
flabel metal2 s 24966 22 25011 1168 1 FreeSans 2000 0 0 0 C[44]
port 49 nsew
flabel metal2 s 26854 22 26899 1168 1 FreeSans 2000 0 0 0 C[45]
port 50 nsew
flabel metal2 s 28742 22 28787 1168 1 FreeSans 2000 0 0 0 C[46]
port 51 nsew
flabel metal2 s 30630 22 30675 1168 1 FreeSans 2000 0 0 0 C[47]
port 52 nsew
flabel metal2 s 32518 22 32563 1168 1 FreeSans 2000 0 0 0 C[48]
port 53 nsew
flabel metal2 s 34406 22 34451 1168 1 FreeSans 2000 0 0 0 C[49]
port 54 nsew
flabel metal2 s 36294 22 36339 1168 1 FreeSans 2000 0 0 0 C[50]
port 55 nsew
flabel metal2 s 38182 22 38227 1168 1 FreeSans 2000 0 0 0 C[51]
port 56 nsew
flabel metal2 s 40070 22 40115 1168 1 FreeSans 2000 0 0 0 C[52]
port 57 nsew
flabel metal2 s 41958 22 42003 1168 1 FreeSans 2000 0 0 0 C[53]
port 58 nsew
flabel metal2 s 43846 22 43891 1168 1 FreeSans 2000 0 0 0 C[54]
port 59 nsew
flabel metal2 s 45734 22 45779 1168 1 FreeSans 2000 0 0 0 C[55]
port 60 nsew
flabel metal2 s 47622 22 47667 1168 1 FreeSans 2000 0 0 0 C[56]
port 61 nsew
flabel metal2 s 49510 22 49555 1168 1 FreeSans 2000 0 0 0 C[57]
port 62 nsew
flabel metal2 s 51398 22 51443 1168 1 FreeSans 2000 0 0 0 C[58]
port 63 nsew
flabel metal2 s 53286 22 53331 1168 1 FreeSans 2000 0 0 0 C[59]
port 64 nsew
flabel metal2 s 55174 22 55219 1168 1 FreeSans 2000 0 0 0 C[60]
port 65 nsew
flabel metal2 s 57062 22 57107 1168 1 FreeSans 2000 0 0 0 C[61]
port 66 nsew
flabel metal2 s 58950 22 58995 1168 1 FreeSans 2000 0 0 0 C[62]
port 67 nsew
flabel metal2 s 60827 0 60883 1486 1 FreeSans 2000 0 0 0 C[63]
port 68 nsew
<< end >>
