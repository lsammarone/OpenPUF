magic
tech sky130A
magscale 1 2
timestamp 1483428465
<< checkpaint >>
rect -2434 -1440 2433 1440
<< metal3 >>
rect -1174 152 1173 180
rect -1174 -152 -1152 152
rect 1152 -152 1173 152
rect -1174 -180 1173 -152
<< via3 >>
rect -1152 -152 1152 152
<< metal4 >>
rect -1174 152 1173 180
rect -1174 -152 -1152 152
rect 1152 -152 1173 152
rect -1174 -180 1173 -152
<< end >>
