magic
tech sky130A
magscale 1 2
timestamp 1654736712
<< metal4 >>
rect -169 918 169 1000
rect -169 682 -118 918
rect 118 682 169 918
rect -169 598 169 682
rect -169 362 -118 598
rect 118 362 169 598
rect -169 278 169 362
rect -169 42 -118 278
rect 118 42 169 278
rect -169 -42 169 42
rect -169 -278 -118 -42
rect 118 -278 169 -42
rect -169 -362 169 -278
rect -169 -598 -118 -362
rect 118 -598 169 -362
rect -169 -682 169 -598
rect -169 -918 -118 -682
rect 118 -918 169 -682
rect -169 -1000 169 -918
<< via4 >>
rect -118 682 118 918
rect -118 362 118 598
rect -118 42 118 278
rect -118 -278 118 -42
rect -118 -598 118 -362
rect -118 -918 118 -682
<< metal5 >>
rect -169 918 169 1000
rect -169 682 -118 918
rect 118 682 169 918
rect -169 598 169 682
rect -169 362 -118 598
rect 118 362 169 598
rect -169 278 169 362
rect -169 42 -118 278
rect 118 42 169 278
rect -169 -42 169 42
rect -169 -278 -118 -42
rect 118 -278 169 -42
rect -169 -362 169 -278
rect -169 -598 -118 -362
rect 118 -598 169 -362
rect -169 -682 169 -598
rect -169 -918 -118 -682
rect 118 -918 169 -682
rect -169 -1000 169 -918
<< end >>
