magic
tech sky130A
magscale 1 2
timestamp 1656715967
<< nwell >>
rect 33226 5925 34010 6074
rect 33246 4847 33624 5925
rect 32979 4818 33624 4847
rect 32979 4526 33515 4818
rect 17259 4150 17641 4471
rect 47401 4310 47783 4631
<< nsubdiff >>
rect 47526 4483 47660 4502
rect 47526 4449 47598 4483
rect 47632 4449 47660 4483
rect 47526 4432 47660 4449
rect 17384 4323 17518 4342
rect 17384 4289 17456 4323
rect 17490 4289 17518 4323
rect 17384 4272 17518 4289
<< nsubdiffcont >>
rect 47598 4449 47632 4483
rect 17456 4289 17490 4323
<< locali >>
rect 32221 4524 32577 4530
rect 32221 4490 32268 4524
rect 32302 4490 32356 4524
rect 32390 4490 32577 4524
rect 32221 4480 32577 4490
rect 47323 4483 47866 4503
rect 47323 4449 47598 4483
rect 47632 4449 47866 4483
rect 47323 4431 47866 4449
rect 46192 4409 46226 4415
rect 46024 4402 46058 4408
rect 46528 4411 46562 4417
rect 46192 4370 46226 4375
rect 46360 4399 46394 4405
rect 46024 4363 46058 4368
rect 46528 4372 46562 4377
rect 46694 4409 46728 4415
rect 46694 4370 46728 4375
rect 46860 4411 46894 4417
rect 46860 4372 46894 4377
rect 47028 4411 47062 4417
rect 47028 4372 47062 4377
rect 47202 4409 47236 4415
rect 47202 4370 47236 4375
rect 47958 4403 47992 4409
rect 46360 4360 46394 4365
rect 47958 4364 47992 4369
rect 48120 4407 48154 4413
rect 48120 4368 48154 4373
rect 48290 4411 48324 4417
rect 48290 4372 48324 4377
rect 48454 4407 48488 4413
rect 48454 4368 48488 4373
rect 48624 4407 48658 4413
rect 48624 4368 48658 4373
rect 48792 4403 48826 4409
rect 48792 4364 48826 4369
rect 48960 4407 48994 4413
rect 48960 4368 48994 4373
rect 49134 4403 49168 4409
rect 49134 4364 49168 4369
rect 17181 4323 17724 4343
rect 17181 4289 17456 4323
rect 17490 4289 17724 4323
rect 17181 4271 17724 4289
rect 16050 4249 16084 4255
rect 15882 4242 15916 4248
rect 16386 4251 16420 4257
rect 16050 4210 16084 4215
rect 16218 4239 16252 4245
rect 15882 4203 15916 4208
rect 16386 4212 16420 4217
rect 16552 4249 16586 4255
rect 16552 4210 16586 4215
rect 16718 4251 16752 4257
rect 16718 4212 16752 4217
rect 16886 4251 16920 4257
rect 16886 4212 16920 4217
rect 17060 4249 17094 4255
rect 17060 4210 17094 4215
rect 17816 4243 17850 4249
rect 16218 4200 16252 4205
rect 17816 4204 17850 4209
rect 17978 4247 18012 4253
rect 17978 4208 18012 4213
rect 18148 4251 18182 4257
rect 18148 4212 18182 4217
rect 18312 4247 18346 4253
rect 18312 4208 18346 4213
rect 18482 4247 18516 4253
rect 18482 4208 18516 4213
rect 18650 4243 18684 4249
rect 18650 4204 18684 4209
rect 18818 4247 18852 4253
rect 18818 4208 18852 4213
rect 18992 4243 19026 4249
rect 18992 4204 19026 4209
<< viali >>
rect 32268 4490 32302 4524
rect 32356 4490 32390 4524
rect 32933 4522 32967 4556
rect 33204 4486 33238 4520
rect 33292 4486 33326 4520
rect 33380 4486 33414 4520
rect 33468 4486 33502 4520
rect 33556 4486 33590 4520
rect 33644 4486 33678 4520
rect 33732 4486 33766 4520
rect 33820 4486 33854 4520
rect 32933 4442 32967 4476
rect 33558 4384 33592 4418
rect 33724 4380 33758 4414
rect 33892 4386 33926 4420
rect 34059 4384 34093 4418
rect 34229 4385 34263 4419
rect 34393 4386 34427 4420
rect 46024 4368 46058 4402
rect 46192 4375 46226 4409
rect 46360 4365 46394 4399
rect 46528 4377 46562 4411
rect 46694 4375 46728 4409
rect 46860 4377 46894 4411
rect 47028 4377 47062 4411
rect 47202 4375 47236 4409
rect 47958 4369 47992 4403
rect 48120 4373 48154 4407
rect 48290 4377 48324 4411
rect 48454 4373 48488 4407
rect 48624 4373 48658 4407
rect 48792 4369 48826 4403
rect 48960 4373 48994 4407
rect 49134 4369 49168 4403
rect 46224 4272 46258 4306
rect 46324 4272 46358 4306
rect 46424 4272 46458 4306
rect 46524 4272 46558 4306
rect 46624 4272 46658 4306
rect 46724 4272 46758 4306
rect 46824 4272 46858 4306
rect 46924 4272 46958 4306
rect 47884 4272 47918 4306
rect 47984 4272 48018 4306
rect 48084 4272 48118 4306
rect 48184 4272 48218 4306
rect 48284 4272 48318 4306
rect 48384 4272 48418 4306
rect 48484 4272 48518 4306
rect 48584 4272 48618 4306
rect 15882 4208 15916 4242
rect 16050 4215 16084 4249
rect 16218 4205 16252 4239
rect 16386 4217 16420 4251
rect 16552 4215 16586 4249
rect 16718 4217 16752 4251
rect 16886 4217 16920 4251
rect 17060 4215 17094 4249
rect 17816 4209 17850 4243
rect 17978 4213 18012 4247
rect 18148 4217 18182 4251
rect 18312 4213 18346 4247
rect 18482 4213 18516 4247
rect 18650 4209 18684 4243
rect 18818 4213 18852 4247
rect 18992 4209 19026 4243
rect 16082 4112 16116 4146
rect 16182 4112 16216 4146
rect 16282 4112 16316 4146
rect 16382 4112 16416 4146
rect 16482 4112 16516 4146
rect 16582 4112 16616 4146
rect 16682 4112 16716 4146
rect 16782 4112 16816 4146
rect 17742 4112 17776 4146
rect 17842 4112 17876 4146
rect 17942 4112 17976 4146
rect 18042 4112 18076 4146
rect 18142 4112 18176 4146
rect 18242 4112 18276 4146
rect 18342 4112 18376 4146
rect 18442 4112 18476 4146
<< metal1 >>
rect 16933 5441 17188 5797
rect 32869 5464 33203 5788
rect 16933 5389 16953 5441
rect 17005 5389 17031 5441
rect 17083 5389 17124 5441
rect 17176 5389 17188 5441
rect 16933 5359 17188 5389
rect 32869 5412 32912 5464
rect 32964 5412 33025 5464
rect 33077 5412 33126 5464
rect 33178 5412 33203 5464
rect 32869 5368 33203 5412
rect 47073 5441 47300 5809
rect 47073 5389 47104 5441
rect 47156 5389 47187 5441
rect 47239 5389 47300 5441
rect 47073 5355 47300 5389
rect 9589 5224 10125 5308
rect 24623 5233 25231 5291
rect 39727 5241 40351 5299
rect 54733 5247 55466 5305
rect 32997 4844 33105 4857
rect 32997 4792 33027 4844
rect 33079 4792 33105 4844
rect 32997 4761 33105 4792
rect 34537 4761 34572 4857
rect 220 4690 19603 4691
rect 219 4626 19603 4690
rect 220 4625 19603 4626
rect 19537 4539 19603 4625
rect 47242 4617 47909 4626
rect 32918 4556 32997 4584
rect 47252 4568 47909 4617
rect 19537 4524 32484 4539
rect 19537 4490 32268 4524
rect 32302 4490 32356 4524
rect 32390 4490 32484 4524
rect 19537 4473 32484 4490
rect 32918 4522 32933 4556
rect 32967 4528 32997 4556
rect 32967 4522 33916 4528
rect 32918 4520 33916 4522
rect 32918 4486 33204 4520
rect 33238 4486 33292 4520
rect 33326 4486 33380 4520
rect 33414 4486 33468 4520
rect 33502 4486 33556 4520
rect 33590 4486 33644 4520
rect 33678 4486 33732 4520
rect 33766 4486 33820 4520
rect 33854 4486 33916 4520
rect 32918 4480 33916 4486
rect 32918 4476 33000 4480
rect 17152 4412 17801 4462
rect 32918 4442 32933 4476
rect 32967 4442 33000 4476
rect 32918 4424 33000 4442
rect 33489 4435 34434 4448
rect 17100 4404 17801 4412
rect 33489 4418 33705 4435
rect 33489 4384 33558 4418
rect 33592 4384 33705 4418
rect 33757 4414 33865 4435
rect 33917 4420 33998 4435
rect 33489 4383 33705 4384
rect 33758 4383 33865 4414
rect 33926 4386 33998 4420
rect 33917 4383 33998 4386
rect 34050 4418 34111 4435
rect 34050 4384 34059 4418
rect 34093 4384 34111 4418
rect 34050 4383 34111 4384
rect 34163 4420 34434 4435
rect 34163 4419 34393 4420
rect 34163 4385 34229 4419
rect 34263 4386 34393 4419
rect 34427 4386 34434 4420
rect 34263 4385 34434 4386
rect 34163 4383 34434 4385
rect 33489 4380 33724 4383
rect 33758 4380 34434 4383
rect 33489 4365 34434 4380
rect 39891 4411 55326 4427
rect 39891 4409 46528 4411
rect 39891 4408 46192 4409
rect 39891 4407 40073 4408
rect 39891 4355 39970 4407
rect 40022 4356 40073 4407
rect 40125 4402 46192 4408
rect 40125 4368 46024 4402
rect 46058 4375 46192 4402
rect 46226 4399 46528 4409
rect 46226 4375 46360 4399
rect 46058 4368 46360 4375
rect 40125 4365 46360 4368
rect 46394 4377 46528 4399
rect 46562 4409 46860 4411
rect 46562 4377 46694 4409
rect 46394 4375 46694 4377
rect 46728 4377 46860 4409
rect 46894 4377 47028 4411
rect 47062 4409 48290 4411
rect 47062 4377 47202 4409
rect 46728 4375 47202 4377
rect 47236 4407 48290 4409
rect 47236 4403 48120 4407
rect 47236 4375 47958 4403
rect 46394 4369 47958 4375
rect 47992 4373 48120 4403
rect 48154 4377 48290 4407
rect 48324 4408 55326 4411
rect 48324 4407 55174 4408
rect 48324 4377 48454 4407
rect 48154 4373 48454 4377
rect 48488 4373 48624 4407
rect 48658 4403 48960 4407
rect 48658 4373 48792 4403
rect 47992 4369 48792 4373
rect 48826 4373 48960 4403
rect 48994 4403 55174 4407
rect 48994 4373 49134 4403
rect 48826 4369 49134 4373
rect 49168 4369 55083 4403
rect 46394 4365 55083 4369
rect 40125 4356 55083 4365
rect 40022 4355 55083 4356
rect 39891 4351 55083 4355
rect 55135 4356 55174 4403
rect 55226 4356 55326 4408
rect 55135 4351 55326 4356
rect 39891 4346 55326 4351
rect 32997 4294 33100 4313
rect 32997 4291 33087 4294
rect 9734 4252 25100 4267
rect 9734 4200 9775 4252
rect 9827 4200 9871 4252
rect 9923 4251 25100 4252
rect 9923 4249 16386 4251
rect 9923 4242 16050 4249
rect 9923 4208 15882 4242
rect 15916 4215 16050 4242
rect 16084 4239 16386 4249
rect 16084 4215 16218 4239
rect 15916 4208 16218 4215
rect 9923 4205 16218 4208
rect 16252 4217 16386 4239
rect 16420 4249 16718 4251
rect 16420 4217 16552 4249
rect 16252 4215 16552 4217
rect 16586 4217 16718 4249
rect 16752 4217 16886 4251
rect 16920 4249 18148 4251
rect 16920 4217 17060 4249
rect 16586 4215 17060 4217
rect 17094 4247 18148 4249
rect 17094 4243 17978 4247
rect 17094 4215 17816 4243
rect 16252 4209 17816 4215
rect 17850 4213 17978 4243
rect 18012 4217 18148 4247
rect 18182 4250 25100 4251
rect 18182 4247 24985 4250
rect 18182 4217 18312 4247
rect 18012 4213 18312 4217
rect 18346 4213 18482 4247
rect 18516 4243 18818 4247
rect 18516 4213 18650 4243
rect 17850 4209 18650 4213
rect 18684 4213 18818 4243
rect 18852 4243 24985 4247
rect 18852 4213 18992 4243
rect 18684 4209 18992 4213
rect 19026 4209 24886 4243
rect 16252 4205 24886 4209
rect 9923 4200 24886 4205
rect 9734 4191 24886 4200
rect 24938 4198 24985 4243
rect 25037 4198 25100 4250
rect 33028 4242 33087 4291
rect 33028 4239 33100 4242
rect 32997 4217 33100 4239
rect 34537 4217 34572 4313
rect 46192 4306 48795 4312
rect 46192 4272 46224 4306
rect 46258 4272 46324 4306
rect 46358 4272 46424 4306
rect 46458 4272 46524 4306
rect 46558 4272 46624 4306
rect 46658 4272 46724 4306
rect 46758 4272 46824 4306
rect 46858 4272 46924 4306
rect 46958 4272 47884 4306
rect 47918 4272 47984 4306
rect 48018 4272 48084 4306
rect 48118 4272 48184 4306
rect 48218 4272 48284 4306
rect 48318 4272 48384 4306
rect 48418 4272 48484 4306
rect 48518 4272 48584 4306
rect 48618 4272 48795 4306
rect 46192 4267 48795 4272
rect 46192 4264 47638 4267
rect 47488 4263 47638 4264
rect 24938 4191 25100 4198
rect 9734 4186 25100 4191
rect 47488 4211 47533 4263
rect 47585 4215 47638 4263
rect 47690 4264 48795 4267
rect 47690 4215 47716 4264
rect 47585 4211 47716 4215
rect 47488 4172 47716 4211
rect 16050 4146 18653 4152
rect 16050 4112 16082 4146
rect 16116 4112 16182 4146
rect 16216 4112 16282 4146
rect 16316 4112 16382 4146
rect 16416 4112 16482 4146
rect 16516 4112 16582 4146
rect 16616 4112 16682 4146
rect 16716 4112 16782 4146
rect 16816 4112 17742 4146
rect 17776 4112 17842 4146
rect 17876 4112 17942 4146
rect 17976 4112 18042 4146
rect 18076 4112 18142 4146
rect 18176 4112 18242 4146
rect 18276 4112 18342 4146
rect 18376 4112 18442 4146
rect 18476 4112 18653 4146
rect 16050 4107 18653 4112
rect 16050 4104 17496 4107
rect 17346 4103 17496 4104
rect 17346 4051 17391 4103
rect 17443 4055 17496 4103
rect 17548 4104 18653 4107
rect 17548 4055 17574 4104
rect 17443 4051 17574 4055
rect 17346 4012 17574 4051
rect 47242 4020 47994 4078
rect 15712 3842 15763 3938
rect 17100 3866 17781 3924
rect 22231 3869 47742 3913
rect 22231 3867 47630 3869
rect 15712 3841 15762 3842
rect 22231 3815 33694 3867
rect 33746 3815 33838 3867
rect 33890 3815 33982 3867
rect 34034 3866 47630 3867
rect 34034 3815 47541 3866
rect 22231 3814 47541 3815
rect 47593 3817 47630 3866
rect 47682 3817 47742 3869
rect 47593 3814 47742 3817
rect 22231 3790 47742 3814
rect 22231 3783 47541 3790
rect 22231 3731 33693 3783
rect 33745 3731 33837 3783
rect 33889 3731 33981 3783
rect 34033 3738 47541 3783
rect 47593 3738 47634 3790
rect 47686 3738 47742 3790
rect 34033 3731 47742 3738
rect 17358 3707 47742 3731
rect 17358 3686 22437 3707
rect 17358 3634 17395 3686
rect 17447 3681 22437 3686
rect 17447 3634 17489 3681
rect 17358 3629 17489 3634
rect 17541 3629 22437 3681
rect 17358 3608 22437 3629
rect 17358 3606 17489 3608
rect 9525 3532 10188 3590
rect 17358 3554 17395 3606
rect 17447 3556 17489 3606
rect 17541 3556 22437 3608
rect 17447 3554 22437 3556
rect 17358 3525 22437 3554
rect 24623 3544 25251 3602
rect 39635 3544 40398 3602
rect 54825 3535 55476 3593
rect 62892 1474 63114 1552
<< via1 >>
rect 9774 5455 9826 5507
rect 9855 5454 9907 5506
rect 24890 5452 24942 5504
rect 24985 5452 25037 5504
rect 16953 5389 17005 5441
rect 17031 5389 17083 5441
rect 17124 5389 17176 5441
rect 32912 5412 32964 5464
rect 33025 5412 33077 5464
rect 33126 5412 33178 5464
rect 39967 5454 40019 5506
rect 40069 5454 40121 5506
rect 47104 5389 47156 5441
rect 47187 5389 47239 5441
rect 55085 5427 55137 5479
rect 55180 5427 55232 5479
rect 8782 5233 8834 5285
rect 8889 5235 8941 5287
rect 8991 5235 9043 5287
rect 9091 5236 9143 5288
rect 23812 5239 23864 5291
rect 23915 5239 23967 5291
rect 23998 5239 24050 5291
rect 24099 5239 24151 5291
rect 24186 5239 24238 5291
rect 38944 5235 38996 5287
rect 39032 5235 39084 5287
rect 39117 5240 39169 5292
rect 55860 5232 55912 5284
rect 55954 5232 56006 5284
rect 56031 5232 56083 5284
rect 56111 5231 56163 5283
rect 56185 5232 56237 5284
rect 32924 4789 32976 4841
rect 33027 4792 33079 4844
rect 33128 4792 33180 4844
rect 47110 4564 47162 4616
rect 47200 4565 47252 4617
rect 16977 4412 17029 4464
rect 17100 4412 17152 4464
rect 33705 4414 33757 4435
rect 33865 4420 33917 4435
rect 33705 4383 33724 4414
rect 33724 4383 33757 4414
rect 33865 4386 33892 4420
rect 33892 4386 33917 4420
rect 33865 4383 33917 4386
rect 33998 4383 34050 4435
rect 34111 4383 34163 4435
rect 39970 4355 40022 4407
rect 40073 4356 40125 4408
rect 55083 4351 55135 4403
rect 55174 4356 55226 4408
rect 9775 4200 9827 4252
rect 9871 4200 9923 4252
rect 24886 4191 24938 4243
rect 24985 4198 25037 4250
rect 32880 4237 32932 4289
rect 32976 4239 33028 4291
rect 33087 4242 33139 4294
rect 33179 4239 33231 4291
rect 47533 4211 47585 4263
rect 47638 4215 47690 4267
rect 17391 4051 17443 4103
rect 17496 4055 17548 4107
rect 48545 4024 48597 4076
rect 48637 4025 48689 4077
rect 48727 4024 48779 4076
rect 48815 4023 48867 4075
rect 16190 3863 16242 3915
rect 16274 3863 16326 3915
rect 16367 3864 16419 3916
rect 33694 3815 33746 3867
rect 33838 3815 33890 3867
rect 33982 3815 34034 3867
rect 47541 3814 47593 3866
rect 47630 3817 47682 3869
rect 33693 3731 33745 3783
rect 33837 3731 33889 3783
rect 33981 3731 34033 3783
rect 47541 3738 47593 3790
rect 47634 3738 47686 3790
rect 17395 3634 17447 3686
rect 17489 3629 17541 3681
rect 8776 3535 8828 3587
rect 8874 3535 8926 3587
rect 8969 3535 9021 3587
rect 9074 3535 9126 3587
rect 17395 3554 17447 3606
rect 17489 3556 17541 3608
rect 23826 3540 23878 3592
rect 23926 3540 23978 3592
rect 24025 3540 24077 3592
rect 24128 3540 24180 3592
rect 38934 3534 38986 3586
rect 39022 3534 39074 3586
rect 39120 3530 39172 3582
rect 55856 3531 55908 3583
rect 55944 3531 55996 3583
rect 56027 3531 56079 3583
rect 56114 3531 56166 3583
rect 9775 3317 9827 3369
rect 9855 3315 9907 3367
rect 24891 3332 24943 3384
rect 24974 3332 25026 3384
rect 39969 3322 40021 3374
rect 40060 3322 40112 3374
rect 55086 3307 55138 3359
rect 55169 3307 55221 3359
<< metal2 >>
rect 5788 7342 5832 8498
rect 7676 7342 7720 8498
rect 9564 7342 9608 8498
rect 11452 7342 11496 8498
rect 13340 7342 13384 8498
rect 15228 7342 15272 8498
rect 17116 7342 17160 8498
rect 19004 7342 19048 8498
rect 20892 7342 20936 8498
rect 22780 7342 22824 8498
rect 24668 7342 24712 8498
rect 26556 7342 26600 8498
rect 28444 7342 28488 8498
rect 30332 7342 30376 8498
rect 32220 7342 32264 8498
rect 34108 7342 34152 8498
rect 35996 7342 36040 8498
rect 37884 7342 37928 8498
rect 39772 7342 39816 8498
rect 41660 7342 41704 8498
rect 43548 7342 43592 8498
rect 45436 7342 45480 8498
rect 47324 7342 47368 8498
rect 49212 7342 49256 8498
rect 51100 7342 51144 8498
rect 52988 7342 53032 8498
rect 54876 7342 54920 8498
rect 56764 7342 56808 8498
rect 58652 7342 58696 8498
rect 60540 7342 60584 8498
rect 62428 7342 62472 8498
rect 0 7137 114 7141
rect 0 7101 4047 7137
rect 64807 7136 64921 7162
rect 0 1707 114 7101
rect 62457 7100 64921 7136
rect 427 6660 541 6695
rect 64449 6660 64563 6699
rect 427 6624 4040 6660
rect 62448 6624 64563 6660
rect 427 2204 541 6624
rect 9750 5507 9939 5537
rect 9750 5455 9774 5507
rect 9826 5506 9939 5507
rect 9826 5455 9855 5506
rect 9750 5454 9855 5455
rect 9907 5454 9939 5506
rect 8718 5288 9202 5413
rect 8718 5287 9091 5288
rect 8718 5285 8889 5287
rect 8718 5233 8782 5285
rect 8834 5235 8889 5285
rect 8941 5235 8991 5287
rect 9043 5236 9091 5287
rect 9143 5236 9202 5288
rect 9043 5235 9202 5236
rect 8834 5233 9202 5235
rect 8718 4066 9202 5233
rect 8718 4010 8785 4066
rect 8841 4010 8899 4066
rect 8955 4010 9013 4066
rect 9069 4010 9202 4066
rect 8718 3951 9202 4010
rect 8718 3895 8785 3951
rect 8841 3895 8899 3951
rect 8955 3895 9013 3951
rect 9069 3895 9202 3951
rect 8718 3836 9202 3895
rect 8718 3780 8785 3836
rect 8841 3780 8899 3836
rect 8955 3780 9013 3836
rect 9069 3780 9202 3836
rect 8718 3587 9202 3780
rect 8718 3535 8776 3587
rect 8828 3535 8874 3587
rect 8926 3535 8969 3587
rect 9021 3535 9074 3587
rect 9126 3535 9202 3587
rect 8718 3423 9202 3535
rect 9750 4252 9939 5454
rect 16933 5441 17193 5512
rect 16933 5389 16953 5441
rect 17005 5389 17031 5441
rect 17083 5389 17124 5441
rect 17176 5389 17193 5441
rect 24861 5504 25050 5527
rect 24861 5452 24890 5504
rect 24942 5452 24985 5504
rect 25037 5452 25050 5504
rect 16933 4464 17193 5389
rect 16933 4412 16977 4464
rect 17029 4412 17100 4464
rect 17152 4412 17193 4464
rect 16933 4368 17193 4412
rect 23774 5291 24241 5391
rect 23774 5239 23812 5291
rect 23864 5239 23915 5291
rect 23967 5239 23998 5291
rect 24050 5239 24099 5291
rect 24151 5239 24186 5291
rect 24238 5239 24241 5291
rect 9750 4200 9775 4252
rect 9827 4200 9871 4252
rect 9923 4200 9939 4252
rect 9750 3369 9939 4200
rect 17358 4107 17564 4152
rect 17358 4103 17496 4107
rect 17358 4051 17391 4103
rect 17443 4055 17496 4103
rect 17548 4055 17564 4107
rect 17443 4051 17564 4055
rect 9750 3317 9775 3369
rect 9827 3367 9939 3369
rect 9827 3317 9855 3367
rect 9750 3315 9855 3317
rect 9907 3315 9939 3367
rect 16139 3916 16492 3962
rect 16139 3915 16367 3916
rect 16139 3863 16190 3915
rect 16242 3863 16274 3915
rect 16326 3864 16367 3915
rect 16419 3864 16492 3916
rect 16326 3863 16492 3864
rect 16139 3505 16492 3863
rect 17358 3686 17564 4051
rect 17358 3634 17395 3686
rect 17447 3681 17564 3686
rect 17447 3634 17489 3681
rect 17358 3629 17489 3634
rect 17541 3629 17564 3681
rect 17358 3608 17564 3629
rect 17358 3606 17489 3608
rect 17358 3554 17395 3606
rect 17447 3556 17489 3606
rect 17541 3556 17564 3608
rect 17447 3554 17564 3556
rect 17358 3525 17564 3554
rect 23774 3976 24241 5239
rect 23774 3920 23824 3976
rect 23880 3920 23928 3976
rect 23984 3920 24032 3976
rect 24088 3920 24136 3976
rect 24192 3920 24241 3976
rect 23774 3860 24241 3920
rect 23774 3804 23824 3860
rect 23880 3804 23928 3860
rect 23984 3804 24032 3860
rect 24088 3804 24136 3860
rect 24192 3804 24241 3860
rect 23774 3744 24241 3804
rect 23774 3688 23824 3744
rect 23880 3688 23928 3744
rect 23984 3688 24032 3744
rect 24088 3688 24136 3744
rect 24192 3688 24241 3744
rect 23774 3592 24241 3688
rect 23774 3540 23826 3592
rect 23878 3540 23926 3592
rect 23978 3540 24025 3592
rect 24077 3540 24128 3592
rect 24180 3540 24241 3592
rect 16139 3449 16179 3505
rect 16235 3449 16287 3505
rect 16343 3449 16395 3505
rect 16451 3449 16492 3505
rect 16139 3411 16492 3449
rect 23774 3440 24241 3540
rect 24861 4250 25050 5452
rect 32866 5464 33201 5507
rect 32866 5412 32912 5464
rect 32964 5412 33025 5464
rect 33077 5412 33126 5464
rect 33178 5412 33201 5464
rect 32866 4844 33201 5412
rect 39952 5506 40139 5525
rect 39952 5454 39967 5506
rect 40019 5454 40069 5506
rect 40121 5454 40139 5506
rect 32866 4841 33027 4844
rect 32866 4789 32924 4841
rect 32976 4792 33027 4841
rect 33079 4792 33128 4844
rect 33180 4792 33201 4844
rect 32976 4789 33201 4792
rect 32866 4757 33201 4789
rect 38890 5292 39190 5389
rect 38890 5287 39117 5292
rect 38890 5235 38944 5287
rect 38996 5235 39032 5287
rect 39084 5240 39117 5287
rect 39169 5240 39190 5292
rect 39084 5235 39190 5240
rect 33637 4435 34176 4458
rect 33637 4383 33705 4435
rect 33757 4383 33865 4435
rect 33917 4383 33998 4435
rect 34050 4383 34111 4435
rect 34163 4383 34176 4435
rect 24861 4243 24985 4250
rect 24861 4191 24886 4243
rect 24938 4198 24985 4243
rect 25037 4198 25050 4250
rect 24938 4191 25050 4198
rect 16139 3355 16179 3411
rect 16235 3355 16287 3411
rect 16343 3355 16395 3411
rect 16451 3355 16492 3411
rect 16139 3329 16492 3355
rect 24861 3384 25050 4191
rect 32828 4294 33253 4312
rect 32828 4291 33087 4294
rect 32828 4289 32976 4291
rect 32828 4237 32880 4289
rect 32932 4239 32976 4289
rect 33028 4242 33087 4291
rect 33139 4291 33253 4294
rect 33139 4242 33179 4291
rect 33028 4239 33179 4242
rect 33231 4239 33253 4291
rect 32932 4237 33253 4239
rect 32828 3625 33253 4237
rect 33637 3867 34176 4383
rect 33637 3815 33694 3867
rect 33746 3815 33838 3867
rect 33890 3815 33982 3867
rect 34034 3815 34176 3867
rect 33637 3783 34176 3815
rect 33637 3731 33693 3783
rect 33745 3731 33837 3783
rect 33889 3731 33981 3783
rect 34033 3731 34176 3783
rect 33637 3657 34176 3731
rect 38890 4325 39190 5235
rect 38890 4269 38911 4325
rect 38967 4269 39005 4325
rect 39061 4269 39099 4325
rect 39155 4269 39190 4325
rect 38890 4237 39190 4269
rect 38890 4181 38911 4237
rect 38967 4181 39005 4237
rect 39061 4181 39099 4237
rect 39155 4181 39190 4237
rect 38890 4149 39190 4181
rect 38890 4093 38911 4149
rect 38967 4093 39005 4149
rect 39061 4093 39099 4149
rect 39155 4093 39190 4149
rect 32828 3569 32874 3625
rect 32930 3569 32999 3625
rect 33055 3569 33124 3625
rect 33180 3569 33253 3625
rect 32828 3529 33253 3569
rect 32828 3473 32874 3529
rect 32930 3473 32999 3529
rect 33055 3473 33124 3529
rect 33180 3473 33253 3529
rect 32828 3441 33253 3473
rect 38890 3586 39190 4093
rect 38890 3534 38934 3586
rect 38986 3534 39022 3586
rect 39074 3582 39190 3586
rect 39074 3534 39120 3582
rect 38890 3530 39120 3534
rect 39172 3530 39190 3582
rect 38890 3437 39190 3530
rect 39952 4408 40139 5454
rect 47081 5441 47300 5494
rect 47081 5389 47104 5441
rect 47156 5389 47187 5441
rect 47239 5389 47300 5441
rect 47081 4617 47300 5389
rect 47081 4616 47200 4617
rect 47081 4564 47110 4616
rect 47162 4565 47200 4616
rect 47252 4565 47300 4617
rect 47162 4564 47300 4565
rect 47081 4529 47300 4564
rect 55056 5479 55245 5502
rect 55056 5427 55085 5479
rect 55137 5427 55180 5479
rect 55232 5427 55245 5479
rect 39952 4407 40073 4408
rect 39952 4355 39970 4407
rect 40022 4356 40073 4407
rect 40125 4356 40139 4408
rect 40022 4355 40139 4356
rect 24861 3332 24891 3384
rect 24943 3332 24974 3384
rect 25026 3332 25050 3384
rect 24861 3319 25050 3332
rect 39952 3374 40139 4355
rect 55056 4408 55245 5427
rect 55056 4403 55174 4408
rect 55056 4351 55083 4403
rect 55135 4356 55174 4403
rect 55226 4356 55245 4408
rect 55135 4351 55245 4356
rect 47500 4267 47706 4312
rect 47500 4263 47638 4267
rect 47500 4211 47533 4263
rect 47585 4215 47638 4263
rect 47690 4215 47706 4267
rect 47585 4211 47706 4215
rect 47500 3869 47706 4211
rect 47500 3866 47630 3869
rect 47500 3814 47541 3866
rect 47593 3817 47630 3866
rect 47682 3817 47706 3869
rect 47593 3814 47706 3817
rect 47500 3790 47706 3814
rect 47500 3738 47541 3790
rect 47593 3738 47634 3790
rect 47686 3738 47706 3790
rect 47500 3695 47706 3738
rect 48508 4077 48922 4099
rect 48508 4076 48637 4077
rect 48508 4024 48545 4076
rect 48597 4025 48637 4076
rect 48689 4076 48922 4077
rect 48689 4025 48727 4076
rect 48597 4024 48727 4025
rect 48779 4075 48922 4076
rect 48779 4024 48815 4075
rect 48508 4023 48815 4024
rect 48867 4023 48922 4075
rect 39952 3322 39969 3374
rect 40021 3322 40060 3374
rect 40112 3322 40139 3374
rect 9750 3297 9939 3315
rect 39952 3314 40139 3322
rect 48508 3478 48922 4023
rect 48508 3422 48545 3478
rect 48601 3422 48638 3478
rect 48694 3422 48731 3478
rect 48787 3422 48824 3478
rect 48880 3422 48922 3478
rect 48508 3396 48922 3422
rect 48508 3340 48545 3396
rect 48601 3340 48638 3396
rect 48694 3340 48731 3396
rect 48787 3340 48824 3396
rect 48880 3340 48922 3396
rect 48508 3303 48922 3340
rect 55056 3359 55245 4351
rect 55821 5284 56242 5389
rect 55821 5232 55860 5284
rect 55912 5232 55954 5284
rect 56006 5232 56031 5284
rect 56083 5283 56185 5284
rect 56083 5232 56111 5283
rect 55821 5231 56111 5232
rect 56163 5232 56185 5283
rect 56237 5232 56242 5284
rect 56163 5231 56242 5232
rect 55821 3870 56242 5231
rect 55821 3814 55858 3870
rect 55914 3814 55962 3870
rect 56018 3814 56066 3870
rect 56122 3814 56170 3870
rect 56226 3814 56242 3870
rect 55821 3780 56242 3814
rect 55821 3724 55858 3780
rect 55914 3724 55962 3780
rect 56018 3724 56066 3780
rect 56122 3724 56170 3780
rect 56226 3724 56242 3780
rect 55821 3583 56242 3724
rect 55821 3531 55856 3583
rect 55908 3531 55944 3583
rect 55996 3531 56027 3583
rect 56079 3531 56114 3583
rect 56166 3531 56242 3583
rect 55821 3439 56242 3531
rect 55056 3307 55086 3359
rect 55138 3307 55169 3359
rect 55221 3307 55245 3359
rect 55056 3294 55245 3307
rect 1151 3058 2579 3248
rect 1151 2804 2037 3058
rect 1151 2718 2559 2804
rect 1151 2710 2037 2718
rect 64449 2204 64563 6624
rect 427 2168 822 2204
rect 1971 2168 2561 2204
rect 62797 2168 64563 2204
rect 427 2156 541 2168
rect 64449 2160 64563 2168
rect 64807 1722 64921 7100
rect 0 1671 734 1707
rect 62872 1686 64921 1722
rect 0 1665 114 1671
rect 64807 1665 64921 1686
rect 2530 1168 2574 1486
rect 4418 1168 4462 1486
rect 6306 1168 6350 1486
rect 8194 1168 8238 1486
rect 10082 1168 10126 1486
rect 11970 1168 12014 1486
rect 13858 1168 13902 1486
rect 15746 1168 15790 1486
rect 17634 1168 17678 1486
rect 19522 1168 19566 1486
rect 21410 1168 21454 1486
rect 23298 1168 23342 1486
rect 25186 1168 25230 1486
rect 27074 1168 27118 1486
rect 28962 1168 29006 1486
rect 30850 1168 30894 1486
rect 32738 1168 32782 1486
rect 34626 1168 34670 1486
rect 36514 1168 36558 1486
rect 38402 1168 38446 1486
rect 40290 1168 40334 1486
rect 42178 1168 42222 1486
rect 44066 1168 44110 1486
rect 45954 1168 45998 1486
rect 47842 1168 47886 1486
rect 49730 1168 49774 1486
rect 51618 1168 51662 1486
rect 53506 1168 53550 1486
rect 55394 1168 55438 1486
rect 57282 1168 57326 1486
rect 59170 1366 59214 1486
rect 59170 1168 59216 1366
rect 641 22 686 1168
rect 2529 22 2574 1168
rect 4417 22 4462 1168
rect 6305 22 6350 1168
rect 8193 22 8238 1168
rect 10081 22 10126 1168
rect 11969 22 12014 1168
rect 13857 22 13902 1168
rect 15745 22 15790 1168
rect 17633 22 17678 1168
rect 19521 22 19566 1168
rect 21409 22 21454 1168
rect 23297 22 23342 1168
rect 25185 22 25230 1168
rect 27073 22 27118 1168
rect 28961 22 29006 1168
rect 30849 22 30894 1168
rect 32737 22 32782 1168
rect 34625 22 34670 1168
rect 36513 22 36558 1168
rect 38401 22 38446 1168
rect 40289 22 40334 1168
rect 42177 22 42222 1168
rect 44065 22 44110 1168
rect 45953 22 45998 1168
rect 47841 22 47886 1168
rect 49729 22 49774 1168
rect 51617 22 51662 1168
rect 53505 22 53550 1168
rect 55393 22 55438 1168
rect 57281 22 57326 1168
rect 59169 468 59216 1168
rect 59169 22 59214 468
rect 61046 0 61102 1486
<< via2 >>
rect 8785 4010 8841 4066
rect 8899 4010 8955 4066
rect 9013 4010 9069 4066
rect 8785 3895 8841 3951
rect 8899 3895 8955 3951
rect 9013 3895 9069 3951
rect 8785 3780 8841 3836
rect 8899 3780 8955 3836
rect 9013 3780 9069 3836
rect 23824 3920 23880 3976
rect 23928 3920 23984 3976
rect 24032 3920 24088 3976
rect 24136 3920 24192 3976
rect 23824 3804 23880 3860
rect 23928 3804 23984 3860
rect 24032 3804 24088 3860
rect 24136 3804 24192 3860
rect 23824 3688 23880 3744
rect 23928 3688 23984 3744
rect 24032 3688 24088 3744
rect 24136 3688 24192 3744
rect 16179 3449 16235 3505
rect 16287 3449 16343 3505
rect 16395 3449 16451 3505
rect 16179 3355 16235 3411
rect 16287 3355 16343 3411
rect 16395 3355 16451 3411
rect 38911 4269 38967 4325
rect 39005 4269 39061 4325
rect 39099 4269 39155 4325
rect 38911 4181 38967 4237
rect 39005 4181 39061 4237
rect 39099 4181 39155 4237
rect 38911 4093 38967 4149
rect 39005 4093 39061 4149
rect 39099 4093 39155 4149
rect 32874 3569 32930 3625
rect 32999 3569 33055 3625
rect 33124 3569 33180 3625
rect 32874 3473 32930 3529
rect 32999 3473 33055 3529
rect 33124 3473 33180 3529
rect 48545 3422 48601 3478
rect 48638 3422 48694 3478
rect 48731 3422 48787 3478
rect 48824 3422 48880 3478
rect 48545 3340 48601 3396
rect 48638 3340 48694 3396
rect 48731 3340 48787 3396
rect 48824 3340 48880 3396
rect 55858 3814 55914 3870
rect 55962 3814 56018 3870
rect 56066 3814 56122 3870
rect 56170 3814 56226 3870
rect 55858 3724 55914 3780
rect 55962 3724 56018 3780
rect 56066 3724 56122 3780
rect 56170 3724 56226 3780
<< metal3 >>
rect 5028 8066 5134 8083
rect 5028 8002 5049 8066
rect 5113 8002 5134 8066
rect 5028 7986 5134 8002
rect 5028 7922 5049 7986
rect 5113 7922 5134 7986
rect 5028 7905 5134 7922
rect 5237 8065 5343 8082
rect 5237 8001 5258 8065
rect 5322 8001 5343 8065
rect 5237 7985 5343 8001
rect 5237 7921 5258 7985
rect 5322 7921 5343 7985
rect 5237 7904 5343 7921
rect 5403 8065 5509 8082
rect 5403 8001 5424 8065
rect 5488 8001 5509 8065
rect 5403 7985 5509 8001
rect 5403 7921 5424 7985
rect 5488 7921 5509 7985
rect 5403 7904 5509 7921
rect 5583 8067 5689 8084
rect 5583 8003 5604 8067
rect 5668 8003 5689 8067
rect 5583 7987 5689 8003
rect 5583 7923 5604 7987
rect 5668 7923 5689 7987
rect 5583 7906 5689 7923
rect 21657 8083 21763 8100
rect 21657 8019 21678 8083
rect 21742 8019 21763 8083
rect 21657 8003 21763 8019
rect 21657 7939 21678 8003
rect 21742 7939 21763 8003
rect 21657 7922 21763 7939
rect 21873 8083 21979 8100
rect 21873 8019 21894 8083
rect 21958 8019 21979 8083
rect 21873 8003 21979 8019
rect 21873 7939 21894 8003
rect 21958 7939 21979 8003
rect 21873 7922 21979 7939
rect 22089 8083 22195 8100
rect 22089 8019 22110 8083
rect 22174 8019 22195 8083
rect 22089 8003 22195 8019
rect 22089 7939 22110 8003
rect 22174 7939 22195 8003
rect 22089 7922 22195 7939
rect 30149 8082 30255 8099
rect 30149 8018 30170 8082
rect 30234 8018 30255 8082
rect 30149 8002 30255 8018
rect 30149 7938 30170 8002
rect 30234 7938 30255 8002
rect 30149 7921 30255 7938
rect 30365 8082 30471 8099
rect 30365 8018 30386 8082
rect 30450 8018 30471 8082
rect 30365 8002 30471 8018
rect 30365 7938 30386 8002
rect 30450 7938 30471 8002
rect 30365 7921 30471 7938
rect 30581 8082 30687 8099
rect 30581 8018 30602 8082
rect 30666 8018 30687 8082
rect 30581 8002 30687 8018
rect 30581 7938 30602 8002
rect 30666 7938 30687 8002
rect 30581 7921 30687 7938
rect 43677 8088 43783 8105
rect 43677 8024 43698 8088
rect 43762 8024 43783 8088
rect 43677 8008 43783 8024
rect 43677 7944 43698 8008
rect 43762 7944 43783 8008
rect 43677 7927 43783 7944
rect 43893 8088 43999 8105
rect 43893 8024 43914 8088
rect 43978 8024 43999 8088
rect 43893 8008 43999 8024
rect 43893 7944 43914 8008
rect 43978 7944 43999 8008
rect 43893 7927 43999 7944
rect 44109 8088 44215 8105
rect 44109 8024 44130 8088
rect 44194 8024 44215 8088
rect 44109 8008 44215 8024
rect 44109 7944 44130 8008
rect 44194 7944 44215 8008
rect 44109 7927 44215 7944
rect 60162 8081 60268 8098
rect 60162 8017 60183 8081
rect 60247 8017 60268 8081
rect 60162 8001 60268 8017
rect 60162 7937 60183 8001
rect 60247 7937 60268 8001
rect 60162 7920 60268 7937
rect 60378 8081 60484 8098
rect 60378 8017 60399 8081
rect 60463 8017 60484 8081
rect 60378 8001 60484 8017
rect 60378 7937 60399 8001
rect 60463 7937 60484 8001
rect 60378 7920 60484 7937
rect 60594 8081 60700 8098
rect 60594 8017 60615 8081
rect 60679 8017 60700 8081
rect 60594 8001 60700 8017
rect 60594 7937 60615 8001
rect 60679 7937 60700 8001
rect 60594 7920 60700 7937
rect 3682 5949 4577 6012
rect 3682 5948 3987 5949
rect 3682 5884 3815 5948
rect 3879 5885 3987 5948
rect 4051 5948 4577 5949
rect 4051 5885 4161 5948
rect 3879 5884 4161 5885
rect 4225 5884 4577 5948
rect 3682 5869 4577 5884
rect 3682 5868 3987 5869
rect 3682 5804 3815 5868
rect 3879 5805 3987 5868
rect 4051 5868 4577 5869
rect 4051 5805 4161 5868
rect 3879 5804 4161 5805
rect 4225 5804 4577 5868
rect 20122 5969 20228 5986
rect 20122 5905 20143 5969
rect 20207 5905 20228 5969
rect 20122 5889 20228 5905
rect 20122 5825 20143 5889
rect 20207 5825 20228 5889
rect 20122 5808 20228 5825
rect 20338 5969 20444 5986
rect 20338 5905 20359 5969
rect 20423 5905 20444 5969
rect 20338 5889 20444 5905
rect 20338 5825 20359 5889
rect 20423 5825 20444 5889
rect 20338 5808 20444 5825
rect 20554 5969 20660 5986
rect 20554 5905 20575 5969
rect 20639 5905 20660 5969
rect 20554 5889 20660 5905
rect 20554 5825 20575 5889
rect 20639 5825 20660 5889
rect 20554 5808 20660 5825
rect 28630 5961 28736 5978
rect 28630 5897 28651 5961
rect 28715 5897 28736 5961
rect 28630 5881 28736 5897
rect 28630 5817 28651 5881
rect 28715 5817 28736 5881
rect 3682 5758 4577 5804
rect 28630 5800 28736 5817
rect 28846 5961 28952 5978
rect 28846 5897 28867 5961
rect 28931 5897 28952 5961
rect 28846 5881 28952 5897
rect 28846 5817 28867 5881
rect 28931 5817 28952 5881
rect 28846 5800 28952 5817
rect 29062 5961 29168 5978
rect 29062 5897 29083 5961
rect 29147 5897 29168 5961
rect 29062 5881 29168 5897
rect 29062 5817 29083 5881
rect 29147 5817 29168 5881
rect 29062 5800 29168 5817
rect 42102 5956 42208 5973
rect 42102 5892 42123 5956
rect 42187 5892 42208 5956
rect 42102 5876 42208 5892
rect 42102 5812 42123 5876
rect 42187 5812 42208 5876
rect 42102 5795 42208 5812
rect 42318 5956 42424 5973
rect 42318 5892 42339 5956
rect 42403 5892 42424 5956
rect 42318 5876 42424 5892
rect 42318 5812 42339 5876
rect 42403 5812 42424 5876
rect 42318 5795 42424 5812
rect 42534 5956 42640 5973
rect 42534 5892 42555 5956
rect 42619 5892 42640 5956
rect 42534 5876 42640 5892
rect 42534 5812 42555 5876
rect 42619 5812 42640 5876
rect 42534 5795 42640 5812
rect 58653 5948 58759 5965
rect 58653 5884 58674 5948
rect 58738 5884 58759 5948
rect 58653 5868 58759 5884
rect 58653 5804 58674 5868
rect 58738 5804 58759 5868
rect 58653 5787 58759 5804
rect 58869 5948 58975 5965
rect 58869 5884 58890 5948
rect 58954 5884 58975 5948
rect 58869 5868 58975 5884
rect 58869 5804 58890 5868
rect 58954 5804 58975 5868
rect 58869 5787 58975 5804
rect 59085 5948 59191 5965
rect 59085 5884 59106 5948
rect 59170 5884 59191 5948
rect 59085 5868 59191 5884
rect 59085 5804 59106 5868
rect 59170 5804 59191 5868
rect 59085 5787 59191 5804
rect 38888 4325 39192 4339
rect 38888 4269 38911 4325
rect 38967 4269 39005 4325
rect 39061 4269 39099 4325
rect 39155 4269 39192 4325
rect 38888 4237 39192 4269
rect 38888 4181 38911 4237
rect 38967 4202 39005 4237
rect 38999 4181 39005 4202
rect 39061 4203 39099 4237
rect 39061 4181 39089 4203
rect 39155 4181 39192 4237
rect 38888 4149 38935 4181
rect 38999 4149 39089 4181
rect 39153 4149 39192 4181
rect 8784 4092 9126 4125
rect 38888 4093 38911 4149
rect 38999 4138 39005 4149
rect 38967 4093 39005 4138
rect 39061 4139 39089 4149
rect 39061 4093 39099 4139
rect 39155 4093 39192 4149
rect 8716 4066 9205 4092
rect 38888 4073 39192 4093
rect 8716 4010 8785 4066
rect 8841 4010 8899 4066
rect 8955 4010 9013 4066
rect 9069 4010 9205 4066
rect 8716 3951 9205 4010
rect 8716 3895 8785 3951
rect 8841 3909 8899 3951
rect 8955 3915 9013 3951
rect 8857 3895 8899 3909
rect 9008 3895 9013 3915
rect 9069 3915 9205 3951
rect 9069 3895 9089 3915
rect 8716 3845 8793 3895
rect 8857 3851 8944 3895
rect 9008 3851 9089 3895
rect 9153 3851 9205 3915
rect 8857 3845 9205 3851
rect 8716 3836 9205 3845
rect 8716 3780 8785 3836
rect 8841 3780 8899 3836
rect 8955 3780 9013 3836
rect 9069 3780 9205 3836
rect 8716 3725 9205 3780
rect 23774 3976 24241 4030
rect 23774 3920 23824 3976
rect 23880 3923 23928 3976
rect 23900 3920 23928 3923
rect 23984 3923 24032 3976
rect 23984 3920 24003 3923
rect 24088 3920 24136 3976
rect 24192 3920 24241 3976
rect 23774 3860 23836 3920
rect 23900 3860 24003 3920
rect 24067 3860 24241 3920
rect 23774 3804 23824 3860
rect 23900 3859 23928 3860
rect 23880 3804 23928 3859
rect 23984 3859 24003 3860
rect 23984 3804 24032 3859
rect 24088 3804 24136 3860
rect 24192 3804 24241 3860
rect 23774 3762 24241 3804
rect 23774 3744 23836 3762
rect 23900 3744 24003 3762
rect 24067 3744 24241 3762
rect 23774 3688 23824 3744
rect 23900 3698 23928 3744
rect 23880 3688 23928 3698
rect 23984 3698 24003 3744
rect 23984 3688 24032 3698
rect 24088 3688 24136 3744
rect 24192 3688 24241 3744
rect 55821 3870 56243 3898
rect 55821 3814 55858 3870
rect 55939 3814 55962 3870
rect 56060 3814 56066 3870
rect 56122 3814 56134 3870
rect 56226 3814 56243 3870
rect 55821 3806 55875 3814
rect 55939 3806 55996 3814
rect 56060 3806 56134 3814
rect 56198 3806 56243 3814
rect 55821 3790 56243 3806
rect 55821 3780 55875 3790
rect 55939 3780 55996 3790
rect 56060 3780 56134 3790
rect 56198 3780 56243 3790
rect 55821 3724 55858 3780
rect 55939 3726 55962 3780
rect 56060 3726 56066 3780
rect 55914 3724 55962 3726
rect 56018 3724 56066 3726
rect 56122 3726 56134 3780
rect 56122 3724 56170 3726
rect 56226 3724 56243 3780
rect 55821 3690 56243 3724
rect 23774 3644 24241 3688
rect 32826 3625 33251 3663
rect 32826 3569 32874 3625
rect 32930 3569 32999 3625
rect 33055 3569 33124 3625
rect 33180 3569 33251 3625
rect 32826 3562 33251 3569
rect 32826 3529 32883 3562
rect 32947 3529 33002 3562
rect 16139 3505 16492 3528
rect 16139 3454 16179 3505
rect 16235 3454 16287 3505
rect 16343 3454 16395 3505
rect 16139 3390 16169 3454
rect 16235 3449 16272 3454
rect 16343 3449 16375 3454
rect 16451 3449 16492 3505
rect 16233 3411 16272 3449
rect 16336 3411 16375 3449
rect 16439 3411 16492 3449
rect 32826 3473 32874 3529
rect 32947 3498 32999 3529
rect 33066 3498 33121 3562
rect 33185 3498 33251 3562
rect 32930 3473 32999 3498
rect 33055 3473 33124 3498
rect 33180 3473 33251 3498
rect 32826 3436 33251 3473
rect 48508 3495 48923 3545
rect 48508 3494 48696 3495
rect 48508 3478 48556 3494
rect 48620 3478 48696 3494
rect 48760 3478 48824 3495
rect 16235 3390 16272 3411
rect 16343 3390 16375 3411
rect 16139 3355 16179 3390
rect 16235 3355 16287 3390
rect 16343 3355 16395 3390
rect 16451 3355 16492 3411
rect 16139 3329 16492 3355
rect 48508 3422 48545 3478
rect 48620 3430 48638 3478
rect 48601 3422 48638 3430
rect 48694 3431 48696 3478
rect 48694 3422 48731 3431
rect 48787 3422 48824 3478
rect 48888 3431 48923 3495
rect 48880 3422 48923 3431
rect 48508 3415 48923 3422
rect 48508 3414 48696 3415
rect 48508 3396 48556 3414
rect 48620 3396 48696 3414
rect 48760 3396 48824 3415
rect 48508 3340 48545 3396
rect 48620 3350 48638 3396
rect 48601 3340 48638 3350
rect 48694 3351 48696 3396
rect 48694 3340 48731 3351
rect 48787 3340 48824 3396
rect 48888 3351 48923 3415
rect 48880 3340 48923 3351
rect 48508 3304 48923 3340
rect 3796 3000 3902 3017
rect 3796 2936 3817 3000
rect 3881 2936 3902 3000
rect 3796 2920 3902 2936
rect 3796 2856 3817 2920
rect 3881 2856 3902 2920
rect 3796 2839 3902 2856
rect 4001 3002 4107 3019
rect 4001 2938 4022 3002
rect 4086 2938 4107 3002
rect 4001 2922 4107 2938
rect 4001 2858 4022 2922
rect 4086 2858 4107 2922
rect 4001 2841 4107 2858
rect 4200 3002 4306 3019
rect 4200 2938 4221 3002
rect 4285 2938 4306 3002
rect 4200 2922 4306 2938
rect 4200 2858 4221 2922
rect 4285 2858 4306 2922
rect 4200 2841 4306 2858
rect 20113 3018 20219 3035
rect 20113 2954 20134 3018
rect 20198 2954 20219 3018
rect 20113 2938 20219 2954
rect 20113 2874 20134 2938
rect 20198 2874 20219 2938
rect 20113 2857 20219 2874
rect 20329 3018 20435 3035
rect 20329 2954 20350 3018
rect 20414 2954 20435 3018
rect 20329 2938 20435 2954
rect 20329 2874 20350 2938
rect 20414 2874 20435 2938
rect 20329 2857 20435 2874
rect 20545 3018 20651 3035
rect 20545 2954 20566 3018
rect 20630 2954 20651 3018
rect 20545 2938 20651 2954
rect 20545 2874 20566 2938
rect 20630 2874 20651 2938
rect 20545 2857 20651 2874
rect 28635 3013 28741 3030
rect 28635 2949 28656 3013
rect 28720 2949 28741 3013
rect 28635 2933 28741 2949
rect 28635 2869 28656 2933
rect 28720 2869 28741 2933
rect 28635 2852 28741 2869
rect 28851 3013 28957 3030
rect 28851 2949 28872 3013
rect 28936 2949 28957 3013
rect 28851 2933 28957 2949
rect 28851 2869 28872 2933
rect 28936 2869 28957 2933
rect 28851 2852 28957 2869
rect 29067 3013 29173 3030
rect 29067 2949 29088 3013
rect 29152 2949 29173 3013
rect 29067 2933 29173 2949
rect 29067 2869 29088 2933
rect 29152 2869 29173 2933
rect 29067 2852 29173 2869
rect 42138 3015 42244 3032
rect 42138 2951 42159 3015
rect 42223 2951 42244 3015
rect 42138 2935 42244 2951
rect 42138 2871 42159 2935
rect 42223 2871 42244 2935
rect 42138 2854 42244 2871
rect 42354 3015 42460 3032
rect 42354 2951 42375 3015
rect 42439 2951 42460 3015
rect 42354 2935 42460 2951
rect 42354 2871 42375 2935
rect 42439 2871 42460 2935
rect 42354 2854 42460 2871
rect 42570 3015 42676 3032
rect 42570 2951 42591 3015
rect 42655 2951 42676 3015
rect 42570 2935 42676 2951
rect 42570 2871 42591 2935
rect 42655 2871 42676 2935
rect 42570 2854 42676 2871
rect 58633 3026 58739 3043
rect 58633 2962 58654 3026
rect 58718 2962 58739 3026
rect 58633 2946 58739 2962
rect 58633 2882 58654 2946
rect 58718 2882 58739 2946
rect 58633 2865 58739 2882
rect 58849 3026 58955 3043
rect 58849 2962 58870 3026
rect 58934 2962 58955 3026
rect 58849 2946 58955 2962
rect 58849 2882 58870 2946
rect 58934 2882 58955 2946
rect 58849 2865 58955 2882
rect 59065 3026 59171 3043
rect 59065 2962 59086 3026
rect 59150 2962 59171 3026
rect 59065 2946 59171 2962
rect 59065 2882 59086 2946
rect 59150 2882 59171 2946
rect 59065 2865 59171 2882
rect 5042 889 5148 906
rect 5042 825 5063 889
rect 5127 825 5148 889
rect 5042 809 5148 825
rect 5042 745 5063 809
rect 5127 745 5148 809
rect 5042 728 5148 745
rect 5263 889 5369 906
rect 5263 825 5284 889
rect 5348 825 5369 889
rect 5263 809 5369 825
rect 5263 745 5284 809
rect 5348 745 5369 809
rect 5263 728 5369 745
rect 5472 889 5578 906
rect 5472 825 5493 889
rect 5557 825 5578 889
rect 5472 809 5578 825
rect 5472 745 5493 809
rect 5557 745 5578 809
rect 5472 728 5578 745
rect 5646 889 5752 906
rect 5646 825 5667 889
rect 5731 825 5752 889
rect 16289 900 16366 903
rect 5646 809 5752 825
rect 5646 745 5667 809
rect 5731 745 5752 809
rect 8770 837 8856 851
rect 8770 773 8781 837
rect 8845 773 8856 837
rect 8770 760 8856 773
rect 8918 837 9004 851
rect 8918 773 8929 837
rect 8993 773 9004 837
rect 8918 760 9004 773
rect 9066 837 9152 851
rect 9066 773 9077 837
rect 9141 773 9152 837
rect 16289 836 16295 900
rect 16359 836 16366 900
rect 16289 834 16366 836
rect 21675 888 21781 905
rect 21675 824 21696 888
rect 21760 824 21781 888
rect 21675 808 21781 824
rect 9066 760 9152 773
rect 16312 781 16389 784
rect 5646 728 5752 745
rect 16312 717 16318 781
rect 16382 717 16389 781
rect 21675 744 21696 808
rect 21760 744 21781 808
rect 21675 727 21781 744
rect 21891 888 21997 905
rect 21891 824 21912 888
rect 21976 824 21997 888
rect 21891 808 21997 824
rect 21891 744 21912 808
rect 21976 744 21997 808
rect 21891 727 21997 744
rect 22107 888 22213 905
rect 22107 824 22128 888
rect 22192 824 22213 888
rect 30104 893 30210 910
rect 22107 808 22213 824
rect 22107 744 22128 808
rect 22192 744 22213 808
rect 23827 841 23923 863
rect 23827 777 23843 841
rect 23907 777 23923 841
rect 23827 755 23923 777
rect 23960 841 24056 863
rect 23960 777 23976 841
rect 24040 777 24056 841
rect 23960 755 24056 777
rect 24093 841 24189 863
rect 24093 777 24109 841
rect 24173 777 24189 841
rect 24093 755 24189 777
rect 30104 829 30125 893
rect 30189 829 30210 893
rect 30104 813 30210 829
rect 22107 727 22213 744
rect 30104 749 30125 813
rect 30189 749 30210 813
rect 30104 732 30210 749
rect 30320 893 30426 910
rect 30320 829 30341 893
rect 30405 829 30426 893
rect 30320 813 30426 829
rect 30320 749 30341 813
rect 30405 749 30426 813
rect 30320 732 30426 749
rect 30536 893 30642 910
rect 30536 829 30557 893
rect 30621 829 30642 893
rect 43622 883 43728 900
rect 30536 813 30642 829
rect 30536 749 30557 813
rect 30621 749 30642 813
rect 30536 732 30642 749
rect 32893 830 32980 854
rect 32893 766 32904 830
rect 32968 766 32980 830
rect 32893 742 32980 766
rect 33016 830 33103 854
rect 33016 766 33027 830
rect 33091 766 33103 830
rect 33016 742 33103 766
rect 33148 830 33235 854
rect 33148 766 33159 830
rect 33223 766 33235 830
rect 33148 742 33235 766
rect 38922 827 39009 851
rect 38922 763 38933 827
rect 38997 763 39009 827
rect 38922 739 39009 763
rect 39091 827 39178 851
rect 39091 763 39102 827
rect 39166 763 39178 827
rect 39091 739 39178 763
rect 43622 819 43643 883
rect 43707 819 43728 883
rect 43622 803 43728 819
rect 43622 739 43643 803
rect 43707 739 43728 803
rect 43622 722 43728 739
rect 43838 883 43944 900
rect 43838 819 43859 883
rect 43923 819 43944 883
rect 43838 803 43944 819
rect 43838 739 43859 803
rect 43923 739 43944 803
rect 43838 722 43944 739
rect 44054 883 44160 900
rect 55871 887 55955 894
rect 44054 819 44075 883
rect 44139 819 44160 883
rect 44054 803 44160 819
rect 44054 739 44075 803
rect 44139 739 44160 803
rect 44054 722 44160 739
rect 48548 877 48632 884
rect 48548 813 48558 877
rect 48622 813 48632 877
rect 48548 797 48632 813
rect 48548 733 48558 797
rect 48622 733 48632 797
rect 48548 726 48632 733
rect 48661 877 48745 884
rect 48661 813 48671 877
rect 48735 813 48745 877
rect 48661 797 48745 813
rect 48661 733 48671 797
rect 48735 733 48745 797
rect 48661 726 48745 733
rect 48776 877 48860 884
rect 48776 813 48786 877
rect 48850 813 48860 877
rect 48776 797 48860 813
rect 48776 733 48786 797
rect 48850 733 48860 797
rect 55871 823 55881 887
rect 55945 823 55955 887
rect 55871 807 55955 823
rect 55871 743 55881 807
rect 55945 743 55955 807
rect 55871 736 55955 743
rect 55990 887 56074 894
rect 55990 823 56000 887
rect 56064 823 56074 887
rect 55990 807 56074 823
rect 55990 743 56000 807
rect 56064 743 56074 807
rect 55990 736 56074 743
rect 56119 887 56203 894
rect 56119 823 56129 887
rect 56193 823 56203 887
rect 56119 807 56203 823
rect 56119 743 56129 807
rect 56193 743 56203 807
rect 56119 736 56203 743
rect 60134 878 60240 895
rect 60134 814 60155 878
rect 60219 814 60240 878
rect 60134 798 60240 814
rect 48776 726 48860 733
rect 60134 734 60155 798
rect 60219 734 60240 798
rect 60134 717 60240 734
rect 60350 878 60456 895
rect 60350 814 60371 878
rect 60435 814 60456 878
rect 60350 798 60456 814
rect 60350 734 60371 798
rect 60435 734 60456 798
rect 60350 717 60456 734
rect 60566 878 60672 895
rect 60566 814 60587 878
rect 60651 814 60672 878
rect 60566 798 60672 814
rect 60566 734 60587 798
rect 60651 734 60672 798
rect 60566 717 60672 734
rect 16312 715 16389 717
<< via3 >>
rect 5049 8002 5113 8066
rect 5049 7922 5113 7986
rect 5258 8001 5322 8065
rect 5258 7921 5322 7985
rect 5424 8001 5488 8065
rect 5424 7921 5488 7985
rect 5604 8003 5668 8067
rect 5604 7923 5668 7987
rect 21678 8019 21742 8083
rect 21678 7939 21742 8003
rect 21894 8019 21958 8083
rect 21894 7939 21958 8003
rect 22110 8019 22174 8083
rect 22110 7939 22174 8003
rect 30170 8018 30234 8082
rect 30170 7938 30234 8002
rect 30386 8018 30450 8082
rect 30386 7938 30450 8002
rect 30602 8018 30666 8082
rect 30602 7938 30666 8002
rect 43698 8024 43762 8088
rect 43698 7944 43762 8008
rect 43914 8024 43978 8088
rect 43914 7944 43978 8008
rect 44130 8024 44194 8088
rect 44130 7944 44194 8008
rect 60183 8017 60247 8081
rect 60183 7937 60247 8001
rect 60399 8017 60463 8081
rect 60399 7937 60463 8001
rect 60615 8017 60679 8081
rect 60615 7937 60679 8001
rect 3815 5884 3879 5948
rect 3987 5885 4051 5949
rect 4161 5884 4225 5948
rect 3815 5804 3879 5868
rect 3987 5805 4051 5869
rect 4161 5804 4225 5868
rect 20143 5905 20207 5969
rect 20143 5825 20207 5889
rect 20359 5905 20423 5969
rect 20359 5825 20423 5889
rect 20575 5905 20639 5969
rect 20575 5825 20639 5889
rect 28651 5897 28715 5961
rect 28651 5817 28715 5881
rect 28867 5897 28931 5961
rect 28867 5817 28931 5881
rect 29083 5897 29147 5961
rect 29083 5817 29147 5881
rect 42123 5892 42187 5956
rect 42123 5812 42187 5876
rect 42339 5892 42403 5956
rect 42339 5812 42403 5876
rect 42555 5892 42619 5956
rect 42555 5812 42619 5876
rect 58674 5884 58738 5948
rect 58674 5804 58738 5868
rect 58890 5884 58954 5948
rect 58890 5804 58954 5868
rect 59106 5884 59170 5948
rect 59106 5804 59170 5868
rect 38935 4181 38967 4202
rect 38967 4181 38999 4202
rect 39089 4181 39099 4203
rect 39099 4181 39153 4203
rect 38935 4149 38999 4181
rect 39089 4149 39153 4181
rect 38935 4138 38967 4149
rect 38967 4138 38999 4149
rect 39089 4139 39099 4149
rect 39099 4139 39153 4149
rect 8793 3895 8841 3909
rect 8841 3895 8857 3909
rect 8944 3895 8955 3915
rect 8955 3895 9008 3915
rect 8793 3845 8857 3895
rect 8944 3851 9008 3895
rect 9089 3851 9153 3915
rect 23836 3920 23880 3923
rect 23880 3920 23900 3923
rect 24003 3920 24032 3923
rect 24032 3920 24067 3923
rect 23836 3860 23900 3920
rect 24003 3860 24067 3920
rect 23836 3859 23880 3860
rect 23880 3859 23900 3860
rect 24003 3859 24032 3860
rect 24032 3859 24067 3860
rect 23836 3744 23900 3762
rect 24003 3744 24067 3762
rect 23836 3698 23880 3744
rect 23880 3698 23900 3744
rect 24003 3698 24032 3744
rect 24032 3698 24067 3744
rect 55875 3814 55914 3870
rect 55914 3814 55939 3870
rect 55996 3814 56018 3870
rect 56018 3814 56060 3870
rect 56134 3814 56170 3870
rect 56170 3814 56198 3870
rect 55875 3806 55939 3814
rect 55996 3806 56060 3814
rect 56134 3806 56198 3814
rect 55875 3780 55939 3790
rect 55996 3780 56060 3790
rect 56134 3780 56198 3790
rect 55875 3726 55914 3780
rect 55914 3726 55939 3780
rect 55996 3726 56018 3780
rect 56018 3726 56060 3780
rect 56134 3726 56170 3780
rect 56170 3726 56198 3780
rect 32883 3529 32947 3562
rect 33002 3529 33066 3562
rect 16169 3449 16179 3454
rect 16179 3449 16233 3454
rect 16272 3449 16287 3454
rect 16287 3449 16336 3454
rect 16375 3449 16395 3454
rect 16395 3449 16439 3454
rect 16169 3411 16233 3449
rect 16272 3411 16336 3449
rect 16375 3411 16439 3449
rect 32883 3498 32930 3529
rect 32930 3498 32947 3529
rect 33002 3498 33055 3529
rect 33055 3498 33066 3529
rect 33121 3529 33185 3562
rect 33121 3498 33124 3529
rect 33124 3498 33180 3529
rect 33180 3498 33185 3529
rect 48556 3478 48620 3494
rect 48696 3478 48760 3495
rect 48824 3478 48888 3495
rect 16169 3390 16179 3411
rect 16179 3390 16233 3411
rect 16272 3390 16287 3411
rect 16287 3390 16336 3411
rect 16375 3390 16395 3411
rect 16395 3390 16439 3411
rect 48556 3430 48601 3478
rect 48601 3430 48620 3478
rect 48696 3431 48731 3478
rect 48731 3431 48760 3478
rect 48824 3431 48880 3478
rect 48880 3431 48888 3478
rect 48556 3396 48620 3414
rect 48696 3396 48760 3415
rect 48824 3396 48888 3415
rect 48556 3350 48601 3396
rect 48601 3350 48620 3396
rect 48696 3351 48731 3396
rect 48731 3351 48760 3396
rect 48824 3351 48880 3396
rect 48880 3351 48888 3396
rect 3817 2936 3881 3000
rect 3817 2856 3881 2920
rect 4022 2938 4086 3002
rect 4022 2858 4086 2922
rect 4221 2938 4285 3002
rect 4221 2858 4285 2922
rect 20134 2954 20198 3018
rect 20134 2874 20198 2938
rect 20350 2954 20414 3018
rect 20350 2874 20414 2938
rect 20566 2954 20630 3018
rect 20566 2874 20630 2938
rect 28656 2949 28720 3013
rect 28656 2869 28720 2933
rect 28872 2949 28936 3013
rect 28872 2869 28936 2933
rect 29088 2949 29152 3013
rect 29088 2869 29152 2933
rect 42159 2951 42223 3015
rect 42159 2871 42223 2935
rect 42375 2951 42439 3015
rect 42375 2871 42439 2935
rect 42591 2951 42655 3015
rect 42591 2871 42655 2935
rect 58654 2962 58718 3026
rect 58654 2882 58718 2946
rect 58870 2962 58934 3026
rect 58870 2882 58934 2946
rect 59086 2962 59150 3026
rect 59086 2882 59150 2946
rect 5063 825 5127 889
rect 5063 745 5127 809
rect 5284 825 5348 889
rect 5284 745 5348 809
rect 5493 825 5557 889
rect 5493 745 5557 809
rect 5667 825 5731 889
rect 5667 745 5731 809
rect 8781 773 8845 837
rect 8929 773 8993 837
rect 9077 773 9141 837
rect 16295 836 16359 900
rect 21696 824 21760 888
rect 16318 717 16382 781
rect 21696 744 21760 808
rect 21912 824 21976 888
rect 21912 744 21976 808
rect 22128 824 22192 888
rect 22128 744 22192 808
rect 23843 777 23907 841
rect 23976 777 24040 841
rect 24109 777 24173 841
rect 30125 829 30189 893
rect 30125 749 30189 813
rect 30341 829 30405 893
rect 30341 749 30405 813
rect 30557 829 30621 893
rect 30557 749 30621 813
rect 32904 766 32968 830
rect 33027 766 33091 830
rect 33159 766 33223 830
rect 38933 763 38997 827
rect 39102 763 39166 827
rect 43643 819 43707 883
rect 43643 739 43707 803
rect 43859 819 43923 883
rect 43859 739 43923 803
rect 44075 819 44139 883
rect 44075 739 44139 803
rect 48558 813 48622 877
rect 48558 733 48622 797
rect 48671 813 48735 877
rect 48671 733 48735 797
rect 48786 813 48850 877
rect 48786 733 48850 797
rect 55881 823 55945 887
rect 55881 743 55945 807
rect 56000 823 56064 887
rect 56000 743 56064 807
rect 56129 823 56193 887
rect 56129 743 56193 807
rect 60155 814 60219 878
rect 60155 734 60219 798
rect 60371 814 60435 878
rect 60371 734 60435 798
rect 60587 814 60651 878
rect 60587 734 60651 798
<< metal4 >>
rect 3650 5949 4456 8265
rect 3650 5948 3987 5949
rect 3650 5884 3815 5948
rect 3879 5885 3987 5948
rect 4051 5948 4456 5949
rect 4051 5885 4161 5948
rect 3879 5884 4161 5885
rect 4225 5884 4456 5948
rect 3650 5869 4456 5884
rect 3650 5868 3987 5869
rect 3650 5804 3815 5868
rect 3879 5805 3987 5868
rect 4051 5868 4456 5869
rect 4051 5805 4161 5868
rect 3879 5804 4161 5805
rect 4225 5804 4456 5868
rect 3650 3002 4456 5804
rect 3650 3000 4022 3002
rect 3650 2936 3817 3000
rect 3881 2938 4022 3000
rect 4086 2938 4221 3002
rect 4285 2938 4456 3002
rect 3881 2936 4456 2938
rect 3650 2922 4456 2936
rect 3650 2920 4022 2922
rect 3650 2856 3817 2920
rect 3881 2858 4022 2920
rect 4086 2858 4221 2922
rect 4285 2858 4456 2922
rect 3881 2856 4456 2858
rect 3650 559 4456 2856
rect 4993 8067 5799 8266
rect 4993 8066 5604 8067
rect 4993 8002 5049 8066
rect 5113 8065 5604 8066
rect 5113 8002 5258 8065
rect 4993 8001 5258 8002
rect 5322 8001 5424 8065
rect 5488 8003 5604 8065
rect 5668 8003 5799 8067
rect 5488 8001 5799 8003
rect 4993 7987 5799 8001
rect 4993 7986 5604 7987
rect 4993 7922 5049 7986
rect 5113 7985 5604 7986
rect 5113 7922 5258 7985
rect 4993 7921 5258 7922
rect 5322 7921 5424 7985
rect 5488 7923 5604 7985
rect 5668 7923 5799 7987
rect 5488 7921 5799 7923
rect 4993 889 5799 7921
rect 19993 5969 20799 8266
rect 19993 5905 20143 5969
rect 20207 5905 20359 5969
rect 20423 5905 20575 5969
rect 20639 5905 20799 5969
rect 19993 5889 20799 5905
rect 19993 5825 20143 5889
rect 20207 5825 20359 5889
rect 20423 5825 20575 5889
rect 20639 5825 20799 5889
rect 4993 825 5063 889
rect 5127 825 5284 889
rect 5348 825 5493 889
rect 5557 825 5667 889
rect 5731 825 5799 889
rect 4993 809 5799 825
rect 4993 745 5063 809
rect 5127 745 5284 809
rect 5348 745 5493 809
rect 5557 745 5667 809
rect 5731 745 5799 809
rect 4993 560 5799 745
rect 8724 3915 9193 4044
rect 8724 3909 8944 3915
rect 8724 3845 8793 3909
rect 8857 3851 8944 3909
rect 9008 3851 9089 3915
rect 9153 3851 9193 3915
rect 8857 3845 9193 3851
rect 8724 837 9193 3845
rect 16139 3454 16493 3529
rect 16139 3390 16169 3454
rect 16233 3390 16272 3454
rect 16336 3390 16375 3454
rect 16439 3390 16493 3454
rect 16139 3328 16493 3390
rect 8724 773 8781 837
rect 8845 773 8929 837
rect 8993 773 9077 837
rect 9141 773 9193 837
rect 8724 661 9193 773
rect 16215 900 16416 3328
rect 16215 836 16295 900
rect 16359 836 16416 900
rect 16215 781 16416 836
rect 16215 717 16318 781
rect 16382 717 16416 781
rect 16215 636 16416 717
rect 19993 3018 20799 5825
rect 19993 2954 20134 3018
rect 20198 2954 20350 3018
rect 20414 2954 20566 3018
rect 20630 2954 20799 3018
rect 19993 2938 20799 2954
rect 19993 2874 20134 2938
rect 20198 2874 20350 2938
rect 20414 2874 20566 2938
rect 20630 2874 20799 2938
rect 19993 560 20799 2874
rect 21493 8083 22299 8266
rect 21493 8019 21678 8083
rect 21742 8019 21894 8083
rect 21958 8019 22110 8083
rect 22174 8019 22299 8083
rect 21493 8003 22299 8019
rect 21493 7939 21678 8003
rect 21742 7939 21894 8003
rect 21958 7939 22110 8003
rect 22174 7939 22299 8003
rect 21493 888 22299 7939
rect 28493 5961 29299 8266
rect 28493 5897 28651 5961
rect 28715 5897 28867 5961
rect 28931 5897 29083 5961
rect 29147 5897 29299 5961
rect 28493 5881 29299 5897
rect 28493 5817 28651 5881
rect 28715 5817 28867 5881
rect 28931 5817 29083 5881
rect 29147 5817 29299 5881
rect 21493 824 21696 888
rect 21760 824 21912 888
rect 21976 824 22128 888
rect 22192 824 22299 888
rect 21493 808 22299 824
rect 21493 744 21696 808
rect 21760 744 21912 808
rect 21976 744 22128 808
rect 22192 744 22299 808
rect 21493 560 22299 744
rect 23774 3923 24241 4058
rect 23774 3859 23836 3923
rect 23900 3859 24003 3923
rect 24067 3859 24241 3923
rect 23774 3762 24241 3859
rect 23774 3698 23836 3762
rect 23900 3698 24003 3762
rect 24067 3698 24241 3762
rect 23774 841 24241 3698
rect 23774 777 23843 841
rect 23907 777 23976 841
rect 24040 777 24109 841
rect 24173 777 24241 841
rect 23774 686 24241 777
rect 28493 3013 29299 5817
rect 28493 2949 28656 3013
rect 28720 2949 28872 3013
rect 28936 2949 29088 3013
rect 29152 2949 29299 3013
rect 28493 2933 29299 2949
rect 28493 2869 28656 2933
rect 28720 2869 28872 2933
rect 28936 2869 29088 2933
rect 29152 2869 29299 2933
rect 28493 560 29299 2869
rect 29993 8082 30799 8266
rect 29993 8018 30170 8082
rect 30234 8018 30386 8082
rect 30450 8018 30602 8082
rect 30666 8018 30799 8082
rect 29993 8002 30799 8018
rect 29993 7938 30170 8002
rect 30234 7938 30386 8002
rect 30450 7938 30602 8002
rect 30666 7938 30799 8002
rect 29993 893 30799 7938
rect 41993 5956 42799 8266
rect 41993 5892 42123 5956
rect 42187 5892 42339 5956
rect 42403 5892 42555 5956
rect 42619 5892 42799 5956
rect 41993 5876 42799 5892
rect 41993 5812 42123 5876
rect 42187 5812 42339 5876
rect 42403 5812 42555 5876
rect 42619 5812 42799 5876
rect 38888 4203 39193 4384
rect 38888 4202 39089 4203
rect 38888 4138 38935 4202
rect 38999 4139 39089 4202
rect 39153 4139 39193 4203
rect 38999 4138 39193 4139
rect 29993 829 30125 893
rect 30189 829 30341 893
rect 30405 829 30557 893
rect 30621 829 30799 893
rect 29993 813 30799 829
rect 29993 749 30125 813
rect 30189 749 30341 813
rect 30405 749 30557 813
rect 30621 749 30799 813
rect 29993 560 30799 749
rect 32826 3562 33251 3665
rect 32826 3498 32883 3562
rect 32947 3498 33002 3562
rect 33066 3498 33121 3562
rect 33185 3498 33251 3562
rect 32826 830 33251 3498
rect 32826 766 32904 830
rect 32968 766 33027 830
rect 33091 766 33159 830
rect 33223 766 33251 830
rect 32826 700 33251 766
rect 38888 827 39193 4138
rect 38888 763 38933 827
rect 38997 763 39102 827
rect 39166 763 39193 827
rect 38888 691 39193 763
rect 41993 3015 42799 5812
rect 41993 2951 42159 3015
rect 42223 2951 42375 3015
rect 42439 2951 42591 3015
rect 42655 2951 42799 3015
rect 41993 2935 42799 2951
rect 41993 2871 42159 2935
rect 42223 2871 42375 2935
rect 42439 2871 42591 2935
rect 42655 2871 42799 2935
rect 41993 560 42799 2871
rect 43493 8088 44299 8266
rect 43493 8024 43698 8088
rect 43762 8024 43914 8088
rect 43978 8024 44130 8088
rect 44194 8024 44299 8088
rect 43493 8008 44299 8024
rect 43493 7944 43698 8008
rect 43762 7944 43914 8008
rect 43978 7944 44130 8008
rect 44194 7944 44299 8008
rect 43493 883 44299 7944
rect 58493 5948 59299 8266
rect 58493 5884 58674 5948
rect 58738 5884 58890 5948
rect 58954 5884 59106 5948
rect 59170 5884 59299 5948
rect 58493 5868 59299 5884
rect 58493 5804 58674 5868
rect 58738 5804 58890 5868
rect 58954 5804 59106 5868
rect 59170 5804 59299 5868
rect 55821 3870 56246 3900
rect 55821 3806 55875 3870
rect 55939 3806 55996 3870
rect 56060 3806 56134 3870
rect 56198 3806 56246 3870
rect 55821 3790 56246 3806
rect 55821 3726 55875 3790
rect 55939 3726 55996 3790
rect 56060 3726 56134 3790
rect 56198 3726 56246 3790
rect 43493 819 43643 883
rect 43707 819 43859 883
rect 43923 819 44075 883
rect 44139 819 44299 883
rect 43493 803 44299 819
rect 43493 739 43643 803
rect 43707 739 43859 803
rect 43923 739 44075 803
rect 44139 739 44299 803
rect 43493 560 44299 739
rect 48508 3495 48922 3591
rect 48508 3494 48696 3495
rect 48508 3430 48556 3494
rect 48620 3431 48696 3494
rect 48760 3431 48824 3495
rect 48888 3431 48922 3495
rect 48620 3430 48922 3431
rect 48508 3415 48922 3430
rect 48508 3414 48696 3415
rect 48508 3350 48556 3414
rect 48620 3351 48696 3414
rect 48760 3351 48824 3415
rect 48888 3351 48922 3415
rect 48620 3350 48922 3351
rect 48508 877 48922 3350
rect 48508 813 48558 877
rect 48622 813 48671 877
rect 48735 813 48786 877
rect 48850 813 48922 877
rect 48508 797 48922 813
rect 48508 733 48558 797
rect 48622 733 48671 797
rect 48735 733 48786 797
rect 48850 733 48922 797
rect 48508 638 48922 733
rect 55821 887 56246 3726
rect 55821 823 55881 887
rect 55945 823 56000 887
rect 56064 823 56129 887
rect 56193 823 56246 887
rect 55821 807 56246 823
rect 55821 743 55881 807
rect 55945 743 56000 807
rect 56064 743 56129 807
rect 56193 743 56246 807
rect 55821 650 56246 743
rect 58493 3026 59299 5804
rect 58493 2962 58654 3026
rect 58718 2962 58870 3026
rect 58934 2962 59086 3026
rect 59150 2962 59299 3026
rect 58493 2946 59299 2962
rect 58493 2882 58654 2946
rect 58718 2882 58870 2946
rect 58934 2882 59086 2946
rect 59150 2882 59299 2946
rect 58493 560 59299 2882
rect 59993 8081 60799 8266
rect 59993 8017 60183 8081
rect 60247 8017 60399 8081
rect 60463 8017 60615 8081
rect 60679 8017 60799 8081
rect 59993 8001 60799 8017
rect 59993 7937 60183 8001
rect 60247 7937 60399 8001
rect 60463 7937 60615 8001
rect 60679 7937 60799 8001
rect 59993 878 60799 7937
rect 59993 814 60155 878
rect 60219 814 60371 878
rect 60435 814 60587 878
rect 60651 814 60799 878
rect 59993 798 60799 814
rect 59993 734 60155 798
rect 60219 734 60371 798
rect 60435 734 60587 798
rect 60651 734 60799 798
rect 59993 560 60799 734
use nbrhalf  nbrhalf_0
timestamp 1656715967
transform -1 0 58940 0 -1 10662
box -3552 2527 26658 5446
use nbrhalf  nbrhalf_1
timestamp 1656715967
transform 1 0 36264 0 1 -1834
box -3552 2527 26658 5446
use nbrhalf  nbrhalf_2
timestamp 1656715967
transform 1 0 6062 0 1 -1834
box -3552 2527 26658 5446
use nbrhalf_64  nbrhalf_64_0
timestamp 1656715967
transform -1 0 28738 0 -1 10662
box -3552 2527 26308 5446
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0
timestamp 1656715967
transform 1 0 32537 0 1 4265
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0
timestamp 1656715967
transform 1 0 33085 0 1 4265
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1656715967
transform 1 0 47821 0 1 4049
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_2
timestamp 1656715967
transform 1 0 45891 0 1 4049
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_3
timestamp 1656715967
transform 1 0 17679 0 1 3889
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_4
timestamp 1656715967
transform 1 0 15749 0 1 3889
box -38 -48 1510 592
use unitcell_nbr  unitcell_nbr_0
timestamp 1656715967
transform 1 0 1196 0 1 1878
box -574 -1185 1322 1192
<< labels >>
flabel metal1 s 62892 1474 63114 1552 1 FreeSans 2000 0 0 0 OUT
port 1 nsew
flabel metal4 s 3650 559 4456 8265 1 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal4 s 19993 560 20799 8266 1 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal4 s 28493 560 29299 8266 1 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal4 s 41993 560 42799 8266 1 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal4 s 58493 560 59299 8266 1 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal4 s 4993 560 5799 8266 1 FreeSans 2000 0 0 0 VSS
port 3 nsew
flabel metal4 s 21493 560 22299 8266 1 FreeSans 2000 0 0 0 VSS
port 3 nsew
flabel metal4 s 29993 560 30799 8266 1 FreeSans 2000 0 0 0 VSS
port 3 nsew
flabel metal4 s 43493 560 44299 8266 1 FreeSans 2000 0 0 0 VSS
port 3 nsew
flabel metal4 s 59993 560 60799 8266 1 FreeSans 2000 0 0 0 VSS
port 3 nsew
flabel metal1 s 219 4626 753 4690 1 FreeSans 2000 0 0 0 RESET
port 4 nsew
flabel metal2 s 62428 7342 62472 8498 1 FreeSans 2000 0 0 0 C[0]
port 5 nsew
flabel metal2 s 60540 7342 60584 8498 1 FreeSans 2000 0 0 0 C[1]
port 6 nsew
flabel metal2 s 58652 7342 58696 8498 1 FreeSans 2000 0 0 0 C[2]
port 7 nsew
flabel metal2 s 56764 7342 56808 8498 1 FreeSans 2000 0 0 0 C[3]
port 8 nsew
flabel metal2 s 54876 7342 54920 8498 1 FreeSans 2000 0 0 0 C[4]
port 9 nsew
flabel metal2 s 52988 7342 53032 8498 1 FreeSans 2000 0 0 0 C[5]
port 10 nsew
flabel metal2 s 51100 7342 51144 8498 1 FreeSans 2000 0 0 0 C[6]
port 11 nsew
flabel metal2 s 49212 7342 49256 8498 1 FreeSans 2000 0 0 0 C[7]
port 12 nsew
flabel metal2 s 47324 7342 47368 8498 1 FreeSans 2000 0 0 0 C[8]
port 13 nsew
flabel metal2 s 45436 7342 45480 8498 1 FreeSans 2000 0 0 0 C[9]
port 14 nsew
flabel metal2 s 43548 7342 43592 8498 1 FreeSans 2000 0 0 0 C[10]
port 15 nsew
flabel metal2 s 41660 7342 41704 8498 1 FreeSans 2000 0 0 0 C[11]
port 16 nsew
flabel metal2 s 39772 7342 39816 8498 1 FreeSans 2000 0 0 0 C[12]
port 17 nsew
flabel metal2 s 37884 7342 37928 8498 1 FreeSans 2000 0 0 0 C[13]
port 18 nsew
flabel metal2 s 35996 7342 36040 8498 1 FreeSans 2000 0 0 0 C[14]
port 19 nsew
flabel metal2 s 34108 7342 34152 8498 1 FreeSans 2000 0 0 0 C[15]
port 20 nsew
flabel metal2 s 32220 7342 32264 8498 1 FreeSans 2000 0 0 0 C[16]
port 21 nsew
flabel metal2 s 30332 7342 30376 8498 1 FreeSans 2000 0 0 0 C[17]
port 22 nsew
flabel metal2 s 28444 7342 28488 8498 1 FreeSans 2000 0 0 0 C[18]
port 23 nsew
flabel metal2 s 26556 7342 26600 8498 1 FreeSans 2000 0 0 0 C[19]
port 24 nsew
flabel metal2 s 24668 7342 24712 8498 1 FreeSans 2000 0 0 0 C[20]
port 25 nsew
flabel metal2 s 22780 7342 22824 8498 1 FreeSans 2000 0 0 0 C[21]
port 26 nsew
flabel metal2 s 20892 7342 20936 8498 1 FreeSans 2000 0 0 0 C[22]
port 27 nsew
flabel metal2 s 19004 7342 19048 8498 1 FreeSans 2000 0 0 0 C[23]
port 28 nsew
flabel metal2 s 17116 7342 17160 8498 1 FreeSans 2000 0 0 0 C[24]
port 29 nsew
flabel metal2 s 15228 7342 15272 8498 1 FreeSans 2000 0 0 0 C[25]
port 30 nsew
flabel metal2 s 13340 7342 13384 8498 1 FreeSans 2000 0 0 0 C[26]
port 31 nsew
flabel metal2 s 11452 7342 11496 8498 1 FreeSans 2000 0 0 0 C[27]
port 32 nsew
flabel metal2 s 9564 7342 9608 8498 1 FreeSans 2000 0 0 0 C[28]
port 33 nsew
flabel metal2 s 7676 7342 7720 8498 1 FreeSans 2000 0 0 0 C[29]
port 34 nsew
flabel metal2 s 5788 7342 5832 8498 1 FreeSans 2000 0 0 0 C[30]
port 35 nsew
flabel metal2 s 641 22 686 1168 1 FreeSans 2000 0 0 0 C[31]
port 36 nsew
flabel metal2 s 2529 22 2574 1168 1 FreeSans 2000 0 0 0 C[32]
port 37 nsew
flabel metal2 s 4417 22 4462 1168 1 FreeSans 2000 0 0 0 C[33]
port 38 nsew
flabel metal2 s 6305 22 6350 1168 1 FreeSans 2000 0 0 0 C[34]
port 39 nsew
flabel metal2 s 8193 22 8238 1168 1 FreeSans 2000 0 0 0 C[35]
port 40 nsew
flabel metal2 s 10081 22 10126 1168 1 FreeSans 2000 0 0 0 C[36]
port 41 nsew
flabel metal2 s 11969 22 12014 1168 1 FreeSans 2000 0 0 0 C[37]
port 42 nsew
flabel metal2 s 13857 22 13902 1168 1 FreeSans 2000 0 0 0 C[38]
port 43 nsew
flabel metal2 s 15745 22 15790 1168 1 FreeSans 2000 0 0 0 C[39]
port 44 nsew
flabel metal2 s 17633 22 17678 1168 1 FreeSans 2000 0 0 0 C[40]
port 45 nsew
flabel metal2 s 19521 22 19566 1168 1 FreeSans 2000 0 0 0 C[41]
port 46 nsew
flabel metal2 s 21409 22 21454 1168 1 FreeSans 2000 0 0 0 C[42]
port 47 nsew
flabel metal2 s 23297 22 23342 1168 1 FreeSans 2000 0 0 0 C[43]
port 48 nsew
flabel metal2 s 25185 22 25230 1168 1 FreeSans 2000 0 0 0 C[44]
port 49 nsew
flabel metal2 s 27073 22 27118 1168 1 FreeSans 2000 0 0 0 C[45]
port 50 nsew
flabel metal2 s 28961 22 29006 1168 1 FreeSans 2000 0 0 0 C[46]
port 51 nsew
flabel metal2 s 30849 22 30894 1168 1 FreeSans 2000 0 0 0 C[47]
port 52 nsew
flabel metal2 s 32737 22 32782 1168 1 FreeSans 2000 0 0 0 C[48]
port 53 nsew
flabel metal2 s 34625 22 34670 1168 1 FreeSans 2000 0 0 0 C[49]
port 54 nsew
flabel metal2 s 36513 22 36558 1168 1 FreeSans 2000 0 0 0 C[50]
port 55 nsew
flabel metal2 s 38401 22 38446 1168 1 FreeSans 2000 0 0 0 C[51]
port 56 nsew
flabel metal2 s 40289 22 40334 1168 1 FreeSans 2000 0 0 0 C[52]
port 57 nsew
flabel metal2 s 42177 22 42222 1168 1 FreeSans 2000 0 0 0 C[53]
port 58 nsew
flabel metal2 s 44065 22 44110 1168 1 FreeSans 2000 0 0 0 C[54]
port 59 nsew
flabel metal2 s 45953 22 45998 1168 1 FreeSans 2000 0 0 0 C[55]
port 60 nsew
flabel metal2 s 47841 22 47886 1168 1 FreeSans 2000 0 0 0 C[56]
port 61 nsew
flabel metal2 s 49729 22 49774 1168 1 FreeSans 2000 0 0 0 C[57]
port 62 nsew
flabel metal2 s 51617 22 51662 1168 1 FreeSans 2000 0 0 0 C[58]
port 63 nsew
flabel metal2 s 53505 22 53550 1168 1 FreeSans 2000 0 0 0 C[59]
port 64 nsew
flabel metal2 s 55393 22 55438 1168 1 FreeSans 2000 0 0 0 C[60]
port 65 nsew
flabel metal2 s 57281 22 57326 1168 1 FreeSans 2000 0 0 0 C[61]
port 66 nsew
flabel metal2 s 59169 22 59214 1168 1 FreeSans 2000 0 0 0 C[62]
port 67 nsew
flabel metal2 s 61046 0 61102 1486 1 FreeSans 2000 0 0 0 C[63]
port 68 nsew
<< properties >>
string GDS_END 9171932
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/design_merged.gds
string GDS_START 9106060
<< end >>
