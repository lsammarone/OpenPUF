magic
tech sky130A
magscale 1 2
timestamp 1656715967
<< error_p >>
rect -38 261 866 582
rect 60 47 112 177
rect 142 47 196 177
rect 226 47 280 177
rect 310 47 364 177
rect 394 47 448 177
rect 478 47 532 177
rect 562 47 616 177
rect 646 47 700 177
rect 730 47 782 177
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 34 21 808 203
rect 34 17 63 21
rect 29 -17 63 17
<< scnmos >>
rect 112 47 142 177
rect 196 47 226 177
rect 280 47 310 177
rect 364 47 394 177
rect 448 47 478 177
rect 532 47 562 177
rect 616 47 646 177
rect 700 47 730 177
<< scpmoshvt >>
rect 112 297 142 497
rect 196 297 226 497
rect 280 297 310 497
rect 364 297 394 497
rect 448 297 478 497
rect 532 297 562 497
rect 616 297 646 497
rect 700 297 730 497
<< ndiff >>
rect 60 93 112 177
rect 60 59 68 93
rect 102 59 112 93
rect 60 47 112 59
rect 142 161 196 177
rect 142 127 152 161
rect 186 127 196 161
rect 142 93 196 127
rect 142 59 152 93
rect 186 59 196 93
rect 142 47 196 59
rect 226 93 280 177
rect 226 59 236 93
rect 270 59 280 93
rect 226 47 280 59
rect 310 161 364 177
rect 310 127 320 161
rect 354 127 364 161
rect 310 93 364 127
rect 310 59 320 93
rect 354 59 364 93
rect 310 47 364 59
rect 394 93 448 177
rect 394 59 404 93
rect 438 59 448 93
rect 394 47 448 59
rect 478 161 532 177
rect 478 127 488 161
rect 522 127 532 161
rect 478 93 532 127
rect 478 59 488 93
rect 522 59 532 93
rect 478 47 532 59
rect 562 93 616 177
rect 562 59 572 93
rect 606 59 616 93
rect 562 47 616 59
rect 646 161 700 177
rect 646 127 656 161
rect 690 127 700 161
rect 646 93 700 127
rect 646 59 656 93
rect 690 59 700 93
rect 646 47 700 59
rect 730 93 782 177
rect 730 59 740 93
rect 774 59 782 93
rect 730 47 782 59
<< pdiff >>
rect 60 485 112 497
rect 60 451 68 485
rect 102 451 112 485
rect 60 417 112 451
rect 60 383 68 417
rect 102 383 112 417
rect 60 297 112 383
rect 142 485 196 497
rect 142 451 152 485
rect 186 451 196 485
rect 142 417 196 451
rect 142 383 152 417
rect 186 383 196 417
rect 142 349 196 383
rect 142 315 152 349
rect 186 315 196 349
rect 142 297 196 315
rect 226 485 280 497
rect 226 451 236 485
rect 270 451 280 485
rect 226 417 280 451
rect 226 383 236 417
rect 270 383 280 417
rect 226 297 280 383
rect 310 485 364 497
rect 310 451 320 485
rect 354 451 364 485
rect 310 417 364 451
rect 310 383 320 417
rect 354 383 364 417
rect 310 349 364 383
rect 310 315 320 349
rect 354 315 364 349
rect 310 297 364 315
rect 394 485 448 497
rect 394 451 404 485
rect 438 451 448 485
rect 394 417 448 451
rect 394 383 404 417
rect 438 383 448 417
rect 394 297 448 383
rect 478 485 532 497
rect 478 451 488 485
rect 522 451 532 485
rect 478 417 532 451
rect 478 383 488 417
rect 522 383 532 417
rect 478 349 532 383
rect 478 315 488 349
rect 522 315 532 349
rect 478 297 532 315
rect 562 485 616 497
rect 562 451 572 485
rect 606 451 616 485
rect 562 417 616 451
rect 562 383 572 417
rect 606 383 616 417
rect 562 297 616 383
rect 646 485 700 497
rect 646 451 656 485
rect 690 451 700 485
rect 646 417 700 451
rect 646 383 656 417
rect 690 383 700 417
rect 646 349 700 383
rect 646 315 656 349
rect 690 315 700 349
rect 646 297 700 315
rect 730 485 782 497
rect 730 451 740 485
rect 774 451 782 485
rect 730 417 782 451
rect 730 383 740 417
rect 774 383 782 417
rect 730 297 782 383
<< ndiffc >>
rect 68 59 102 93
rect 152 127 186 161
rect 152 59 186 93
rect 236 59 270 93
rect 320 127 354 161
rect 320 59 354 93
rect 404 59 438 93
rect 488 127 522 161
rect 488 59 522 93
rect 572 59 606 93
rect 656 127 690 161
rect 656 59 690 93
rect 740 59 774 93
<< pdiffc >>
rect 68 451 102 485
rect 68 383 102 417
rect 152 451 186 485
rect 152 383 186 417
rect 152 315 186 349
rect 236 451 270 485
rect 236 383 270 417
rect 320 451 354 485
rect 320 383 354 417
rect 320 315 354 349
rect 404 451 438 485
rect 404 383 438 417
rect 488 451 522 485
rect 488 383 522 417
rect 488 315 522 349
rect 572 451 606 485
rect 572 383 606 417
rect 656 451 690 485
rect 656 383 690 417
rect 656 315 690 349
rect 740 451 774 485
rect 740 383 774 417
<< poly >>
rect 112 497 142 523
rect 196 497 226 523
rect 280 497 310 523
rect 364 497 394 523
rect 448 497 478 523
rect 532 497 562 523
rect 616 497 646 523
rect 700 497 730 523
rect 112 265 142 297
rect 196 265 226 297
rect 280 265 310 297
rect 364 265 394 297
rect 448 265 478 297
rect 532 265 562 297
rect 616 265 646 297
rect 700 265 730 297
rect 112 249 730 265
rect 112 215 152 249
rect 186 215 236 249
rect 270 215 320 249
rect 354 215 404 249
rect 438 215 488 249
rect 522 215 572 249
rect 606 215 656 249
rect 690 215 730 249
rect 112 199 730 215
rect 112 177 142 199
rect 196 177 226 199
rect 280 177 310 199
rect 364 177 394 199
rect 448 177 478 199
rect 532 177 562 199
rect 616 177 646 199
rect 700 177 730 199
rect 112 21 142 47
rect 196 21 226 47
rect 280 21 310 47
rect 364 21 394 47
rect 448 21 478 47
rect 532 21 562 47
rect 616 21 646 47
rect 700 21 730 47
<< polycont >>
rect 152 215 186 249
rect 236 215 270 249
rect 320 215 354 249
rect 404 215 438 249
rect 488 215 522 249
rect 572 215 606 249
rect 656 215 690 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 51 485 102 527
rect 51 451 68 485
rect 51 417 102 451
rect 51 383 68 417
rect 51 367 102 383
rect 136 485 202 493
rect 136 451 152 485
rect 186 451 202 485
rect 136 417 202 451
rect 136 383 152 417
rect 186 383 202 417
rect 136 349 202 383
rect 236 485 270 527
rect 236 417 270 451
rect 236 367 270 383
rect 304 485 370 493
rect 304 451 320 485
rect 354 451 370 485
rect 304 417 370 451
rect 304 383 320 417
rect 354 383 370 417
rect 136 333 152 349
rect 17 315 152 333
rect 186 333 202 349
rect 304 349 370 383
rect 404 485 438 527
rect 404 417 438 451
rect 404 367 438 383
rect 472 485 538 493
rect 472 451 488 485
rect 522 451 538 485
rect 472 417 538 451
rect 472 383 488 417
rect 522 383 538 417
rect 304 333 320 349
rect 186 315 320 333
rect 354 333 370 349
rect 472 349 538 383
rect 572 485 606 527
rect 572 417 606 451
rect 572 367 606 383
rect 640 485 706 493
rect 640 451 656 485
rect 690 451 706 485
rect 640 417 706 451
rect 640 383 656 417
rect 690 383 706 417
rect 472 333 488 349
rect 354 315 488 333
rect 522 333 538 349
rect 640 349 706 383
rect 740 485 800 527
rect 774 451 800 485
rect 740 417 800 451
rect 774 383 800 417
rect 740 367 800 383
rect 640 333 656 349
rect 522 315 656 333
rect 690 333 706 349
rect 690 315 811 333
rect 17 299 811 315
rect 17 181 86 299
rect 136 249 707 265
rect 136 215 152 249
rect 186 215 236 249
rect 270 215 320 249
rect 354 215 404 249
rect 438 215 488 249
rect 522 215 572 249
rect 606 215 656 249
rect 690 215 707 249
rect 747 181 811 299
rect 17 161 811 181
rect 17 143 152 161
rect 136 127 152 143
rect 186 143 320 161
rect 186 127 202 143
rect 51 93 102 109
rect 51 59 68 93
rect 51 17 102 59
rect 136 93 202 127
rect 304 127 320 143
rect 354 143 488 161
rect 354 127 370 143
rect 136 59 152 93
rect 186 59 202 93
rect 136 51 202 59
rect 236 93 270 109
rect 236 17 270 59
rect 304 93 370 127
rect 472 127 488 143
rect 522 143 656 161
rect 522 127 538 143
rect 304 59 320 93
rect 354 59 370 93
rect 304 51 370 59
rect 404 93 438 109
rect 404 17 438 59
rect 472 93 538 127
rect 640 127 656 143
rect 690 143 811 161
rect 690 127 706 143
rect 472 59 488 93
rect 522 59 538 93
rect 472 51 538 59
rect 572 93 606 109
rect 572 17 606 59
rect 640 93 706 127
rect 640 59 656 93
rect 690 59 706 93
rect 640 51 706 59
rect 740 93 801 109
rect 774 59 801 93
rect 740 17 801 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 213 221 247 255 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 305 221 339 255 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 397 221 431 255 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 489 221 523 255 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 581 221 615 255 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 673 221 707 255 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 765 221 799 255 0 FreeSans 487 0 0 0 Y
port 2 nsew
flabel locali s 29 221 63 255 0 FreeSans 487 0 0 0 Y
port 2 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 390 0 0 0 VNB
port 3 nsew
flabel nwell s 29 527 63 561 0 FreeSans 390 0 0 0 VPB
port 4 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 390 0 0 0 VGND
port 5 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 390 0 0 0 VPWR
port 6 nsew
flabel locali s 230 238 230 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 322 238 322 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 414 238 414 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 506 238 506 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 598 238 598 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 690 238 690 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 782 238 782 238 0 FreeSans 487 0 0 0 Y
port 2 nsew
flabel locali s 46 238 46 238 0 FreeSans 487 0 0 0 Y
port 2 nsew
flabel pwell s 46 0 46 0 0 FreeSans 390 0 0 0 VNB
port 3 nsew
flabel nwell s 46 544 46 544 0 FreeSans 390 0 0 0 VPB
port 4 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 390 0 0 0 VGND
port 5 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 390 0 0 0 VPWR
port 6 nsew
flabel locali s 230 238 230 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 322 238 322 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 414 238 414 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 506 238 506 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 598 238 598 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 690 238 690 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 782 238 782 238 0 FreeSans 487 0 0 0 Y
port 2 nsew
flabel locali s 46 238 46 238 0 FreeSans 487 0 0 0 Y
port 2 nsew
flabel pwell s 46 0 46 0 0 FreeSans 390 0 0 0 VNB
port 3 nsew
flabel nwell s 46 544 46 544 0 FreeSans 390 0 0 0 VPB
port 4 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 390 0 0 0 VGND
port 5 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 390 0 0 0 VPWR
port 6 nsew
flabel locali s 230 238 230 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 322 238 322 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 414 238 414 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 506 238 506 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 598 238 598 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 690 238 690 238 0 FreeSans 487 0 0 0 A
port 1 nsew
flabel locali s 782 238 782 238 0 FreeSans 487 0 0 0 Y
port 2 nsew
flabel locali s 46 238 46 238 0 FreeSans 487 0 0 0 Y
port 2 nsew
flabel pwell s 46 0 46 0 0 FreeSans 390 0 0 0 VNB
port 3 nsew
flabel nwell s 46 544 46 544 0 FreeSans 390 0 0 0 VPB
port 4 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 390 0 0 0 VGND
port 5 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 390 0 0 0 VPWR
port 6 nsew
flabel locali s 230 238 230 238 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel locali s 322 238 322 238 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel locali s 414 238 414 238 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel locali s 506 238 506 238 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel locali s 598 238 598 238 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel locali s 690 238 690 238 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel locali s 782 238 782 238 0 FreeSans 250 0 0 0 Y
port 2 nsew
flabel locali s 46 238 46 238 0 FreeSans 250 0 0 0 Y
port 2 nsew
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
rlabel comment s 0 0 0 0 4 inv_8
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 9627510
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/design_merged.gds
string GDS_START 9585002
string path 0.000 0.000 20.700 0.000 
<< end >>
