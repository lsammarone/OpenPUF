magic
tech sky130A
magscale 1 2
timestamp 1656715967
<< nwell >>
rect 14749 3456 15131 3777
rect 44891 3616 45273 3937
<< nsubdiff >>
rect 45016 3789 45150 3808
rect 45016 3755 45088 3789
rect 45122 3755 45150 3789
rect 45016 3738 45150 3755
rect 14874 3629 15008 3648
rect 14874 3595 14946 3629
rect 14980 3595 15008 3629
rect 14874 3578 15008 3595
<< nsubdiffcont >>
rect 45088 3755 45122 3789
rect 14946 3595 14980 3629
<< locali >>
rect 44813 3789 45356 3809
rect 44813 3755 45088 3789
rect 45122 3755 45356 3789
rect 44813 3737 45356 3755
rect 43682 3715 43716 3721
rect 43514 3708 43548 3714
rect 44018 3717 44052 3723
rect 43682 3676 43716 3681
rect 43850 3705 43884 3711
rect 43514 3669 43548 3674
rect 44018 3678 44052 3683
rect 44184 3715 44218 3721
rect 44184 3676 44218 3681
rect 44350 3717 44384 3723
rect 44350 3678 44384 3683
rect 44518 3717 44552 3723
rect 44518 3678 44552 3683
rect 44692 3715 44726 3721
rect 44692 3676 44726 3681
rect 45448 3709 45482 3715
rect 43850 3666 43884 3671
rect 45448 3670 45482 3675
rect 45610 3713 45644 3719
rect 45610 3674 45644 3679
rect 45780 3717 45814 3723
rect 45780 3678 45814 3683
rect 45944 3713 45978 3719
rect 45944 3674 45978 3679
rect 46114 3713 46148 3719
rect 46114 3674 46148 3679
rect 46282 3709 46316 3715
rect 46282 3670 46316 3675
rect 46450 3713 46484 3719
rect 46450 3674 46484 3679
rect 46624 3709 46658 3715
rect 46624 3670 46658 3675
rect 14671 3629 15214 3649
rect 14671 3595 14946 3629
rect 14980 3595 15214 3629
rect 14671 3577 15214 3595
rect 13540 3555 13574 3561
rect 13372 3548 13406 3554
rect 13876 3557 13910 3563
rect 13540 3516 13574 3521
rect 13708 3545 13742 3551
rect 13372 3509 13406 3514
rect 13876 3518 13910 3523
rect 14042 3555 14076 3561
rect 14042 3516 14076 3521
rect 14208 3557 14242 3563
rect 14208 3518 14242 3523
rect 14376 3557 14410 3563
rect 14376 3518 14410 3523
rect 14550 3555 14584 3561
rect 14550 3516 14584 3521
rect 15306 3549 15340 3555
rect 13708 3506 13742 3511
rect 15306 3510 15340 3515
rect 15468 3553 15502 3559
rect 15468 3514 15502 3519
rect 15638 3557 15672 3563
rect 15638 3518 15672 3523
rect 15802 3553 15836 3559
rect 15802 3514 15836 3519
rect 15972 3553 16006 3559
rect 15972 3514 16006 3519
rect 16140 3549 16174 3555
rect 16140 3510 16174 3515
rect 16308 3553 16342 3559
rect 16308 3514 16342 3519
rect 16482 3549 16516 3555
rect 16482 3510 16516 3515
<< viali >>
rect 43514 3674 43548 3708
rect 43682 3681 43716 3715
rect 43850 3671 43884 3705
rect 44018 3683 44052 3717
rect 44184 3681 44218 3715
rect 44350 3683 44384 3717
rect 44518 3683 44552 3717
rect 44692 3681 44726 3715
rect 45448 3675 45482 3709
rect 45610 3679 45644 3713
rect 45780 3683 45814 3717
rect 45944 3679 45978 3713
rect 46114 3679 46148 3713
rect 46282 3675 46316 3709
rect 46450 3679 46484 3713
rect 46624 3675 46658 3709
rect 43714 3578 43748 3612
rect 43814 3578 43848 3612
rect 43914 3578 43948 3612
rect 44014 3578 44048 3612
rect 44114 3578 44148 3612
rect 44214 3578 44248 3612
rect 44314 3578 44348 3612
rect 44414 3578 44448 3612
rect 45374 3578 45408 3612
rect 45474 3578 45508 3612
rect 45574 3578 45608 3612
rect 45674 3578 45708 3612
rect 45774 3578 45808 3612
rect 45874 3578 45908 3612
rect 45974 3578 46008 3612
rect 46074 3578 46108 3612
rect 13372 3514 13406 3548
rect 13540 3521 13574 3555
rect 13708 3511 13742 3545
rect 13876 3523 13910 3557
rect 14042 3521 14076 3555
rect 14208 3523 14242 3557
rect 14376 3523 14410 3557
rect 14550 3521 14584 3555
rect 15306 3515 15340 3549
rect 15468 3519 15502 3553
rect 15638 3523 15672 3557
rect 15802 3519 15836 3553
rect 15972 3519 16006 3553
rect 16140 3515 16174 3549
rect 16308 3519 16342 3553
rect 16482 3515 16516 3549
rect 13572 3418 13606 3452
rect 13672 3418 13706 3452
rect 13772 3418 13806 3452
rect 13872 3418 13906 3452
rect 13972 3418 14006 3452
rect 14072 3418 14106 3452
rect 14172 3418 14206 3452
rect 14272 3418 14306 3452
rect 15232 3418 15266 3452
rect 15332 3418 15366 3452
rect 15432 3418 15466 3452
rect 15532 3418 15566 3452
rect 15632 3418 15666 3452
rect 15732 3418 15766 3452
rect 15832 3418 15866 3452
rect 15932 3418 15966 3452
<< metal1 >>
rect 14423 4747 14678 5103
rect 14423 4695 14443 4747
rect 14495 4695 14521 4747
rect 14573 4695 14614 4747
rect 14666 4695 14678 4747
rect 14423 4665 14678 4695
rect 44563 4747 44790 5115
rect 44563 4695 44594 4747
rect 44646 4695 44677 4747
rect 44729 4695 44790 4747
rect 44563 4661 44790 4695
rect 7079 4528 7615 4612
rect 22113 4537 22721 4595
rect 37217 4545 37841 4603
rect 52223 4551 52956 4609
rect 44732 3923 45399 3932
rect 44742 3874 45399 3923
rect 14642 3718 15291 3768
rect 14590 3710 15291 3718
rect 37381 3717 52816 3733
rect 37381 3715 44018 3717
rect 37381 3714 43682 3715
rect 37381 3713 37563 3714
rect 37381 3661 37460 3713
rect 37512 3662 37563 3713
rect 37615 3708 43682 3714
rect 37615 3674 43514 3708
rect 43548 3681 43682 3708
rect 43716 3705 44018 3715
rect 43716 3681 43850 3705
rect 43548 3674 43850 3681
rect 37615 3671 43850 3674
rect 43884 3683 44018 3705
rect 44052 3715 44350 3717
rect 44052 3683 44184 3715
rect 43884 3681 44184 3683
rect 44218 3683 44350 3715
rect 44384 3683 44518 3717
rect 44552 3715 45780 3717
rect 44552 3683 44692 3715
rect 44218 3681 44692 3683
rect 44726 3713 45780 3715
rect 44726 3709 45610 3713
rect 44726 3681 45448 3709
rect 43884 3675 45448 3681
rect 45482 3679 45610 3709
rect 45644 3683 45780 3713
rect 45814 3714 52816 3717
rect 45814 3713 52664 3714
rect 45814 3683 45944 3713
rect 45644 3679 45944 3683
rect 45978 3679 46114 3713
rect 46148 3709 46450 3713
rect 46148 3679 46282 3709
rect 45482 3675 46282 3679
rect 46316 3679 46450 3709
rect 46484 3709 52664 3713
rect 46484 3679 46624 3709
rect 46316 3675 46624 3679
rect 46658 3675 52573 3709
rect 43884 3671 52573 3675
rect 37615 3662 52573 3671
rect 37512 3661 52573 3662
rect 37381 3657 52573 3661
rect 52625 3662 52664 3709
rect 52716 3662 52816 3714
rect 52625 3657 52816 3662
rect 37381 3652 52816 3657
rect 43682 3612 46285 3618
rect 43682 3578 43714 3612
rect 43748 3578 43814 3612
rect 43848 3578 43914 3612
rect 43948 3578 44014 3612
rect 44048 3578 44114 3612
rect 44148 3578 44214 3612
rect 44248 3578 44314 3612
rect 44348 3578 44414 3612
rect 44448 3578 45374 3612
rect 45408 3578 45474 3612
rect 45508 3578 45574 3612
rect 45608 3578 45674 3612
rect 45708 3578 45774 3612
rect 45808 3578 45874 3612
rect 45908 3578 45974 3612
rect 46008 3578 46074 3612
rect 46108 3578 46285 3612
rect 43682 3573 46285 3578
rect 7224 3558 22590 3573
rect 43682 3570 45128 3573
rect 7224 3506 7265 3558
rect 7317 3506 7361 3558
rect 7413 3557 22590 3558
rect 7413 3555 13876 3557
rect 7413 3548 13540 3555
rect 7413 3514 13372 3548
rect 13406 3521 13540 3548
rect 13574 3545 13876 3555
rect 13574 3521 13708 3545
rect 13406 3514 13708 3521
rect 7413 3511 13708 3514
rect 13742 3523 13876 3545
rect 13910 3555 14208 3557
rect 13910 3523 14042 3555
rect 13742 3521 14042 3523
rect 14076 3523 14208 3555
rect 14242 3523 14376 3557
rect 14410 3555 15638 3557
rect 14410 3523 14550 3555
rect 14076 3521 14550 3523
rect 14584 3553 15638 3555
rect 14584 3549 15468 3553
rect 14584 3521 15306 3549
rect 13742 3515 15306 3521
rect 15340 3519 15468 3549
rect 15502 3523 15638 3553
rect 15672 3556 22590 3557
rect 15672 3553 22475 3556
rect 15672 3523 15802 3553
rect 15502 3519 15802 3523
rect 15836 3519 15972 3553
rect 16006 3549 16308 3553
rect 16006 3519 16140 3549
rect 15340 3515 16140 3519
rect 16174 3519 16308 3549
rect 16342 3549 22475 3553
rect 16342 3519 16482 3549
rect 16174 3515 16482 3519
rect 16516 3515 22376 3549
rect 13742 3511 22376 3515
rect 7413 3506 22376 3511
rect 7224 3497 22376 3506
rect 22428 3504 22475 3549
rect 22527 3504 22590 3556
rect 22428 3497 22590 3504
rect 7224 3492 22590 3497
rect 44978 3569 45128 3570
rect 44978 3517 45023 3569
rect 45075 3521 45128 3569
rect 45180 3570 46285 3573
rect 45180 3521 45206 3570
rect 45075 3517 45206 3521
rect 44978 3478 45206 3517
rect 13540 3452 16143 3458
rect 13540 3418 13572 3452
rect 13606 3418 13672 3452
rect 13706 3418 13772 3452
rect 13806 3418 13872 3452
rect 13906 3418 13972 3452
rect 14006 3418 14072 3452
rect 14106 3418 14172 3452
rect 14206 3418 14272 3452
rect 14306 3418 15232 3452
rect 15266 3418 15332 3452
rect 15366 3418 15432 3452
rect 15466 3418 15532 3452
rect 15566 3418 15632 3452
rect 15666 3418 15732 3452
rect 15766 3418 15832 3452
rect 15866 3418 15932 3452
rect 15966 3418 16143 3452
rect 13540 3413 16143 3418
rect 13540 3410 14986 3413
rect 14836 3409 14986 3410
rect 14836 3357 14881 3409
rect 14933 3361 14986 3409
rect 15038 3410 16143 3413
rect 15038 3361 15064 3410
rect 14933 3357 15064 3361
rect 14836 3318 15064 3357
rect 44732 3326 45484 3384
rect 13202 3148 13253 3244
rect 14590 3172 15271 3230
rect 19721 3175 45232 3219
rect 19721 3172 45120 3175
rect 13202 3147 13252 3148
rect 19721 3120 45031 3172
rect 45083 3123 45120 3172
rect 45172 3123 45232 3175
rect 45083 3120 45232 3123
rect 19721 3096 45232 3120
rect 19721 3044 45031 3096
rect 45083 3044 45124 3096
rect 45176 3044 45232 3096
rect 19721 3037 45232 3044
rect 14848 3013 45232 3037
rect 14848 2992 19927 3013
rect 14848 2940 14885 2992
rect 14937 2987 19927 2992
rect 14937 2940 14979 2987
rect 14848 2935 14979 2940
rect 15031 2935 19927 2987
rect 14848 2914 19927 2935
rect 14848 2912 14979 2914
rect 7015 2840 7678 2898
rect 14848 2860 14885 2912
rect 14937 2862 14979 2912
rect 15031 2862 19927 2914
rect 14937 2860 19927 2862
rect 14848 2831 19927 2860
rect 22113 2852 22741 2910
rect 37125 2852 37888 2910
rect 52315 2843 52966 2901
rect 60382 780 60604 858
<< via1 >>
rect 7264 4761 7316 4813
rect 7345 4760 7397 4812
rect 22380 4758 22432 4810
rect 22475 4758 22527 4810
rect 37457 4760 37509 4812
rect 37559 4760 37611 4812
rect 14443 4695 14495 4747
rect 14521 4695 14573 4747
rect 14614 4695 14666 4747
rect 44594 4695 44646 4747
rect 44677 4695 44729 4747
rect 52575 4733 52627 4785
rect 52670 4733 52722 4785
rect 6272 4537 6324 4589
rect 6379 4539 6431 4591
rect 6481 4539 6533 4591
rect 6581 4540 6633 4592
rect 21302 4543 21354 4595
rect 21405 4543 21457 4595
rect 21488 4543 21540 4595
rect 21589 4543 21641 4595
rect 21676 4543 21728 4595
rect 36434 4539 36486 4591
rect 36522 4539 36574 4591
rect 36607 4544 36659 4596
rect 53350 4536 53402 4588
rect 53444 4536 53496 4588
rect 53521 4536 53573 4588
rect 53601 4535 53653 4587
rect 53675 4536 53727 4588
rect 44600 3870 44652 3922
rect 44690 3871 44742 3923
rect 14467 3718 14519 3770
rect 14590 3718 14642 3770
rect 37460 3661 37512 3713
rect 37563 3662 37615 3714
rect 52573 3657 52625 3709
rect 52664 3662 52716 3714
rect 7265 3506 7317 3558
rect 7361 3506 7413 3558
rect 22376 3497 22428 3549
rect 22475 3504 22527 3556
rect 45023 3517 45075 3569
rect 45128 3521 45180 3573
rect 14881 3357 14933 3409
rect 14986 3361 15038 3413
rect 46035 3330 46087 3382
rect 46127 3331 46179 3383
rect 46217 3330 46269 3382
rect 46305 3329 46357 3381
rect 13680 3169 13732 3221
rect 13764 3169 13816 3221
rect 13857 3170 13909 3222
rect 45031 3120 45083 3172
rect 45120 3123 45172 3175
rect 45031 3044 45083 3096
rect 45124 3044 45176 3096
rect 14885 2940 14937 2992
rect 14979 2935 15031 2987
rect 6266 2843 6318 2895
rect 6364 2843 6416 2895
rect 6459 2843 6511 2895
rect 6564 2843 6616 2895
rect 14885 2860 14937 2912
rect 14979 2862 15031 2914
rect 21316 2848 21368 2900
rect 21416 2848 21468 2900
rect 21515 2848 21567 2900
rect 21618 2848 21670 2900
rect 36424 2842 36476 2894
rect 36512 2842 36564 2894
rect 36610 2838 36662 2890
rect 53346 2839 53398 2891
rect 53434 2839 53486 2891
rect 53517 2839 53569 2891
rect 53604 2839 53656 2891
rect 7265 2623 7317 2675
rect 7345 2621 7397 2673
rect 22381 2638 22433 2690
rect 22464 2638 22516 2690
rect 37459 2628 37511 2680
rect 37550 2628 37602 2680
rect 52576 2613 52628 2665
rect 52659 2613 52711 2665
<< metal2 >>
rect 7240 4813 7429 4843
rect 7240 4761 7264 4813
rect 7316 4812 7429 4813
rect 7316 4761 7345 4812
rect 7240 4760 7345 4761
rect 7397 4760 7429 4812
rect 6208 4592 6692 4719
rect 6208 4591 6581 4592
rect 6208 4589 6379 4591
rect 6208 4537 6272 4589
rect 6324 4539 6379 4589
rect 6431 4539 6481 4591
rect 6533 4540 6581 4591
rect 6633 4540 6692 4592
rect 6533 4539 6692 4540
rect 6324 4537 6692 4539
rect 6208 3372 6692 4537
rect 6208 3316 6275 3372
rect 6331 3316 6389 3372
rect 6445 3316 6503 3372
rect 6559 3316 6692 3372
rect 6208 3257 6692 3316
rect 6208 3201 6275 3257
rect 6331 3201 6389 3257
rect 6445 3201 6503 3257
rect 6559 3201 6692 3257
rect 6208 3142 6692 3201
rect 6208 3086 6275 3142
rect 6331 3086 6389 3142
rect 6445 3086 6503 3142
rect 6559 3086 6692 3142
rect 6208 2895 6692 3086
rect 6208 2843 6266 2895
rect 6318 2843 6364 2895
rect 6416 2843 6459 2895
rect 6511 2843 6564 2895
rect 6616 2843 6692 2895
rect 6208 2729 6692 2843
rect 7240 3558 7429 4760
rect 14423 4747 14683 4818
rect 14423 4695 14443 4747
rect 14495 4695 14521 4747
rect 14573 4695 14614 4747
rect 14666 4695 14683 4747
rect 22351 4810 22540 4833
rect 22351 4758 22380 4810
rect 22432 4758 22475 4810
rect 22527 4758 22540 4810
rect 14423 3770 14683 4695
rect 14423 3718 14467 3770
rect 14519 3718 14590 3770
rect 14642 3718 14683 3770
rect 14423 3674 14683 3718
rect 21264 4595 21731 4697
rect 21264 4543 21302 4595
rect 21354 4543 21405 4595
rect 21457 4543 21488 4595
rect 21540 4543 21589 4595
rect 21641 4543 21676 4595
rect 21728 4543 21731 4595
rect 7240 3506 7265 3558
rect 7317 3506 7361 3558
rect 7413 3506 7429 3558
rect 7240 2675 7429 3506
rect 14848 3413 15054 3458
rect 14848 3409 14986 3413
rect 14848 3357 14881 3409
rect 14933 3361 14986 3409
rect 15038 3361 15054 3413
rect 14933 3357 15054 3361
rect 7240 2623 7265 2675
rect 7317 2673 7429 2675
rect 7317 2623 7345 2673
rect 7240 2621 7345 2623
rect 7397 2621 7429 2673
rect 13629 3222 13982 3268
rect 13629 3221 13857 3222
rect 13629 3169 13680 3221
rect 13732 3169 13764 3221
rect 13816 3170 13857 3221
rect 13909 3170 13982 3222
rect 13816 3169 13982 3170
rect 13629 2811 13982 3169
rect 14848 2992 15054 3357
rect 14848 2940 14885 2992
rect 14937 2987 15054 2992
rect 14937 2940 14979 2987
rect 14848 2935 14979 2940
rect 15031 2935 15054 2987
rect 14848 2914 15054 2935
rect 14848 2912 14979 2914
rect 14848 2860 14885 2912
rect 14937 2862 14979 2912
rect 15031 2862 15054 2914
rect 14937 2860 15054 2862
rect 14848 2831 15054 2860
rect 21264 3282 21731 4543
rect 21264 3226 21314 3282
rect 21370 3226 21418 3282
rect 21474 3226 21522 3282
rect 21578 3226 21626 3282
rect 21682 3226 21731 3282
rect 21264 3166 21731 3226
rect 21264 3110 21314 3166
rect 21370 3110 21418 3166
rect 21474 3110 21522 3166
rect 21578 3110 21626 3166
rect 21682 3110 21731 3166
rect 21264 3050 21731 3110
rect 21264 2994 21314 3050
rect 21370 2994 21418 3050
rect 21474 2994 21522 3050
rect 21578 2994 21626 3050
rect 21682 2994 21731 3050
rect 21264 2900 21731 2994
rect 21264 2848 21316 2900
rect 21368 2848 21416 2900
rect 21468 2848 21515 2900
rect 21567 2848 21618 2900
rect 21670 2848 21731 2900
rect 13629 2755 13669 2811
rect 13725 2755 13777 2811
rect 13833 2755 13885 2811
rect 13941 2755 13982 2811
rect 13629 2717 13982 2755
rect 21264 2746 21731 2848
rect 22351 3556 22540 4758
rect 37442 4812 37629 4831
rect 37442 4760 37457 4812
rect 37509 4760 37559 4812
rect 37611 4760 37629 4812
rect 22351 3549 22475 3556
rect 22351 3497 22376 3549
rect 22428 3504 22475 3549
rect 22527 3504 22540 3556
rect 22428 3497 22540 3504
rect 13629 2661 13669 2717
rect 13725 2661 13777 2717
rect 13833 2661 13885 2717
rect 13941 2661 13982 2717
rect 13629 2635 13982 2661
rect 22351 2690 22540 3497
rect 36380 4596 36680 4695
rect 36380 4591 36607 4596
rect 36380 4539 36434 4591
rect 36486 4539 36522 4591
rect 36574 4544 36607 4591
rect 36659 4544 36680 4596
rect 36574 4539 36680 4544
rect 36380 3631 36680 4539
rect 36380 3575 36401 3631
rect 36457 3575 36495 3631
rect 36551 3575 36589 3631
rect 36645 3575 36680 3631
rect 36380 3543 36680 3575
rect 36380 3487 36401 3543
rect 36457 3487 36495 3543
rect 36551 3487 36589 3543
rect 36645 3487 36680 3543
rect 36380 3455 36680 3487
rect 36380 3399 36401 3455
rect 36457 3399 36495 3455
rect 36551 3399 36589 3455
rect 36645 3399 36680 3455
rect 36380 2894 36680 3399
rect 36380 2842 36424 2894
rect 36476 2842 36512 2894
rect 36564 2890 36680 2894
rect 36564 2842 36610 2890
rect 36380 2838 36610 2842
rect 36662 2838 36680 2890
rect 36380 2743 36680 2838
rect 37442 3714 37629 4760
rect 44571 4747 44790 4800
rect 44571 4695 44594 4747
rect 44646 4695 44677 4747
rect 44729 4695 44790 4747
rect 44571 3923 44790 4695
rect 44571 3922 44690 3923
rect 44571 3870 44600 3922
rect 44652 3871 44690 3922
rect 44742 3871 44790 3923
rect 44652 3870 44790 3871
rect 44571 3835 44790 3870
rect 52546 4785 52735 4808
rect 52546 4733 52575 4785
rect 52627 4733 52670 4785
rect 52722 4733 52735 4785
rect 37442 3713 37563 3714
rect 37442 3661 37460 3713
rect 37512 3662 37563 3713
rect 37615 3662 37629 3714
rect 37512 3661 37629 3662
rect 22351 2638 22381 2690
rect 22433 2638 22464 2690
rect 22516 2638 22540 2690
rect 22351 2625 22540 2638
rect 37442 2680 37629 3661
rect 52546 3714 52735 4733
rect 52546 3709 52664 3714
rect 52546 3657 52573 3709
rect 52625 3662 52664 3709
rect 52716 3662 52735 3714
rect 52625 3657 52735 3662
rect 44990 3573 45196 3618
rect 44990 3569 45128 3573
rect 44990 3517 45023 3569
rect 45075 3521 45128 3569
rect 45180 3521 45196 3573
rect 45075 3517 45196 3521
rect 44990 3175 45196 3517
rect 44990 3172 45120 3175
rect 44990 3120 45031 3172
rect 45083 3123 45120 3172
rect 45172 3123 45196 3175
rect 45083 3120 45196 3123
rect 44990 3096 45196 3120
rect 44990 3044 45031 3096
rect 45083 3044 45124 3096
rect 45176 3044 45196 3096
rect 44990 3001 45196 3044
rect 45998 3383 46412 3405
rect 45998 3382 46127 3383
rect 45998 3330 46035 3382
rect 46087 3331 46127 3382
rect 46179 3382 46412 3383
rect 46179 3331 46217 3382
rect 46087 3330 46217 3331
rect 46269 3381 46412 3382
rect 46269 3330 46305 3381
rect 45998 3329 46305 3330
rect 46357 3329 46412 3381
rect 37442 2628 37459 2680
rect 37511 2628 37550 2680
rect 37602 2628 37629 2680
rect 7240 2603 7429 2621
rect 37442 2620 37629 2628
rect 45998 2784 46412 3329
rect 45998 2728 46035 2784
rect 46091 2728 46128 2784
rect 46184 2728 46221 2784
rect 46277 2728 46314 2784
rect 46370 2728 46412 2784
rect 45998 2702 46412 2728
rect 45998 2646 46035 2702
rect 46091 2646 46128 2702
rect 46184 2646 46221 2702
rect 46277 2646 46314 2702
rect 46370 2646 46412 2702
rect 45998 2609 46412 2646
rect 52546 2665 52735 3657
rect 53311 4588 53732 4695
rect 53311 4536 53350 4588
rect 53402 4536 53444 4588
rect 53496 4536 53521 4588
rect 53573 4587 53675 4588
rect 53573 4536 53601 4587
rect 53311 4535 53601 4536
rect 53653 4536 53675 4587
rect 53727 4536 53732 4588
rect 53653 4535 53732 4536
rect 53311 3176 53732 4535
rect 53311 3120 53348 3176
rect 53404 3120 53452 3176
rect 53508 3120 53556 3176
rect 53612 3120 53660 3176
rect 53716 3120 53732 3176
rect 53311 3086 53732 3120
rect 53311 3030 53348 3086
rect 53404 3030 53452 3086
rect 53508 3030 53556 3086
rect 53612 3030 53660 3086
rect 53716 3030 53732 3086
rect 53311 2891 53732 3030
rect 53311 2839 53346 2891
rect 53398 2839 53434 2891
rect 53486 2839 53517 2891
rect 53569 2839 53604 2891
rect 53656 2839 53732 2891
rect 53311 2745 53732 2839
rect 52546 2613 52576 2665
rect 52628 2613 52659 2665
rect 52711 2613 52735 2665
rect 52546 2600 52735 2613
<< via2 >>
rect 6275 3316 6331 3372
rect 6389 3316 6445 3372
rect 6503 3316 6559 3372
rect 6275 3201 6331 3257
rect 6389 3201 6445 3257
rect 6503 3201 6559 3257
rect 6275 3086 6331 3142
rect 6389 3086 6445 3142
rect 6503 3086 6559 3142
rect 21314 3226 21370 3282
rect 21418 3226 21474 3282
rect 21522 3226 21578 3282
rect 21626 3226 21682 3282
rect 21314 3110 21370 3166
rect 21418 3110 21474 3166
rect 21522 3110 21578 3166
rect 21626 3110 21682 3166
rect 21314 2994 21370 3050
rect 21418 2994 21474 3050
rect 21522 2994 21578 3050
rect 21626 2994 21682 3050
rect 13669 2755 13725 2811
rect 13777 2755 13833 2811
rect 13885 2755 13941 2811
rect 13669 2661 13725 2717
rect 13777 2661 13833 2717
rect 13885 2661 13941 2717
rect 36401 3575 36457 3631
rect 36495 3575 36551 3631
rect 36589 3575 36645 3631
rect 36401 3487 36457 3543
rect 36495 3487 36551 3543
rect 36589 3487 36645 3543
rect 36401 3399 36457 3455
rect 36495 3399 36551 3455
rect 36589 3399 36645 3455
rect 46035 2728 46091 2784
rect 46128 2728 46184 2784
rect 46221 2728 46277 2784
rect 46314 2728 46370 2784
rect 46035 2646 46091 2702
rect 46128 2646 46184 2702
rect 46221 2646 46277 2702
rect 46314 2646 46370 2702
rect 53348 3120 53404 3176
rect 53452 3120 53508 3176
rect 53556 3120 53612 3176
rect 53660 3120 53716 3176
rect 53348 3030 53404 3086
rect 53452 3030 53508 3086
rect 53556 3030 53612 3086
rect 53660 3030 53716 3086
<< metal3 >>
rect 2518 7372 2624 7389
rect 2518 7308 2539 7372
rect 2603 7308 2624 7372
rect 2518 7292 2624 7308
rect 2518 7228 2539 7292
rect 2603 7228 2624 7292
rect 2518 7211 2624 7228
rect 2727 7371 2833 7388
rect 2727 7307 2748 7371
rect 2812 7307 2833 7371
rect 2727 7291 2833 7307
rect 2727 7227 2748 7291
rect 2812 7227 2833 7291
rect 2727 7210 2833 7227
rect 2893 7371 2999 7388
rect 2893 7307 2914 7371
rect 2978 7307 2999 7371
rect 2893 7291 2999 7307
rect 2893 7227 2914 7291
rect 2978 7227 2999 7291
rect 2893 7210 2999 7227
rect 3073 7373 3179 7390
rect 3073 7309 3094 7373
rect 3158 7309 3179 7373
rect 3073 7293 3179 7309
rect 3073 7229 3094 7293
rect 3158 7229 3179 7293
rect 3073 7212 3179 7229
rect 1284 5254 1390 5271
rect 1284 5190 1305 5254
rect 1369 5190 1390 5254
rect 1284 5174 1390 5190
rect 1284 5110 1305 5174
rect 1369 5110 1390 5174
rect 1284 5093 1390 5110
rect 1456 5255 1562 5272
rect 1456 5191 1477 5255
rect 1541 5191 1562 5255
rect 1456 5175 1562 5191
rect 1456 5111 1477 5175
rect 1541 5111 1562 5175
rect 1456 5094 1562 5111
rect 1630 5254 1736 5271
rect 1630 5190 1651 5254
rect 1715 5190 1736 5254
rect 1630 5174 1736 5190
rect 1630 5110 1651 5174
rect 1715 5110 1736 5174
rect 1630 5093 1736 5110
rect 36378 3631 36682 3645
rect 36378 3575 36401 3631
rect 36457 3575 36495 3631
rect 36551 3575 36589 3631
rect 36645 3575 36682 3631
rect 36378 3543 36682 3575
rect 36378 3487 36401 3543
rect 36457 3508 36495 3543
rect 36489 3487 36495 3508
rect 36551 3509 36589 3543
rect 36551 3487 36579 3509
rect 36645 3487 36682 3543
rect 36378 3455 36425 3487
rect 36489 3455 36579 3487
rect 36643 3455 36682 3487
rect 6274 3398 6616 3431
rect 36378 3399 36401 3455
rect 36489 3444 36495 3455
rect 36457 3399 36495 3444
rect 36551 3445 36579 3455
rect 36551 3399 36589 3445
rect 36645 3399 36682 3455
rect 6206 3372 6695 3398
rect 36378 3379 36682 3399
rect 6206 3316 6275 3372
rect 6331 3316 6389 3372
rect 6445 3316 6503 3372
rect 6559 3316 6695 3372
rect 6206 3257 6695 3316
rect 6206 3201 6275 3257
rect 6331 3215 6389 3257
rect 6445 3221 6503 3257
rect 6347 3201 6389 3215
rect 6498 3201 6503 3221
rect 6559 3221 6695 3257
rect 6559 3201 6579 3221
rect 6206 3151 6283 3201
rect 6347 3157 6434 3201
rect 6498 3157 6579 3201
rect 6643 3157 6695 3221
rect 6347 3151 6695 3157
rect 6206 3142 6695 3151
rect 6206 3086 6275 3142
rect 6331 3086 6389 3142
rect 6445 3086 6503 3142
rect 6559 3086 6695 3142
rect 6206 3031 6695 3086
rect 21264 3282 21731 3336
rect 21264 3226 21314 3282
rect 21370 3229 21418 3282
rect 21390 3226 21418 3229
rect 21474 3229 21522 3282
rect 21474 3226 21493 3229
rect 21578 3226 21626 3282
rect 21682 3226 21731 3282
rect 21264 3166 21326 3226
rect 21390 3166 21493 3226
rect 21557 3166 21731 3226
rect 21264 3110 21314 3166
rect 21390 3165 21418 3166
rect 21370 3110 21418 3165
rect 21474 3165 21493 3166
rect 21474 3110 21522 3165
rect 21578 3110 21626 3166
rect 21682 3110 21731 3166
rect 21264 3068 21731 3110
rect 21264 3050 21326 3068
rect 21390 3050 21493 3068
rect 21557 3050 21731 3068
rect 21264 2994 21314 3050
rect 21390 3004 21418 3050
rect 21370 2994 21418 3004
rect 21474 3004 21493 3050
rect 21474 2994 21522 3004
rect 21578 2994 21626 3050
rect 21682 2994 21731 3050
rect 53311 3176 53733 3204
rect 53311 3120 53348 3176
rect 53429 3120 53452 3176
rect 53550 3120 53556 3176
rect 53612 3120 53624 3176
rect 53716 3120 53733 3176
rect 53311 3112 53365 3120
rect 53429 3112 53486 3120
rect 53550 3112 53624 3120
rect 53688 3112 53733 3120
rect 53311 3096 53733 3112
rect 53311 3086 53365 3096
rect 53429 3086 53486 3096
rect 53550 3086 53624 3096
rect 53688 3086 53733 3096
rect 53311 3030 53348 3086
rect 53429 3032 53452 3086
rect 53550 3032 53556 3086
rect 53404 3030 53452 3032
rect 53508 3030 53556 3032
rect 53612 3032 53624 3086
rect 53612 3030 53660 3032
rect 53716 3030 53733 3086
rect 53311 2996 53733 3030
rect 21264 2950 21731 2994
rect 13629 2811 13982 2834
rect 13629 2760 13669 2811
rect 13725 2760 13777 2811
rect 13833 2760 13885 2811
rect 13629 2696 13659 2760
rect 13725 2755 13762 2760
rect 13833 2755 13865 2760
rect 13941 2755 13982 2811
rect 13723 2717 13762 2755
rect 13826 2717 13865 2755
rect 13929 2717 13982 2755
rect 13725 2696 13762 2717
rect 13833 2696 13865 2717
rect 13629 2661 13669 2696
rect 13725 2661 13777 2696
rect 13833 2661 13885 2696
rect 13941 2661 13982 2717
rect 13629 2635 13982 2661
rect 45998 2801 46413 2851
rect 45998 2800 46186 2801
rect 45998 2784 46046 2800
rect 46110 2784 46186 2800
rect 46250 2784 46314 2801
rect 45998 2728 46035 2784
rect 46110 2736 46128 2784
rect 46091 2728 46128 2736
rect 46184 2737 46186 2784
rect 46184 2728 46221 2737
rect 46277 2728 46314 2784
rect 46378 2737 46413 2801
rect 46370 2728 46413 2737
rect 45998 2721 46413 2728
rect 45998 2720 46186 2721
rect 45998 2702 46046 2720
rect 46110 2702 46186 2720
rect 46250 2702 46314 2721
rect 45998 2646 46035 2702
rect 46110 2656 46128 2702
rect 46091 2646 46128 2656
rect 46184 2657 46186 2702
rect 46184 2646 46221 2657
rect 46277 2646 46314 2702
rect 46378 2657 46413 2721
rect 46370 2646 46413 2657
rect 45998 2610 46413 2646
rect 1286 2306 1392 2323
rect 1286 2242 1307 2306
rect 1371 2242 1392 2306
rect 1286 2226 1392 2242
rect 1286 2162 1307 2226
rect 1371 2162 1392 2226
rect 1286 2145 1392 2162
rect 1491 2308 1597 2325
rect 1491 2244 1512 2308
rect 1576 2244 1597 2308
rect 1491 2228 1597 2244
rect 1491 2164 1512 2228
rect 1576 2164 1597 2228
rect 1491 2147 1597 2164
rect 1690 2308 1796 2325
rect 1690 2244 1711 2308
rect 1775 2244 1796 2308
rect 1690 2228 1796 2244
rect 1690 2164 1711 2228
rect 1775 2164 1796 2228
rect 1690 2147 1796 2164
rect 2532 195 2638 212
rect 2532 131 2553 195
rect 2617 131 2638 195
rect 2532 115 2638 131
rect 2532 51 2553 115
rect 2617 51 2638 115
rect 2532 34 2638 51
rect 2753 195 2859 212
rect 2753 131 2774 195
rect 2838 131 2859 195
rect 2753 115 2859 131
rect 2753 51 2774 115
rect 2838 51 2859 115
rect 2753 34 2859 51
rect 2962 195 3068 212
rect 2962 131 2983 195
rect 3047 131 3068 195
rect 2962 115 3068 131
rect 2962 51 2983 115
rect 3047 51 3068 115
rect 2962 34 3068 51
rect 3136 195 3242 212
rect 3136 131 3157 195
rect 3221 131 3242 195
rect 13779 206 13856 209
rect 3136 115 3242 131
rect 3136 51 3157 115
rect 3221 51 3242 115
rect 6260 143 6346 157
rect 6260 79 6271 143
rect 6335 79 6346 143
rect 6260 66 6346 79
rect 6408 143 6494 157
rect 6408 79 6419 143
rect 6483 79 6494 143
rect 6408 66 6494 79
rect 6556 143 6642 157
rect 6556 79 6567 143
rect 6631 79 6642 143
rect 13779 142 13785 206
rect 13849 142 13856 206
rect 53361 193 53445 200
rect 46038 183 46122 190
rect 13779 140 13856 142
rect 21317 147 21413 169
rect 6556 66 6642 79
rect 13802 87 13879 90
rect 3136 34 3242 51
rect 13802 23 13808 87
rect 13872 23 13879 87
rect 21317 83 21333 147
rect 21397 83 21413 147
rect 21317 61 21413 83
rect 21450 147 21546 169
rect 21450 83 21466 147
rect 21530 83 21546 147
rect 21450 61 21546 83
rect 21583 147 21679 169
rect 21583 83 21599 147
rect 21663 83 21679 147
rect 21583 61 21679 83
rect 36412 133 36499 157
rect 36412 69 36423 133
rect 36487 69 36499 133
rect 36412 45 36499 69
rect 36581 133 36668 157
rect 36581 69 36592 133
rect 36656 69 36668 133
rect 36581 45 36668 69
rect 46038 119 46048 183
rect 46112 119 46122 183
rect 46038 103 46122 119
rect 46038 39 46048 103
rect 46112 39 46122 103
rect 46038 32 46122 39
rect 46151 183 46235 190
rect 46151 119 46161 183
rect 46225 119 46235 183
rect 46151 103 46235 119
rect 46151 39 46161 103
rect 46225 39 46235 103
rect 46151 32 46235 39
rect 46266 183 46350 190
rect 46266 119 46276 183
rect 46340 119 46350 183
rect 46266 103 46350 119
rect 46266 39 46276 103
rect 46340 39 46350 103
rect 53361 129 53371 193
rect 53435 129 53445 193
rect 53361 113 53445 129
rect 53361 49 53371 113
rect 53435 49 53445 113
rect 53361 42 53445 49
rect 53480 193 53564 200
rect 53480 129 53490 193
rect 53554 129 53564 193
rect 53480 113 53564 129
rect 53480 49 53490 113
rect 53554 49 53564 113
rect 53480 42 53564 49
rect 53609 193 53693 200
rect 53609 129 53619 193
rect 53683 129 53693 193
rect 53609 113 53693 129
rect 53609 49 53619 113
rect 53683 49 53693 113
rect 53609 42 53693 49
rect 46266 32 46350 39
rect 13802 21 13879 23
<< via3 >>
rect 2539 7308 2603 7372
rect 2539 7228 2603 7292
rect 2748 7307 2812 7371
rect 2748 7227 2812 7291
rect 2914 7307 2978 7371
rect 2914 7227 2978 7291
rect 3094 7309 3158 7373
rect 3094 7229 3158 7293
rect 1305 5190 1369 5254
rect 1305 5110 1369 5174
rect 1477 5191 1541 5255
rect 1477 5111 1541 5175
rect 1651 5190 1715 5254
rect 1651 5110 1715 5174
rect 36425 3487 36457 3508
rect 36457 3487 36489 3508
rect 36579 3487 36589 3509
rect 36589 3487 36643 3509
rect 36425 3455 36489 3487
rect 36579 3455 36643 3487
rect 36425 3444 36457 3455
rect 36457 3444 36489 3455
rect 36579 3445 36589 3455
rect 36589 3445 36643 3455
rect 6283 3201 6331 3215
rect 6331 3201 6347 3215
rect 6434 3201 6445 3221
rect 6445 3201 6498 3221
rect 6283 3151 6347 3201
rect 6434 3157 6498 3201
rect 6579 3157 6643 3221
rect 21326 3226 21370 3229
rect 21370 3226 21390 3229
rect 21493 3226 21522 3229
rect 21522 3226 21557 3229
rect 21326 3166 21390 3226
rect 21493 3166 21557 3226
rect 21326 3165 21370 3166
rect 21370 3165 21390 3166
rect 21493 3165 21522 3166
rect 21522 3165 21557 3166
rect 21326 3050 21390 3068
rect 21493 3050 21557 3068
rect 21326 3004 21370 3050
rect 21370 3004 21390 3050
rect 21493 3004 21522 3050
rect 21522 3004 21557 3050
rect 53365 3120 53404 3176
rect 53404 3120 53429 3176
rect 53486 3120 53508 3176
rect 53508 3120 53550 3176
rect 53624 3120 53660 3176
rect 53660 3120 53688 3176
rect 53365 3112 53429 3120
rect 53486 3112 53550 3120
rect 53624 3112 53688 3120
rect 53365 3086 53429 3096
rect 53486 3086 53550 3096
rect 53624 3086 53688 3096
rect 53365 3032 53404 3086
rect 53404 3032 53429 3086
rect 53486 3032 53508 3086
rect 53508 3032 53550 3086
rect 53624 3032 53660 3086
rect 53660 3032 53688 3086
rect 13659 2755 13669 2760
rect 13669 2755 13723 2760
rect 13762 2755 13777 2760
rect 13777 2755 13826 2760
rect 13865 2755 13885 2760
rect 13885 2755 13929 2760
rect 13659 2717 13723 2755
rect 13762 2717 13826 2755
rect 13865 2717 13929 2755
rect 13659 2696 13669 2717
rect 13669 2696 13723 2717
rect 13762 2696 13777 2717
rect 13777 2696 13826 2717
rect 13865 2696 13885 2717
rect 13885 2696 13929 2717
rect 46046 2784 46110 2800
rect 46186 2784 46250 2801
rect 46314 2784 46378 2801
rect 46046 2736 46091 2784
rect 46091 2736 46110 2784
rect 46186 2737 46221 2784
rect 46221 2737 46250 2784
rect 46314 2737 46370 2784
rect 46370 2737 46378 2784
rect 46046 2702 46110 2720
rect 46186 2702 46250 2721
rect 46314 2702 46378 2721
rect 46046 2656 46091 2702
rect 46091 2656 46110 2702
rect 46186 2657 46221 2702
rect 46221 2657 46250 2702
rect 46314 2657 46370 2702
rect 46370 2657 46378 2702
rect 1307 2242 1371 2306
rect 1307 2162 1371 2226
rect 1512 2244 1576 2308
rect 1512 2164 1576 2228
rect 1711 2244 1775 2308
rect 1711 2164 1775 2228
rect 2553 131 2617 195
rect 2553 51 2617 115
rect 2774 131 2838 195
rect 2774 51 2838 115
rect 2983 131 3047 195
rect 2983 51 3047 115
rect 3157 131 3221 195
rect 3157 51 3221 115
rect 6271 79 6335 143
rect 6419 79 6483 143
rect 6567 79 6631 143
rect 13785 142 13849 206
rect 13808 23 13872 87
rect 21333 83 21397 147
rect 21466 83 21530 147
rect 21599 83 21663 147
rect 36423 69 36487 133
rect 36592 69 36656 133
rect 46048 119 46112 183
rect 46048 39 46112 103
rect 46161 119 46225 183
rect 46161 39 46225 103
rect 46276 119 46340 183
rect 46276 39 46340 103
rect 53371 129 53435 193
rect 53371 49 53435 113
rect 53490 129 53554 193
rect 53490 49 53554 113
rect 53619 129 53683 193
rect 53619 49 53683 113
<< metal4 >>
rect 2467 7373 3251 7443
rect 2467 7372 3094 7373
rect 2467 7308 2539 7372
rect 2603 7371 3094 7372
rect 2603 7308 2748 7371
rect 2467 7307 2748 7308
rect 2812 7307 2914 7371
rect 2978 7309 3094 7371
rect 3158 7309 3251 7373
rect 2978 7307 3251 7309
rect 2467 7293 3251 7307
rect 2467 7292 3094 7293
rect 2467 7228 2539 7292
rect 2603 7291 3094 7292
rect 2603 7228 2748 7291
rect 2467 7227 2748 7228
rect 2812 7227 2914 7291
rect 2978 7229 3094 7291
rect 3158 7229 3251 7293
rect 2978 7227 3251 7229
rect 1234 5255 1852 5401
rect 1234 5254 1477 5255
rect 1234 5190 1305 5254
rect 1369 5191 1477 5254
rect 1541 5254 1852 5255
rect 1541 5191 1651 5254
rect 1369 5190 1651 5191
rect 1715 5190 1852 5254
rect 1234 5175 1852 5190
rect 1234 5174 1477 5175
rect 1234 5110 1305 5174
rect 1369 5111 1477 5174
rect 1541 5174 1852 5175
rect 1541 5111 1651 5174
rect 1369 5110 1651 5111
rect 1715 5110 1852 5174
rect 1234 2308 1852 5110
rect 1234 2306 1512 2308
rect 1234 2242 1307 2306
rect 1371 2244 1512 2306
rect 1576 2244 1711 2308
rect 1775 2244 1852 2308
rect 1371 2242 1852 2244
rect 1234 2228 1852 2242
rect 1234 2226 1512 2228
rect 1234 2162 1307 2226
rect 1371 2164 1512 2226
rect 1576 2164 1711 2228
rect 1775 2164 1852 2228
rect 1371 2162 1852 2164
rect 1234 2095 1852 2162
rect 2467 195 3251 7227
rect 36378 3509 36683 3690
rect 36378 3508 36579 3509
rect 36378 3444 36425 3508
rect 36489 3445 36579 3508
rect 36643 3445 36683 3509
rect 36489 3444 36683 3445
rect 2467 131 2553 195
rect 2617 131 2774 195
rect 2838 131 2983 195
rect 3047 131 3157 195
rect 3221 131 3251 195
rect 2467 115 3251 131
rect 2467 51 2553 115
rect 2617 51 2774 115
rect 2838 51 2983 115
rect 3047 51 3157 115
rect 3221 51 3251 115
rect 2467 -55 3251 51
rect 6214 3221 6683 3350
rect 6214 3215 6434 3221
rect 6214 3151 6283 3215
rect 6347 3157 6434 3215
rect 6498 3157 6579 3221
rect 6643 3157 6683 3221
rect 6347 3151 6683 3157
rect 6214 143 6683 3151
rect 21264 3229 21731 3364
rect 21264 3165 21326 3229
rect 21390 3165 21493 3229
rect 21557 3165 21731 3229
rect 21264 3068 21731 3165
rect 21264 3004 21326 3068
rect 21390 3004 21493 3068
rect 21557 3004 21731 3068
rect 13629 2760 13983 2835
rect 13629 2696 13659 2760
rect 13723 2696 13762 2760
rect 13826 2696 13865 2760
rect 13929 2696 13983 2760
rect 13629 2634 13983 2696
rect 6214 79 6271 143
rect 6335 79 6419 143
rect 6483 79 6567 143
rect 6631 79 6683 143
rect 6214 -33 6683 79
rect 13705 206 13906 2634
rect 13705 142 13785 206
rect 13849 142 13906 206
rect 13705 87 13906 142
rect 13705 23 13808 87
rect 13872 23 13906 87
rect 13705 -58 13906 23
rect 21264 147 21731 3004
rect 21264 83 21333 147
rect 21397 83 21466 147
rect 21530 83 21599 147
rect 21663 83 21731 147
rect 21264 -8 21731 83
rect 36378 133 36683 3444
rect 53311 3176 53736 3206
rect 53311 3112 53365 3176
rect 53429 3112 53486 3176
rect 53550 3112 53624 3176
rect 53688 3112 53736 3176
rect 53311 3096 53736 3112
rect 53311 3032 53365 3096
rect 53429 3032 53486 3096
rect 53550 3032 53624 3096
rect 53688 3032 53736 3096
rect 36378 69 36423 133
rect 36487 69 36592 133
rect 36656 69 36683 133
rect 36378 -3 36683 69
rect 45998 2801 46412 2897
rect 45998 2800 46186 2801
rect 45998 2736 46046 2800
rect 46110 2737 46186 2800
rect 46250 2737 46314 2801
rect 46378 2737 46412 2801
rect 46110 2736 46412 2737
rect 45998 2721 46412 2736
rect 45998 2720 46186 2721
rect 45998 2656 46046 2720
rect 46110 2657 46186 2720
rect 46250 2657 46314 2721
rect 46378 2657 46412 2721
rect 46110 2656 46412 2657
rect 45998 183 46412 2656
rect 45998 119 46048 183
rect 46112 119 46161 183
rect 46225 119 46276 183
rect 46340 119 46412 183
rect 45998 103 46412 119
rect 45998 39 46048 103
rect 46112 39 46161 103
rect 46225 39 46276 103
rect 46340 39 46412 103
rect 45998 -56 46412 39
rect 53311 193 53736 3032
rect 53311 129 53371 193
rect 53435 129 53490 193
rect 53554 129 53619 193
rect 53683 129 53736 193
rect 53311 113 53736 129
rect 53311 49 53371 113
rect 53435 49 53490 113
rect 53554 49 53619 113
rect 53683 49 53736 113
rect 53311 -44 53736 49
use brbufhalf  brbufhalf_0
timestamp 1656715967
transform -1 0 26228 0 -1 9968
box -3552 2527 26658 5446
use brbufhalf  brbufhalf_1
timestamp 1656715967
transform 1 0 33754 0 1 -2528
box -3552 2527 26658 5446
use brbufhalf  brbufhalf_2
timestamp 1656715967
transform 1 0 3552 0 1 -2528
box -3552 2527 26658 5446
use brbufhalf_128  brbufhalf_128_0
timestamp 1656715967
transform -1 0 56430 0 -1 9968
box -3546 2527 26658 5446
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0
timestamp 1656715967
transform 1 0 15169 0 1 3195
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1656715967
transform 1 0 13239 0 1 3195
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_2
timestamp 1656715967
transform 1 0 45311 0 1 3355
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_3
timestamp 1656715967
transform 1 0 43381 0 1 3355
box -38 -48 1510 592
<< properties >>
string GDS_END 9659582
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/design_merged.gds
string GDS_START 9627558
<< end >>
