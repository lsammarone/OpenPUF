magic
tech sky130A
magscale 1 2
timestamp 1655323538
<< metal3 >>
rect -1052 152 1051 180
rect -1052 -152 -1032 152
rect 1032 -152 1051 152
rect -1052 -180 1051 -152
<< via3 >>
rect -1032 -152 1032 152
<< metal4 >>
rect -1052 152 1051 180
rect -1052 -152 -1032 152
rect 1032 -152 1051 152
rect -1052 -180 1051 -152
<< end >>
