magic
tech sky130A
magscale 1 2
timestamp 1655322987
<< metal4 >>
rect -403 598 403 720
rect -403 -598 -278 598
rect 278 -598 403 598
rect -403 -721 403 -598
<< via4 >>
rect -278 -598 278 598
<< metal5 >>
rect -403 598 403 720
rect -403 -598 -278 598
rect 278 -598 403 598
rect -403 -721 403 -598
<< end >>
