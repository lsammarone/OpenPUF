magic
tech sky130A
magscale 1 2
timestamp 1656715967
<< metal1 >>
rect -500 500 500 557
rect -500 -557 500 -500
<< rmetal1 >>
rect -500 -500 500 500
<< properties >>
string gencell sky130_fd_pr__res_generic_m1
string library sky130
string parameters w 5 l 5 m 1 nx 1 wmin 0.14 lmin 0.14 rho 0.125 val 125.0m dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
