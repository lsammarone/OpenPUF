magic
tech sky130A
magscale 1 2
timestamp 1656729169
<< pwell >>
rect -2704 526 2602 602
rect -2704 -526 2635 526
rect -2704 -996 2602 -526
<< nmoslvt >>
rect -2551 -500 -2351 500
rect -2293 -500 -2093 500
rect -2035 -500 -1835 500
rect -1777 -500 -1577 500
rect -1519 -500 -1319 500
rect -1261 -500 -1061 500
rect -1003 -500 -803 500
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
rect 803 -500 1003 500
rect 1061 -500 1261 500
rect 1319 -500 1519 500
rect 1577 -500 1777 500
rect 1835 -500 2035 500
rect 2093 -500 2293 500
rect 2351 -500 2551 500
<< ndiff >>
rect -2609 459 -2551 500
rect -2609 425 -2597 459
rect -2563 425 -2551 459
rect -2609 391 -2551 425
rect -2609 357 -2597 391
rect -2563 357 -2551 391
rect -2609 323 -2551 357
rect -2609 289 -2597 323
rect -2563 289 -2551 323
rect -2609 255 -2551 289
rect -2609 221 -2597 255
rect -2563 221 -2551 255
rect -2609 187 -2551 221
rect -2609 153 -2597 187
rect -2563 153 -2551 187
rect -2609 119 -2551 153
rect -2609 85 -2597 119
rect -2563 85 -2551 119
rect -2609 51 -2551 85
rect -2609 17 -2597 51
rect -2563 17 -2551 51
rect -2609 -17 -2551 17
rect -2609 -51 -2597 -17
rect -2563 -51 -2551 -17
rect -2609 -85 -2551 -51
rect -2609 -119 -2597 -85
rect -2563 -119 -2551 -85
rect -2609 -153 -2551 -119
rect -2609 -187 -2597 -153
rect -2563 -187 -2551 -153
rect -2609 -221 -2551 -187
rect -2609 -255 -2597 -221
rect -2563 -255 -2551 -221
rect -2609 -289 -2551 -255
rect -2609 -323 -2597 -289
rect -2563 -323 -2551 -289
rect -2609 -357 -2551 -323
rect -2609 -391 -2597 -357
rect -2563 -391 -2551 -357
rect -2609 -425 -2551 -391
rect -2609 -459 -2597 -425
rect -2563 -459 -2551 -425
rect -2609 -500 -2551 -459
rect -2351 459 -2293 500
rect -2351 425 -2339 459
rect -2305 425 -2293 459
rect -2351 391 -2293 425
rect -2351 357 -2339 391
rect -2305 357 -2293 391
rect -2351 323 -2293 357
rect -2351 289 -2339 323
rect -2305 289 -2293 323
rect -2351 255 -2293 289
rect -2351 221 -2339 255
rect -2305 221 -2293 255
rect -2351 187 -2293 221
rect -2351 153 -2339 187
rect -2305 153 -2293 187
rect -2351 119 -2293 153
rect -2351 85 -2339 119
rect -2305 85 -2293 119
rect -2351 51 -2293 85
rect -2351 17 -2339 51
rect -2305 17 -2293 51
rect -2351 -17 -2293 17
rect -2351 -51 -2339 -17
rect -2305 -51 -2293 -17
rect -2351 -85 -2293 -51
rect -2351 -119 -2339 -85
rect -2305 -119 -2293 -85
rect -2351 -153 -2293 -119
rect -2351 -187 -2339 -153
rect -2305 -187 -2293 -153
rect -2351 -221 -2293 -187
rect -2351 -255 -2339 -221
rect -2305 -255 -2293 -221
rect -2351 -289 -2293 -255
rect -2351 -323 -2339 -289
rect -2305 -323 -2293 -289
rect -2351 -357 -2293 -323
rect -2351 -391 -2339 -357
rect -2305 -391 -2293 -357
rect -2351 -425 -2293 -391
rect -2351 -459 -2339 -425
rect -2305 -459 -2293 -425
rect -2351 -500 -2293 -459
rect -2093 459 -2035 500
rect -2093 425 -2081 459
rect -2047 425 -2035 459
rect -2093 391 -2035 425
rect -2093 357 -2081 391
rect -2047 357 -2035 391
rect -2093 323 -2035 357
rect -2093 289 -2081 323
rect -2047 289 -2035 323
rect -2093 255 -2035 289
rect -2093 221 -2081 255
rect -2047 221 -2035 255
rect -2093 187 -2035 221
rect -2093 153 -2081 187
rect -2047 153 -2035 187
rect -2093 119 -2035 153
rect -2093 85 -2081 119
rect -2047 85 -2035 119
rect -2093 51 -2035 85
rect -2093 17 -2081 51
rect -2047 17 -2035 51
rect -2093 -17 -2035 17
rect -2093 -51 -2081 -17
rect -2047 -51 -2035 -17
rect -2093 -85 -2035 -51
rect -2093 -119 -2081 -85
rect -2047 -119 -2035 -85
rect -2093 -153 -2035 -119
rect -2093 -187 -2081 -153
rect -2047 -187 -2035 -153
rect -2093 -221 -2035 -187
rect -2093 -255 -2081 -221
rect -2047 -255 -2035 -221
rect -2093 -289 -2035 -255
rect -2093 -323 -2081 -289
rect -2047 -323 -2035 -289
rect -2093 -357 -2035 -323
rect -2093 -391 -2081 -357
rect -2047 -391 -2035 -357
rect -2093 -425 -2035 -391
rect -2093 -459 -2081 -425
rect -2047 -459 -2035 -425
rect -2093 -500 -2035 -459
rect -1835 459 -1777 500
rect -1835 425 -1823 459
rect -1789 425 -1777 459
rect -1835 391 -1777 425
rect -1835 357 -1823 391
rect -1789 357 -1777 391
rect -1835 323 -1777 357
rect -1835 289 -1823 323
rect -1789 289 -1777 323
rect -1835 255 -1777 289
rect -1835 221 -1823 255
rect -1789 221 -1777 255
rect -1835 187 -1777 221
rect -1835 153 -1823 187
rect -1789 153 -1777 187
rect -1835 119 -1777 153
rect -1835 85 -1823 119
rect -1789 85 -1777 119
rect -1835 51 -1777 85
rect -1835 17 -1823 51
rect -1789 17 -1777 51
rect -1835 -17 -1777 17
rect -1835 -51 -1823 -17
rect -1789 -51 -1777 -17
rect -1835 -85 -1777 -51
rect -1835 -119 -1823 -85
rect -1789 -119 -1777 -85
rect -1835 -153 -1777 -119
rect -1835 -187 -1823 -153
rect -1789 -187 -1777 -153
rect -1835 -221 -1777 -187
rect -1835 -255 -1823 -221
rect -1789 -255 -1777 -221
rect -1835 -289 -1777 -255
rect -1835 -323 -1823 -289
rect -1789 -323 -1777 -289
rect -1835 -357 -1777 -323
rect -1835 -391 -1823 -357
rect -1789 -391 -1777 -357
rect -1835 -425 -1777 -391
rect -1835 -459 -1823 -425
rect -1789 -459 -1777 -425
rect -1835 -500 -1777 -459
rect -1577 459 -1519 500
rect -1577 425 -1565 459
rect -1531 425 -1519 459
rect -1577 391 -1519 425
rect -1577 357 -1565 391
rect -1531 357 -1519 391
rect -1577 323 -1519 357
rect -1577 289 -1565 323
rect -1531 289 -1519 323
rect -1577 255 -1519 289
rect -1577 221 -1565 255
rect -1531 221 -1519 255
rect -1577 187 -1519 221
rect -1577 153 -1565 187
rect -1531 153 -1519 187
rect -1577 119 -1519 153
rect -1577 85 -1565 119
rect -1531 85 -1519 119
rect -1577 51 -1519 85
rect -1577 17 -1565 51
rect -1531 17 -1519 51
rect -1577 -17 -1519 17
rect -1577 -51 -1565 -17
rect -1531 -51 -1519 -17
rect -1577 -85 -1519 -51
rect -1577 -119 -1565 -85
rect -1531 -119 -1519 -85
rect -1577 -153 -1519 -119
rect -1577 -187 -1565 -153
rect -1531 -187 -1519 -153
rect -1577 -221 -1519 -187
rect -1577 -255 -1565 -221
rect -1531 -255 -1519 -221
rect -1577 -289 -1519 -255
rect -1577 -323 -1565 -289
rect -1531 -323 -1519 -289
rect -1577 -357 -1519 -323
rect -1577 -391 -1565 -357
rect -1531 -391 -1519 -357
rect -1577 -425 -1519 -391
rect -1577 -459 -1565 -425
rect -1531 -459 -1519 -425
rect -1577 -500 -1519 -459
rect -1319 459 -1261 500
rect -1319 425 -1307 459
rect -1273 425 -1261 459
rect -1319 391 -1261 425
rect -1319 357 -1307 391
rect -1273 357 -1261 391
rect -1319 323 -1261 357
rect -1319 289 -1307 323
rect -1273 289 -1261 323
rect -1319 255 -1261 289
rect -1319 221 -1307 255
rect -1273 221 -1261 255
rect -1319 187 -1261 221
rect -1319 153 -1307 187
rect -1273 153 -1261 187
rect -1319 119 -1261 153
rect -1319 85 -1307 119
rect -1273 85 -1261 119
rect -1319 51 -1261 85
rect -1319 17 -1307 51
rect -1273 17 -1261 51
rect -1319 -17 -1261 17
rect -1319 -51 -1307 -17
rect -1273 -51 -1261 -17
rect -1319 -85 -1261 -51
rect -1319 -119 -1307 -85
rect -1273 -119 -1261 -85
rect -1319 -153 -1261 -119
rect -1319 -187 -1307 -153
rect -1273 -187 -1261 -153
rect -1319 -221 -1261 -187
rect -1319 -255 -1307 -221
rect -1273 -255 -1261 -221
rect -1319 -289 -1261 -255
rect -1319 -323 -1307 -289
rect -1273 -323 -1261 -289
rect -1319 -357 -1261 -323
rect -1319 -391 -1307 -357
rect -1273 -391 -1261 -357
rect -1319 -425 -1261 -391
rect -1319 -459 -1307 -425
rect -1273 -459 -1261 -425
rect -1319 -500 -1261 -459
rect -1061 459 -1003 500
rect -1061 425 -1049 459
rect -1015 425 -1003 459
rect -1061 391 -1003 425
rect -1061 357 -1049 391
rect -1015 357 -1003 391
rect -1061 323 -1003 357
rect -1061 289 -1049 323
rect -1015 289 -1003 323
rect -1061 255 -1003 289
rect -1061 221 -1049 255
rect -1015 221 -1003 255
rect -1061 187 -1003 221
rect -1061 153 -1049 187
rect -1015 153 -1003 187
rect -1061 119 -1003 153
rect -1061 85 -1049 119
rect -1015 85 -1003 119
rect -1061 51 -1003 85
rect -1061 17 -1049 51
rect -1015 17 -1003 51
rect -1061 -17 -1003 17
rect -1061 -51 -1049 -17
rect -1015 -51 -1003 -17
rect -1061 -85 -1003 -51
rect -1061 -119 -1049 -85
rect -1015 -119 -1003 -85
rect -1061 -153 -1003 -119
rect -1061 -187 -1049 -153
rect -1015 -187 -1003 -153
rect -1061 -221 -1003 -187
rect -1061 -255 -1049 -221
rect -1015 -255 -1003 -221
rect -1061 -289 -1003 -255
rect -1061 -323 -1049 -289
rect -1015 -323 -1003 -289
rect -1061 -357 -1003 -323
rect -1061 -391 -1049 -357
rect -1015 -391 -1003 -357
rect -1061 -425 -1003 -391
rect -1061 -459 -1049 -425
rect -1015 -459 -1003 -425
rect -1061 -500 -1003 -459
rect -803 459 -745 500
rect -803 425 -791 459
rect -757 425 -745 459
rect -803 391 -745 425
rect -803 357 -791 391
rect -757 357 -745 391
rect -803 323 -745 357
rect -803 289 -791 323
rect -757 289 -745 323
rect -803 255 -745 289
rect -803 221 -791 255
rect -757 221 -745 255
rect -803 187 -745 221
rect -803 153 -791 187
rect -757 153 -745 187
rect -803 119 -745 153
rect -803 85 -791 119
rect -757 85 -745 119
rect -803 51 -745 85
rect -803 17 -791 51
rect -757 17 -745 51
rect -803 -17 -745 17
rect -803 -51 -791 -17
rect -757 -51 -745 -17
rect -803 -85 -745 -51
rect -803 -119 -791 -85
rect -757 -119 -745 -85
rect -803 -153 -745 -119
rect -803 -187 -791 -153
rect -757 -187 -745 -153
rect -803 -221 -745 -187
rect -803 -255 -791 -221
rect -757 -255 -745 -221
rect -803 -289 -745 -255
rect -803 -323 -791 -289
rect -757 -323 -745 -289
rect -803 -357 -745 -323
rect -803 -391 -791 -357
rect -757 -391 -745 -357
rect -803 -425 -745 -391
rect -803 -459 -791 -425
rect -757 -459 -745 -425
rect -803 -500 -745 -459
rect -545 459 -487 500
rect -545 425 -533 459
rect -499 425 -487 459
rect -545 391 -487 425
rect -545 357 -533 391
rect -499 357 -487 391
rect -545 323 -487 357
rect -545 289 -533 323
rect -499 289 -487 323
rect -545 255 -487 289
rect -545 221 -533 255
rect -499 221 -487 255
rect -545 187 -487 221
rect -545 153 -533 187
rect -499 153 -487 187
rect -545 119 -487 153
rect -545 85 -533 119
rect -499 85 -487 119
rect -545 51 -487 85
rect -545 17 -533 51
rect -499 17 -487 51
rect -545 -17 -487 17
rect -545 -51 -533 -17
rect -499 -51 -487 -17
rect -545 -85 -487 -51
rect -545 -119 -533 -85
rect -499 -119 -487 -85
rect -545 -153 -487 -119
rect -545 -187 -533 -153
rect -499 -187 -487 -153
rect -545 -221 -487 -187
rect -545 -255 -533 -221
rect -499 -255 -487 -221
rect -545 -289 -487 -255
rect -545 -323 -533 -289
rect -499 -323 -487 -289
rect -545 -357 -487 -323
rect -545 -391 -533 -357
rect -499 -391 -487 -357
rect -545 -425 -487 -391
rect -545 -459 -533 -425
rect -499 -459 -487 -425
rect -545 -500 -487 -459
rect -287 459 -229 500
rect -287 425 -275 459
rect -241 425 -229 459
rect -287 391 -229 425
rect -287 357 -275 391
rect -241 357 -229 391
rect -287 323 -229 357
rect -287 289 -275 323
rect -241 289 -229 323
rect -287 255 -229 289
rect -287 221 -275 255
rect -241 221 -229 255
rect -287 187 -229 221
rect -287 153 -275 187
rect -241 153 -229 187
rect -287 119 -229 153
rect -287 85 -275 119
rect -241 85 -229 119
rect -287 51 -229 85
rect -287 17 -275 51
rect -241 17 -229 51
rect -287 -17 -229 17
rect -287 -51 -275 -17
rect -241 -51 -229 -17
rect -287 -85 -229 -51
rect -287 -119 -275 -85
rect -241 -119 -229 -85
rect -287 -153 -229 -119
rect -287 -187 -275 -153
rect -241 -187 -229 -153
rect -287 -221 -229 -187
rect -287 -255 -275 -221
rect -241 -255 -229 -221
rect -287 -289 -229 -255
rect -287 -323 -275 -289
rect -241 -323 -229 -289
rect -287 -357 -229 -323
rect -287 -391 -275 -357
rect -241 -391 -229 -357
rect -287 -425 -229 -391
rect -287 -459 -275 -425
rect -241 -459 -229 -425
rect -287 -500 -229 -459
rect -29 459 29 500
rect -29 425 -17 459
rect 17 425 29 459
rect -29 391 29 425
rect -29 357 -17 391
rect 17 357 29 391
rect -29 323 29 357
rect -29 289 -17 323
rect 17 289 29 323
rect -29 255 29 289
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -289 29 -255
rect -29 -323 -17 -289
rect 17 -323 29 -289
rect -29 -357 29 -323
rect -29 -391 -17 -357
rect 17 -391 29 -357
rect -29 -425 29 -391
rect -29 -459 -17 -425
rect 17 -459 29 -425
rect -29 -500 29 -459
rect 229 459 287 500
rect 229 425 241 459
rect 275 425 287 459
rect 229 391 287 425
rect 229 357 241 391
rect 275 357 287 391
rect 229 323 287 357
rect 229 289 241 323
rect 275 289 287 323
rect 229 255 287 289
rect 229 221 241 255
rect 275 221 287 255
rect 229 187 287 221
rect 229 153 241 187
rect 275 153 287 187
rect 229 119 287 153
rect 229 85 241 119
rect 275 85 287 119
rect 229 51 287 85
rect 229 17 241 51
rect 275 17 287 51
rect 229 -17 287 17
rect 229 -51 241 -17
rect 275 -51 287 -17
rect 229 -85 287 -51
rect 229 -119 241 -85
rect 275 -119 287 -85
rect 229 -153 287 -119
rect 229 -187 241 -153
rect 275 -187 287 -153
rect 229 -221 287 -187
rect 229 -255 241 -221
rect 275 -255 287 -221
rect 229 -289 287 -255
rect 229 -323 241 -289
rect 275 -323 287 -289
rect 229 -357 287 -323
rect 229 -391 241 -357
rect 275 -391 287 -357
rect 229 -425 287 -391
rect 229 -459 241 -425
rect 275 -459 287 -425
rect 229 -500 287 -459
rect 487 459 545 500
rect 487 425 499 459
rect 533 425 545 459
rect 487 391 545 425
rect 487 357 499 391
rect 533 357 545 391
rect 487 323 545 357
rect 487 289 499 323
rect 533 289 545 323
rect 487 255 545 289
rect 487 221 499 255
rect 533 221 545 255
rect 487 187 545 221
rect 487 153 499 187
rect 533 153 545 187
rect 487 119 545 153
rect 487 85 499 119
rect 533 85 545 119
rect 487 51 545 85
rect 487 17 499 51
rect 533 17 545 51
rect 487 -17 545 17
rect 487 -51 499 -17
rect 533 -51 545 -17
rect 487 -85 545 -51
rect 487 -119 499 -85
rect 533 -119 545 -85
rect 487 -153 545 -119
rect 487 -187 499 -153
rect 533 -187 545 -153
rect 487 -221 545 -187
rect 487 -255 499 -221
rect 533 -255 545 -221
rect 487 -289 545 -255
rect 487 -323 499 -289
rect 533 -323 545 -289
rect 487 -357 545 -323
rect 487 -391 499 -357
rect 533 -391 545 -357
rect 487 -425 545 -391
rect 487 -459 499 -425
rect 533 -459 545 -425
rect 487 -500 545 -459
rect 745 459 803 500
rect 745 425 757 459
rect 791 425 803 459
rect 745 391 803 425
rect 745 357 757 391
rect 791 357 803 391
rect 745 323 803 357
rect 745 289 757 323
rect 791 289 803 323
rect 745 255 803 289
rect 745 221 757 255
rect 791 221 803 255
rect 745 187 803 221
rect 745 153 757 187
rect 791 153 803 187
rect 745 119 803 153
rect 745 85 757 119
rect 791 85 803 119
rect 745 51 803 85
rect 745 17 757 51
rect 791 17 803 51
rect 745 -17 803 17
rect 745 -51 757 -17
rect 791 -51 803 -17
rect 745 -85 803 -51
rect 745 -119 757 -85
rect 791 -119 803 -85
rect 745 -153 803 -119
rect 745 -187 757 -153
rect 791 -187 803 -153
rect 745 -221 803 -187
rect 745 -255 757 -221
rect 791 -255 803 -221
rect 745 -289 803 -255
rect 745 -323 757 -289
rect 791 -323 803 -289
rect 745 -357 803 -323
rect 745 -391 757 -357
rect 791 -391 803 -357
rect 745 -425 803 -391
rect 745 -459 757 -425
rect 791 -459 803 -425
rect 745 -500 803 -459
rect 1003 459 1061 500
rect 1003 425 1015 459
rect 1049 425 1061 459
rect 1003 391 1061 425
rect 1003 357 1015 391
rect 1049 357 1061 391
rect 1003 323 1061 357
rect 1003 289 1015 323
rect 1049 289 1061 323
rect 1003 255 1061 289
rect 1003 221 1015 255
rect 1049 221 1061 255
rect 1003 187 1061 221
rect 1003 153 1015 187
rect 1049 153 1061 187
rect 1003 119 1061 153
rect 1003 85 1015 119
rect 1049 85 1061 119
rect 1003 51 1061 85
rect 1003 17 1015 51
rect 1049 17 1061 51
rect 1003 -17 1061 17
rect 1003 -51 1015 -17
rect 1049 -51 1061 -17
rect 1003 -85 1061 -51
rect 1003 -119 1015 -85
rect 1049 -119 1061 -85
rect 1003 -153 1061 -119
rect 1003 -187 1015 -153
rect 1049 -187 1061 -153
rect 1003 -221 1061 -187
rect 1003 -255 1015 -221
rect 1049 -255 1061 -221
rect 1003 -289 1061 -255
rect 1003 -323 1015 -289
rect 1049 -323 1061 -289
rect 1003 -357 1061 -323
rect 1003 -391 1015 -357
rect 1049 -391 1061 -357
rect 1003 -425 1061 -391
rect 1003 -459 1015 -425
rect 1049 -459 1061 -425
rect 1003 -500 1061 -459
rect 1261 459 1319 500
rect 1261 425 1273 459
rect 1307 425 1319 459
rect 1261 391 1319 425
rect 1261 357 1273 391
rect 1307 357 1319 391
rect 1261 323 1319 357
rect 1261 289 1273 323
rect 1307 289 1319 323
rect 1261 255 1319 289
rect 1261 221 1273 255
rect 1307 221 1319 255
rect 1261 187 1319 221
rect 1261 153 1273 187
rect 1307 153 1319 187
rect 1261 119 1319 153
rect 1261 85 1273 119
rect 1307 85 1319 119
rect 1261 51 1319 85
rect 1261 17 1273 51
rect 1307 17 1319 51
rect 1261 -17 1319 17
rect 1261 -51 1273 -17
rect 1307 -51 1319 -17
rect 1261 -85 1319 -51
rect 1261 -119 1273 -85
rect 1307 -119 1319 -85
rect 1261 -153 1319 -119
rect 1261 -187 1273 -153
rect 1307 -187 1319 -153
rect 1261 -221 1319 -187
rect 1261 -255 1273 -221
rect 1307 -255 1319 -221
rect 1261 -289 1319 -255
rect 1261 -323 1273 -289
rect 1307 -323 1319 -289
rect 1261 -357 1319 -323
rect 1261 -391 1273 -357
rect 1307 -391 1319 -357
rect 1261 -425 1319 -391
rect 1261 -459 1273 -425
rect 1307 -459 1319 -425
rect 1261 -500 1319 -459
rect 1519 459 1577 500
rect 1519 425 1531 459
rect 1565 425 1577 459
rect 1519 391 1577 425
rect 1519 357 1531 391
rect 1565 357 1577 391
rect 1519 323 1577 357
rect 1519 289 1531 323
rect 1565 289 1577 323
rect 1519 255 1577 289
rect 1519 221 1531 255
rect 1565 221 1577 255
rect 1519 187 1577 221
rect 1519 153 1531 187
rect 1565 153 1577 187
rect 1519 119 1577 153
rect 1519 85 1531 119
rect 1565 85 1577 119
rect 1519 51 1577 85
rect 1519 17 1531 51
rect 1565 17 1577 51
rect 1519 -17 1577 17
rect 1519 -51 1531 -17
rect 1565 -51 1577 -17
rect 1519 -85 1577 -51
rect 1519 -119 1531 -85
rect 1565 -119 1577 -85
rect 1519 -153 1577 -119
rect 1519 -187 1531 -153
rect 1565 -187 1577 -153
rect 1519 -221 1577 -187
rect 1519 -255 1531 -221
rect 1565 -255 1577 -221
rect 1519 -289 1577 -255
rect 1519 -323 1531 -289
rect 1565 -323 1577 -289
rect 1519 -357 1577 -323
rect 1519 -391 1531 -357
rect 1565 -391 1577 -357
rect 1519 -425 1577 -391
rect 1519 -459 1531 -425
rect 1565 -459 1577 -425
rect 1519 -500 1577 -459
rect 1777 459 1835 500
rect 1777 425 1789 459
rect 1823 425 1835 459
rect 1777 391 1835 425
rect 1777 357 1789 391
rect 1823 357 1835 391
rect 1777 323 1835 357
rect 1777 289 1789 323
rect 1823 289 1835 323
rect 1777 255 1835 289
rect 1777 221 1789 255
rect 1823 221 1835 255
rect 1777 187 1835 221
rect 1777 153 1789 187
rect 1823 153 1835 187
rect 1777 119 1835 153
rect 1777 85 1789 119
rect 1823 85 1835 119
rect 1777 51 1835 85
rect 1777 17 1789 51
rect 1823 17 1835 51
rect 1777 -17 1835 17
rect 1777 -51 1789 -17
rect 1823 -51 1835 -17
rect 1777 -85 1835 -51
rect 1777 -119 1789 -85
rect 1823 -119 1835 -85
rect 1777 -153 1835 -119
rect 1777 -187 1789 -153
rect 1823 -187 1835 -153
rect 1777 -221 1835 -187
rect 1777 -255 1789 -221
rect 1823 -255 1835 -221
rect 1777 -289 1835 -255
rect 1777 -323 1789 -289
rect 1823 -323 1835 -289
rect 1777 -357 1835 -323
rect 1777 -391 1789 -357
rect 1823 -391 1835 -357
rect 1777 -425 1835 -391
rect 1777 -459 1789 -425
rect 1823 -459 1835 -425
rect 1777 -500 1835 -459
rect 2035 459 2093 500
rect 2035 425 2047 459
rect 2081 425 2093 459
rect 2035 391 2093 425
rect 2035 357 2047 391
rect 2081 357 2093 391
rect 2035 323 2093 357
rect 2035 289 2047 323
rect 2081 289 2093 323
rect 2035 255 2093 289
rect 2035 221 2047 255
rect 2081 221 2093 255
rect 2035 187 2093 221
rect 2035 153 2047 187
rect 2081 153 2093 187
rect 2035 119 2093 153
rect 2035 85 2047 119
rect 2081 85 2093 119
rect 2035 51 2093 85
rect 2035 17 2047 51
rect 2081 17 2093 51
rect 2035 -17 2093 17
rect 2035 -51 2047 -17
rect 2081 -51 2093 -17
rect 2035 -85 2093 -51
rect 2035 -119 2047 -85
rect 2081 -119 2093 -85
rect 2035 -153 2093 -119
rect 2035 -187 2047 -153
rect 2081 -187 2093 -153
rect 2035 -221 2093 -187
rect 2035 -255 2047 -221
rect 2081 -255 2093 -221
rect 2035 -289 2093 -255
rect 2035 -323 2047 -289
rect 2081 -323 2093 -289
rect 2035 -357 2093 -323
rect 2035 -391 2047 -357
rect 2081 -391 2093 -357
rect 2035 -425 2093 -391
rect 2035 -459 2047 -425
rect 2081 -459 2093 -425
rect 2035 -500 2093 -459
rect 2293 459 2351 500
rect 2293 425 2305 459
rect 2339 425 2351 459
rect 2293 391 2351 425
rect 2293 357 2305 391
rect 2339 357 2351 391
rect 2293 323 2351 357
rect 2293 289 2305 323
rect 2339 289 2351 323
rect 2293 255 2351 289
rect 2293 221 2305 255
rect 2339 221 2351 255
rect 2293 187 2351 221
rect 2293 153 2305 187
rect 2339 153 2351 187
rect 2293 119 2351 153
rect 2293 85 2305 119
rect 2339 85 2351 119
rect 2293 51 2351 85
rect 2293 17 2305 51
rect 2339 17 2351 51
rect 2293 -17 2351 17
rect 2293 -51 2305 -17
rect 2339 -51 2351 -17
rect 2293 -85 2351 -51
rect 2293 -119 2305 -85
rect 2339 -119 2351 -85
rect 2293 -153 2351 -119
rect 2293 -187 2305 -153
rect 2339 -187 2351 -153
rect 2293 -221 2351 -187
rect 2293 -255 2305 -221
rect 2339 -255 2351 -221
rect 2293 -289 2351 -255
rect 2293 -323 2305 -289
rect 2339 -323 2351 -289
rect 2293 -357 2351 -323
rect 2293 -391 2305 -357
rect 2339 -391 2351 -357
rect 2293 -425 2351 -391
rect 2293 -459 2305 -425
rect 2339 -459 2351 -425
rect 2293 -500 2351 -459
rect 2551 459 2609 500
rect 2551 425 2563 459
rect 2597 425 2609 459
rect 2551 391 2609 425
rect 2551 357 2563 391
rect 2597 357 2609 391
rect 2551 323 2609 357
rect 2551 289 2563 323
rect 2597 289 2609 323
rect 2551 255 2609 289
rect 2551 221 2563 255
rect 2597 221 2609 255
rect 2551 187 2609 221
rect 2551 153 2563 187
rect 2597 153 2609 187
rect 2551 119 2609 153
rect 2551 85 2563 119
rect 2597 85 2609 119
rect 2551 51 2609 85
rect 2551 17 2563 51
rect 2597 17 2609 51
rect 2551 -17 2609 17
rect 2551 -51 2563 -17
rect 2597 -51 2609 -17
rect 2551 -85 2609 -51
rect 2551 -119 2563 -85
rect 2597 -119 2609 -85
rect 2551 -153 2609 -119
rect 2551 -187 2563 -153
rect 2597 -187 2609 -153
rect 2551 -221 2609 -187
rect 2551 -255 2563 -221
rect 2597 -255 2609 -221
rect 2551 -289 2609 -255
rect 2551 -323 2563 -289
rect 2597 -323 2609 -289
rect 2551 -357 2609 -323
rect 2551 -391 2563 -357
rect 2597 -391 2609 -357
rect 2551 -425 2609 -391
rect 2551 -459 2563 -425
rect 2597 -459 2609 -425
rect 2551 -500 2609 -459
<< ndiffc >>
rect -2597 425 -2563 459
rect -2597 357 -2563 391
rect -2597 289 -2563 323
rect -2597 221 -2563 255
rect -2597 153 -2563 187
rect -2597 85 -2563 119
rect -2597 17 -2563 51
rect -2597 -51 -2563 -17
rect -2597 -119 -2563 -85
rect -2597 -187 -2563 -153
rect -2597 -255 -2563 -221
rect -2597 -323 -2563 -289
rect -2597 -391 -2563 -357
rect -2597 -459 -2563 -425
rect -2339 425 -2305 459
rect -2339 357 -2305 391
rect -2339 289 -2305 323
rect -2339 221 -2305 255
rect -2339 153 -2305 187
rect -2339 85 -2305 119
rect -2339 17 -2305 51
rect -2339 -51 -2305 -17
rect -2339 -119 -2305 -85
rect -2339 -187 -2305 -153
rect -2339 -255 -2305 -221
rect -2339 -323 -2305 -289
rect -2339 -391 -2305 -357
rect -2339 -459 -2305 -425
rect -2081 425 -2047 459
rect -2081 357 -2047 391
rect -2081 289 -2047 323
rect -2081 221 -2047 255
rect -2081 153 -2047 187
rect -2081 85 -2047 119
rect -2081 17 -2047 51
rect -2081 -51 -2047 -17
rect -2081 -119 -2047 -85
rect -2081 -187 -2047 -153
rect -2081 -255 -2047 -221
rect -2081 -323 -2047 -289
rect -2081 -391 -2047 -357
rect -2081 -459 -2047 -425
rect -1823 425 -1789 459
rect -1823 357 -1789 391
rect -1823 289 -1789 323
rect -1823 221 -1789 255
rect -1823 153 -1789 187
rect -1823 85 -1789 119
rect -1823 17 -1789 51
rect -1823 -51 -1789 -17
rect -1823 -119 -1789 -85
rect -1823 -187 -1789 -153
rect -1823 -255 -1789 -221
rect -1823 -323 -1789 -289
rect -1823 -391 -1789 -357
rect -1823 -459 -1789 -425
rect -1565 425 -1531 459
rect -1565 357 -1531 391
rect -1565 289 -1531 323
rect -1565 221 -1531 255
rect -1565 153 -1531 187
rect -1565 85 -1531 119
rect -1565 17 -1531 51
rect -1565 -51 -1531 -17
rect -1565 -119 -1531 -85
rect -1565 -187 -1531 -153
rect -1565 -255 -1531 -221
rect -1565 -323 -1531 -289
rect -1565 -391 -1531 -357
rect -1565 -459 -1531 -425
rect -1307 425 -1273 459
rect -1307 357 -1273 391
rect -1307 289 -1273 323
rect -1307 221 -1273 255
rect -1307 153 -1273 187
rect -1307 85 -1273 119
rect -1307 17 -1273 51
rect -1307 -51 -1273 -17
rect -1307 -119 -1273 -85
rect -1307 -187 -1273 -153
rect -1307 -255 -1273 -221
rect -1307 -323 -1273 -289
rect -1307 -391 -1273 -357
rect -1307 -459 -1273 -425
rect -1049 425 -1015 459
rect -1049 357 -1015 391
rect -1049 289 -1015 323
rect -1049 221 -1015 255
rect -1049 153 -1015 187
rect -1049 85 -1015 119
rect -1049 17 -1015 51
rect -1049 -51 -1015 -17
rect -1049 -119 -1015 -85
rect -1049 -187 -1015 -153
rect -1049 -255 -1015 -221
rect -1049 -323 -1015 -289
rect -1049 -391 -1015 -357
rect -1049 -459 -1015 -425
rect -791 425 -757 459
rect -791 357 -757 391
rect -791 289 -757 323
rect -791 221 -757 255
rect -791 153 -757 187
rect -791 85 -757 119
rect -791 17 -757 51
rect -791 -51 -757 -17
rect -791 -119 -757 -85
rect -791 -187 -757 -153
rect -791 -255 -757 -221
rect -791 -323 -757 -289
rect -791 -391 -757 -357
rect -791 -459 -757 -425
rect -533 425 -499 459
rect -533 357 -499 391
rect -533 289 -499 323
rect -533 221 -499 255
rect -533 153 -499 187
rect -533 85 -499 119
rect -533 17 -499 51
rect -533 -51 -499 -17
rect -533 -119 -499 -85
rect -533 -187 -499 -153
rect -533 -255 -499 -221
rect -533 -323 -499 -289
rect -533 -391 -499 -357
rect -533 -459 -499 -425
rect -275 425 -241 459
rect -275 357 -241 391
rect -275 289 -241 323
rect -275 221 -241 255
rect -275 153 -241 187
rect -275 85 -241 119
rect -275 17 -241 51
rect -275 -51 -241 -17
rect -275 -119 -241 -85
rect -275 -187 -241 -153
rect -275 -255 -241 -221
rect -275 -323 -241 -289
rect -275 -391 -241 -357
rect -275 -459 -241 -425
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect 241 425 275 459
rect 241 357 275 391
rect 241 289 275 323
rect 241 221 275 255
rect 241 153 275 187
rect 241 85 275 119
rect 241 17 275 51
rect 241 -51 275 -17
rect 241 -119 275 -85
rect 241 -187 275 -153
rect 241 -255 275 -221
rect 241 -323 275 -289
rect 241 -391 275 -357
rect 241 -459 275 -425
rect 499 425 533 459
rect 499 357 533 391
rect 499 289 533 323
rect 499 221 533 255
rect 499 153 533 187
rect 499 85 533 119
rect 499 17 533 51
rect 499 -51 533 -17
rect 499 -119 533 -85
rect 499 -187 533 -153
rect 499 -255 533 -221
rect 499 -323 533 -289
rect 499 -391 533 -357
rect 499 -459 533 -425
rect 757 425 791 459
rect 757 357 791 391
rect 757 289 791 323
rect 757 221 791 255
rect 757 153 791 187
rect 757 85 791 119
rect 757 17 791 51
rect 757 -51 791 -17
rect 757 -119 791 -85
rect 757 -187 791 -153
rect 757 -255 791 -221
rect 757 -323 791 -289
rect 757 -391 791 -357
rect 757 -459 791 -425
rect 1015 425 1049 459
rect 1015 357 1049 391
rect 1015 289 1049 323
rect 1015 221 1049 255
rect 1015 153 1049 187
rect 1015 85 1049 119
rect 1015 17 1049 51
rect 1015 -51 1049 -17
rect 1015 -119 1049 -85
rect 1015 -187 1049 -153
rect 1015 -255 1049 -221
rect 1015 -323 1049 -289
rect 1015 -391 1049 -357
rect 1015 -459 1049 -425
rect 1273 425 1307 459
rect 1273 357 1307 391
rect 1273 289 1307 323
rect 1273 221 1307 255
rect 1273 153 1307 187
rect 1273 85 1307 119
rect 1273 17 1307 51
rect 1273 -51 1307 -17
rect 1273 -119 1307 -85
rect 1273 -187 1307 -153
rect 1273 -255 1307 -221
rect 1273 -323 1307 -289
rect 1273 -391 1307 -357
rect 1273 -459 1307 -425
rect 1531 425 1565 459
rect 1531 357 1565 391
rect 1531 289 1565 323
rect 1531 221 1565 255
rect 1531 153 1565 187
rect 1531 85 1565 119
rect 1531 17 1565 51
rect 1531 -51 1565 -17
rect 1531 -119 1565 -85
rect 1531 -187 1565 -153
rect 1531 -255 1565 -221
rect 1531 -323 1565 -289
rect 1531 -391 1565 -357
rect 1531 -459 1565 -425
rect 1789 425 1823 459
rect 1789 357 1823 391
rect 1789 289 1823 323
rect 1789 221 1823 255
rect 1789 153 1823 187
rect 1789 85 1823 119
rect 1789 17 1823 51
rect 1789 -51 1823 -17
rect 1789 -119 1823 -85
rect 1789 -187 1823 -153
rect 1789 -255 1823 -221
rect 1789 -323 1823 -289
rect 1789 -391 1823 -357
rect 1789 -459 1823 -425
rect 2047 425 2081 459
rect 2047 357 2081 391
rect 2047 289 2081 323
rect 2047 221 2081 255
rect 2047 153 2081 187
rect 2047 85 2081 119
rect 2047 17 2081 51
rect 2047 -51 2081 -17
rect 2047 -119 2081 -85
rect 2047 -187 2081 -153
rect 2047 -255 2081 -221
rect 2047 -323 2081 -289
rect 2047 -391 2081 -357
rect 2047 -459 2081 -425
rect 2305 425 2339 459
rect 2305 357 2339 391
rect 2305 289 2339 323
rect 2305 221 2339 255
rect 2305 153 2339 187
rect 2305 85 2339 119
rect 2305 17 2339 51
rect 2305 -51 2339 -17
rect 2305 -119 2339 -85
rect 2305 -187 2339 -153
rect 2305 -255 2339 -221
rect 2305 -323 2339 -289
rect 2305 -391 2339 -357
rect 2305 -459 2339 -425
rect 2563 425 2597 459
rect 2563 357 2597 391
rect 2563 289 2597 323
rect 2563 221 2597 255
rect 2563 153 2597 187
rect 2563 85 2597 119
rect 2563 17 2597 51
rect 2563 -51 2597 -17
rect 2563 -119 2597 -85
rect 2563 -187 2597 -153
rect 2563 -255 2597 -221
rect 2563 -323 2597 -289
rect 2563 -391 2597 -357
rect 2563 -459 2597 -425
<< psubdiff >>
rect -2668 -843 -2628 -800
rect -2668 -877 -2665 -843
rect -2631 -877 -2628 -843
rect -2668 -920 -2628 -877
rect -1610 -873 -1490 -870
rect -1610 -907 -1565 -873
rect -1531 -907 -1490 -873
rect -1610 -920 -1490 -907
rect -310 -873 -190 -870
rect -310 -907 -265 -873
rect -231 -907 -190 -873
rect -310 -920 -190 -907
rect 990 -873 1110 -870
rect 990 -907 1035 -873
rect 1069 -907 1110 -873
rect 990 -920 1110 -907
<< psubdiffcont >>
rect -2665 -877 -2631 -843
rect -1565 -907 -1531 -873
rect -265 -907 -231 -873
rect 1035 -907 1069 -873
<< poly >>
rect -2551 500 -2351 526
rect -2293 500 -2093 526
rect -2035 500 -1835 526
rect -1777 500 -1577 526
rect -1519 500 -1319 526
rect -1261 500 -1061 526
rect -1003 500 -803 526
rect -745 500 -545 526
rect -487 500 -287 526
rect -229 500 -29 526
rect 29 500 229 526
rect 287 500 487 526
rect 545 500 745 526
rect 803 500 1003 526
rect 1061 500 1261 526
rect 1319 500 1519 526
rect 1577 500 1777 526
rect 1835 500 2035 526
rect 2093 500 2293 526
rect 2351 500 2551 526
rect -2551 -526 -2351 -500
rect -2293 -526 -2093 -500
rect -2035 -526 -1835 -500
rect -1777 -526 -1577 -500
rect -1519 -526 -1319 -500
rect -1261 -526 -1061 -500
rect -1003 -526 -803 -500
rect -745 -526 -545 -500
rect -487 -526 -287 -500
rect -229 -526 -29 -500
rect 29 -526 229 -500
rect 287 -526 487 -500
rect 545 -526 745 -500
rect 803 -526 1003 -500
rect 1061 -526 1261 -500
rect 1319 -526 1519 -500
rect 1577 -526 1777 -500
rect 1835 -526 2035 -500
rect 2093 -526 2293 -500
rect 2351 -526 2551 -500
rect -2488 -716 -2368 -526
rect -2232 -716 -2112 -526
rect -1976 -716 -1856 -526
rect -1720 -716 -1600 -526
rect -1464 -716 -1344 -526
rect -1208 -716 -1088 -526
rect -952 -716 -832 -526
rect -696 -716 -576 -526
rect -440 -716 -320 -526
rect -184 -716 -64 -526
rect 72 -716 192 -526
rect 328 -716 448 -526
rect 584 -716 704 -526
rect 840 -716 960 -526
rect 1096 -716 1216 -526
rect 1352 -716 1472 -526
rect 1608 -716 1728 -526
rect 1864 -716 1984 -526
rect 2120 -716 2240 -526
rect 2376 -716 2496 -526
rect -2528 -749 2608 -716
rect -2528 -783 -2425 -749
rect -2391 -783 -2225 -749
rect -2191 -783 -2025 -749
rect -1991 -783 -1825 -749
rect -1791 -783 -1625 -749
rect -1591 -783 -1425 -749
rect -1391 -783 -1225 -749
rect -1191 -783 -1025 -749
rect -991 -783 -825 -749
rect -791 -783 -625 -749
rect -591 -783 -425 -749
rect -391 -783 -225 -749
rect -191 -783 -25 -749
rect 9 -783 175 -749
rect 209 -783 375 -749
rect 409 -783 575 -749
rect 609 -783 775 -749
rect 809 -783 975 -749
rect 1009 -783 1175 -749
rect 1209 -783 1375 -749
rect 1409 -783 1575 -749
rect 1609 -783 1775 -749
rect 1809 -783 1975 -749
rect 2009 -783 2175 -749
rect 2209 -783 2375 -749
rect 2409 -783 2608 -749
rect -2528 -816 2608 -783
<< polycont >>
rect -2425 -783 -2391 -749
rect -2225 -783 -2191 -749
rect -2025 -783 -1991 -749
rect -1825 -783 -1791 -749
rect -1625 -783 -1591 -749
rect -1425 -783 -1391 -749
rect -1225 -783 -1191 -749
rect -1025 -783 -991 -749
rect -825 -783 -791 -749
rect -625 -783 -591 -749
rect -425 -783 -391 -749
rect -225 -783 -191 -749
rect -25 -783 9 -749
rect 175 -783 209 -749
rect 375 -783 409 -749
rect 575 -783 609 -749
rect 775 -783 809 -749
rect 975 -783 1009 -749
rect 1175 -783 1209 -749
rect 1375 -783 1409 -749
rect 1575 -783 1609 -749
rect 1775 -783 1809 -749
rect 1975 -783 2009 -749
rect 2175 -783 2209 -749
rect 2375 -783 2409 -749
<< locali >>
rect -2706 897 2608 910
rect -2706 863 -2425 897
rect -2391 863 -2225 897
rect -2191 863 -2025 897
rect -1991 863 -1825 897
rect -1791 863 -1625 897
rect -1591 863 -1425 897
rect -1391 863 -1225 897
rect -1191 863 -1025 897
rect -991 863 -825 897
rect -791 863 -625 897
rect -591 863 -425 897
rect -391 863 -225 897
rect -191 863 -25 897
rect 9 863 175 897
rect 209 863 375 897
rect 409 863 575 897
rect 609 863 775 897
rect 809 863 975 897
rect 1009 863 1175 897
rect 1209 863 1375 897
rect 1409 863 1575 897
rect 1609 863 1775 897
rect 1809 863 1975 897
rect 2009 863 2175 897
rect 2209 863 2375 897
rect 2409 863 2608 897
rect -2706 850 2608 863
rect -2608 690 2608 750
rect -2597 485 -2563 504
rect -2597 413 -2563 425
rect -2597 341 -2563 357
rect -2597 269 -2563 289
rect -2597 197 -2563 221
rect -2597 125 -2563 153
rect -2597 53 -2563 85
rect -2597 -17 -2563 17
rect -2597 -85 -2563 -53
rect -2597 -153 -2563 -125
rect -2597 -221 -2563 -197
rect -2597 -289 -2563 -269
rect -2597 -357 -2563 -341
rect -2597 -425 -2563 -413
rect -2597 -570 -2563 -485
rect -2339 485 -2305 690
rect -2339 413 -2305 425
rect -2339 341 -2305 357
rect -2339 269 -2305 289
rect -2339 197 -2305 221
rect -2339 125 -2305 153
rect -2339 53 -2305 85
rect -2339 -17 -2305 17
rect -2339 -85 -2305 -53
rect -2339 -153 -2305 -125
rect -2339 -221 -2305 -197
rect -2339 -289 -2305 -269
rect -2339 -357 -2305 -341
rect -2339 -425 -2305 -413
rect -2339 -504 -2305 -485
rect -2081 485 -2047 504
rect -2081 413 -2047 425
rect -2081 341 -2047 357
rect -2081 269 -2047 289
rect -2081 197 -2047 221
rect -2081 125 -2047 153
rect -2081 53 -2047 85
rect -2081 -17 -2047 17
rect -2081 -85 -2047 -53
rect -2081 -153 -2047 -125
rect -2081 -221 -2047 -197
rect -2081 -289 -2047 -269
rect -2081 -357 -2047 -341
rect -2081 -425 -2047 -413
rect -2081 -570 -2047 -485
rect -1823 485 -1789 690
rect -1823 413 -1789 425
rect -1823 341 -1789 357
rect -1823 269 -1789 289
rect -1823 197 -1789 221
rect -1823 125 -1789 153
rect -1823 53 -1789 85
rect -1823 -17 -1789 17
rect -1823 -85 -1789 -53
rect -1823 -153 -1789 -125
rect -1823 -221 -1789 -197
rect -1823 -289 -1789 -269
rect -1823 -357 -1789 -341
rect -1823 -425 -1789 -413
rect -1823 -504 -1789 -485
rect -1565 485 -1531 504
rect -1565 413 -1531 425
rect -1565 341 -1531 357
rect -1565 269 -1531 289
rect -1565 197 -1531 221
rect -1565 125 -1531 153
rect -1565 53 -1531 85
rect -1565 -17 -1531 17
rect -1565 -85 -1531 -53
rect -1565 -153 -1531 -125
rect -1565 -221 -1531 -197
rect -1565 -289 -1531 -269
rect -1565 -357 -1531 -341
rect -1565 -425 -1531 -413
rect -1565 -570 -1531 -485
rect -1307 485 -1273 690
rect -1307 413 -1273 425
rect -1307 341 -1273 357
rect -1307 269 -1273 289
rect -1307 197 -1273 221
rect -1307 125 -1273 153
rect -1307 53 -1273 85
rect -1307 -17 -1273 17
rect -1307 -85 -1273 -53
rect -1307 -153 -1273 -125
rect -1307 -221 -1273 -197
rect -1307 -289 -1273 -269
rect -1307 -357 -1273 -341
rect -1307 -425 -1273 -413
rect -1307 -504 -1273 -485
rect -1049 485 -1015 504
rect -1049 413 -1015 425
rect -1049 341 -1015 357
rect -1049 269 -1015 289
rect -1049 197 -1015 221
rect -1049 125 -1015 153
rect -1049 53 -1015 85
rect -1049 -17 -1015 17
rect -1049 -85 -1015 -53
rect -1049 -153 -1015 -125
rect -1049 -221 -1015 -197
rect -1049 -289 -1015 -269
rect -1049 -357 -1015 -341
rect -1049 -425 -1015 -413
rect -1049 -570 -1015 -485
rect -791 485 -757 690
rect -791 413 -757 425
rect -791 341 -757 357
rect -791 269 -757 289
rect -791 197 -757 221
rect -791 125 -757 153
rect -791 53 -757 85
rect -791 -17 -757 17
rect -791 -85 -757 -53
rect -791 -153 -757 -125
rect -791 -221 -757 -197
rect -791 -289 -757 -269
rect -791 -357 -757 -341
rect -791 -425 -757 -413
rect -791 -504 -757 -485
rect -533 485 -499 504
rect -533 413 -499 425
rect -533 341 -499 357
rect -533 269 -499 289
rect -533 197 -499 221
rect -533 125 -499 153
rect -533 53 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -53
rect -533 -153 -499 -125
rect -533 -221 -499 -197
rect -533 -289 -499 -269
rect -533 -357 -499 -341
rect -533 -425 -499 -413
rect -533 -570 -499 -485
rect -275 485 -241 690
rect -275 413 -241 425
rect -275 341 -241 357
rect -275 269 -241 289
rect -275 197 -241 221
rect -275 125 -241 153
rect -275 53 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -53
rect -275 -153 -241 -125
rect -275 -221 -241 -197
rect -275 -289 -241 -269
rect -275 -357 -241 -341
rect -275 -425 -241 -413
rect -275 -504 -241 -485
rect -17 485 17 504
rect -17 413 17 425
rect -17 341 17 357
rect -17 269 17 289
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -289 17 -269
rect -17 -357 17 -341
rect -17 -425 17 -413
rect -17 -570 17 -485
rect 241 485 275 690
rect 241 413 275 425
rect 241 341 275 357
rect 241 269 275 289
rect 241 197 275 221
rect 241 125 275 153
rect 241 53 275 85
rect 241 -17 275 17
rect 241 -85 275 -53
rect 241 -153 275 -125
rect 241 -221 275 -197
rect 241 -289 275 -269
rect 241 -357 275 -341
rect 241 -425 275 -413
rect 241 -504 275 -485
rect 499 485 533 504
rect 499 413 533 425
rect 499 341 533 357
rect 499 269 533 289
rect 499 197 533 221
rect 499 125 533 153
rect 499 53 533 85
rect 499 -17 533 17
rect 499 -85 533 -53
rect 499 -153 533 -125
rect 499 -221 533 -197
rect 499 -289 533 -269
rect 499 -357 533 -341
rect 499 -425 533 -413
rect 499 -570 533 -485
rect 757 485 791 690
rect 757 413 791 425
rect 757 341 791 357
rect 757 269 791 289
rect 757 197 791 221
rect 757 125 791 153
rect 757 53 791 85
rect 757 -17 791 17
rect 757 -85 791 -53
rect 757 -153 791 -125
rect 757 -221 791 -197
rect 757 -289 791 -269
rect 757 -357 791 -341
rect 757 -425 791 -413
rect 757 -504 791 -485
rect 1015 485 1049 504
rect 1015 413 1049 425
rect 1015 341 1049 357
rect 1015 269 1049 289
rect 1015 197 1049 221
rect 1015 125 1049 153
rect 1015 53 1049 85
rect 1015 -17 1049 17
rect 1015 -85 1049 -53
rect 1015 -153 1049 -125
rect 1015 -221 1049 -197
rect 1015 -289 1049 -269
rect 1015 -357 1049 -341
rect 1015 -425 1049 -413
rect 1015 -570 1049 -485
rect 1273 485 1307 690
rect 1273 413 1307 425
rect 1273 341 1307 357
rect 1273 269 1307 289
rect 1273 197 1307 221
rect 1273 125 1307 153
rect 1273 53 1307 85
rect 1273 -17 1307 17
rect 1273 -85 1307 -53
rect 1273 -153 1307 -125
rect 1273 -221 1307 -197
rect 1273 -289 1307 -269
rect 1273 -357 1307 -341
rect 1273 -425 1307 -413
rect 1273 -504 1307 -485
rect 1531 485 1565 504
rect 1531 413 1565 425
rect 1531 341 1565 357
rect 1531 269 1565 289
rect 1531 197 1565 221
rect 1531 125 1565 153
rect 1531 53 1565 85
rect 1531 -17 1565 17
rect 1531 -85 1565 -53
rect 1531 -153 1565 -125
rect 1531 -221 1565 -197
rect 1531 -289 1565 -269
rect 1531 -357 1565 -341
rect 1531 -425 1565 -413
rect 1531 -570 1565 -485
rect 1789 485 1823 690
rect 1789 413 1823 425
rect 1789 341 1823 357
rect 1789 269 1823 289
rect 1789 197 1823 221
rect 1789 125 1823 153
rect 1789 53 1823 85
rect 1789 -17 1823 17
rect 1789 -85 1823 -53
rect 1789 -153 1823 -125
rect 1789 -221 1823 -197
rect 1789 -289 1823 -269
rect 1789 -357 1823 -341
rect 1789 -425 1823 -413
rect 1789 -504 1823 -485
rect 2047 485 2081 504
rect 2047 413 2081 425
rect 2047 341 2081 357
rect 2047 269 2081 289
rect 2047 197 2081 221
rect 2047 125 2081 153
rect 2047 53 2081 85
rect 2047 -17 2081 17
rect 2047 -85 2081 -53
rect 2047 -153 2081 -125
rect 2047 -221 2081 -197
rect 2047 -289 2081 -269
rect 2047 -357 2081 -341
rect 2047 -425 2081 -413
rect 2047 -570 2081 -485
rect 2305 485 2339 690
rect 2305 413 2339 425
rect 2305 341 2339 357
rect 2305 269 2339 289
rect 2305 197 2339 221
rect 2305 125 2339 153
rect 2305 53 2339 85
rect 2305 -17 2339 17
rect 2305 -85 2339 -53
rect 2305 -153 2339 -125
rect 2305 -221 2339 -197
rect 2305 -289 2339 -269
rect 2305 -357 2339 -341
rect 2305 -425 2339 -413
rect 2305 -504 2339 -485
rect 2563 485 2597 504
rect 2563 413 2597 425
rect 2563 341 2597 357
rect 2563 269 2597 289
rect 2563 197 2597 221
rect 2563 125 2597 153
rect 2563 53 2597 85
rect 2563 -17 2597 17
rect 2563 -85 2597 -53
rect 2563 -153 2597 -125
rect 2563 -221 2597 -197
rect 2563 -289 2597 -269
rect 2563 -357 2597 -341
rect 2563 -425 2597 -413
rect 2563 -570 2597 -485
rect -2608 -630 2608 -570
rect -2528 -749 2608 -736
rect -2678 -843 -2618 -760
rect -2528 -783 -2425 -749
rect -2391 -783 -2225 -749
rect -2191 -783 -2025 -749
rect -1991 -783 -1825 -749
rect -1791 -783 -1625 -749
rect -1591 -783 -1425 -749
rect -1391 -783 -1225 -749
rect -1191 -783 -1025 -749
rect -991 -783 -825 -749
rect -791 -783 -625 -749
rect -591 -783 -425 -749
rect -391 -783 -225 -749
rect -191 -783 -25 -749
rect 9 -783 175 -749
rect 209 -783 375 -749
rect 409 -783 575 -749
rect 609 -783 775 -749
rect 809 -783 975 -749
rect 1009 -783 1175 -749
rect 1209 -783 1375 -749
rect 1409 -783 1575 -749
rect 1609 -783 1775 -749
rect 1809 -783 1975 -749
rect 2009 -783 2175 -749
rect 2209 -783 2375 -749
rect 2409 -783 2608 -749
rect -2528 -796 2608 -783
rect -2678 -877 -2665 -843
rect -2631 -877 -2618 -843
rect -2678 -970 -2618 -877
rect -1630 -873 -1470 -850
rect -1630 -907 -1565 -873
rect -1531 -907 -1470 -873
rect -1630 -970 -1470 -907
rect -330 -873 -170 -850
rect -330 -907 -265 -873
rect -231 -907 -170 -873
rect -330 -970 -170 -907
rect 970 -873 1130 -850
rect 970 -907 1035 -873
rect 1069 -907 1130 -873
rect 970 -970 1130 -907
rect -2706 -983 2608 -970
rect -2706 -1017 -2425 -983
rect -2391 -1017 -2225 -983
rect -2191 -1017 -2025 -983
rect -1991 -1017 -1825 -983
rect -1791 -1017 -1625 -983
rect -1591 -1017 -1425 -983
rect -1391 -1017 -1225 -983
rect -1191 -1017 -1025 -983
rect -991 -1017 -825 -983
rect -791 -1017 -625 -983
rect -591 -1017 -425 -983
rect -391 -1017 -225 -983
rect -191 -1017 -25 -983
rect 9 -1017 175 -983
rect 209 -1017 375 -983
rect 409 -1017 575 -983
rect 609 -1017 775 -983
rect 809 -1017 975 -983
rect 1009 -1017 1175 -983
rect 1209 -1017 1375 -983
rect 1409 -1017 1575 -983
rect 1609 -1017 1775 -983
rect 1809 -1017 1975 -983
rect 2009 -1017 2175 -983
rect 2209 -1017 2375 -983
rect 2409 -1017 2608 -983
rect -2706 -1030 2608 -1017
<< viali >>
rect -2425 863 -2391 897
rect -2225 863 -2191 897
rect -2025 863 -1991 897
rect -1825 863 -1791 897
rect -1625 863 -1591 897
rect -1425 863 -1391 897
rect -1225 863 -1191 897
rect -1025 863 -991 897
rect -825 863 -791 897
rect -625 863 -591 897
rect -425 863 -391 897
rect -225 863 -191 897
rect -25 863 9 897
rect 175 863 209 897
rect 375 863 409 897
rect 575 863 609 897
rect 775 863 809 897
rect 975 863 1009 897
rect 1175 863 1209 897
rect 1375 863 1409 897
rect 1575 863 1609 897
rect 1775 863 1809 897
rect 1975 863 2009 897
rect 2175 863 2209 897
rect 2375 863 2409 897
rect -2597 459 -2563 485
rect -2597 451 -2563 459
rect -2597 391 -2563 413
rect -2597 379 -2563 391
rect -2597 323 -2563 341
rect -2597 307 -2563 323
rect -2597 255 -2563 269
rect -2597 235 -2563 255
rect -2597 187 -2563 197
rect -2597 163 -2563 187
rect -2597 119 -2563 125
rect -2597 91 -2563 119
rect -2597 51 -2563 53
rect -2597 19 -2563 51
rect -2597 -51 -2563 -19
rect -2597 -53 -2563 -51
rect -2597 -119 -2563 -91
rect -2597 -125 -2563 -119
rect -2597 -187 -2563 -163
rect -2597 -197 -2563 -187
rect -2597 -255 -2563 -235
rect -2597 -269 -2563 -255
rect -2597 -323 -2563 -307
rect -2597 -341 -2563 -323
rect -2597 -391 -2563 -379
rect -2597 -413 -2563 -391
rect -2597 -459 -2563 -451
rect -2597 -485 -2563 -459
rect -2339 459 -2305 485
rect -2339 451 -2305 459
rect -2339 391 -2305 413
rect -2339 379 -2305 391
rect -2339 323 -2305 341
rect -2339 307 -2305 323
rect -2339 255 -2305 269
rect -2339 235 -2305 255
rect -2339 187 -2305 197
rect -2339 163 -2305 187
rect -2339 119 -2305 125
rect -2339 91 -2305 119
rect -2339 51 -2305 53
rect -2339 19 -2305 51
rect -2339 -51 -2305 -19
rect -2339 -53 -2305 -51
rect -2339 -119 -2305 -91
rect -2339 -125 -2305 -119
rect -2339 -187 -2305 -163
rect -2339 -197 -2305 -187
rect -2339 -255 -2305 -235
rect -2339 -269 -2305 -255
rect -2339 -323 -2305 -307
rect -2339 -341 -2305 -323
rect -2339 -391 -2305 -379
rect -2339 -413 -2305 -391
rect -2339 -459 -2305 -451
rect -2339 -485 -2305 -459
rect -2081 459 -2047 485
rect -2081 451 -2047 459
rect -2081 391 -2047 413
rect -2081 379 -2047 391
rect -2081 323 -2047 341
rect -2081 307 -2047 323
rect -2081 255 -2047 269
rect -2081 235 -2047 255
rect -2081 187 -2047 197
rect -2081 163 -2047 187
rect -2081 119 -2047 125
rect -2081 91 -2047 119
rect -2081 51 -2047 53
rect -2081 19 -2047 51
rect -2081 -51 -2047 -19
rect -2081 -53 -2047 -51
rect -2081 -119 -2047 -91
rect -2081 -125 -2047 -119
rect -2081 -187 -2047 -163
rect -2081 -197 -2047 -187
rect -2081 -255 -2047 -235
rect -2081 -269 -2047 -255
rect -2081 -323 -2047 -307
rect -2081 -341 -2047 -323
rect -2081 -391 -2047 -379
rect -2081 -413 -2047 -391
rect -2081 -459 -2047 -451
rect -2081 -485 -2047 -459
rect -1823 459 -1789 485
rect -1823 451 -1789 459
rect -1823 391 -1789 413
rect -1823 379 -1789 391
rect -1823 323 -1789 341
rect -1823 307 -1789 323
rect -1823 255 -1789 269
rect -1823 235 -1789 255
rect -1823 187 -1789 197
rect -1823 163 -1789 187
rect -1823 119 -1789 125
rect -1823 91 -1789 119
rect -1823 51 -1789 53
rect -1823 19 -1789 51
rect -1823 -51 -1789 -19
rect -1823 -53 -1789 -51
rect -1823 -119 -1789 -91
rect -1823 -125 -1789 -119
rect -1823 -187 -1789 -163
rect -1823 -197 -1789 -187
rect -1823 -255 -1789 -235
rect -1823 -269 -1789 -255
rect -1823 -323 -1789 -307
rect -1823 -341 -1789 -323
rect -1823 -391 -1789 -379
rect -1823 -413 -1789 -391
rect -1823 -459 -1789 -451
rect -1823 -485 -1789 -459
rect -1565 459 -1531 485
rect -1565 451 -1531 459
rect -1565 391 -1531 413
rect -1565 379 -1531 391
rect -1565 323 -1531 341
rect -1565 307 -1531 323
rect -1565 255 -1531 269
rect -1565 235 -1531 255
rect -1565 187 -1531 197
rect -1565 163 -1531 187
rect -1565 119 -1531 125
rect -1565 91 -1531 119
rect -1565 51 -1531 53
rect -1565 19 -1531 51
rect -1565 -51 -1531 -19
rect -1565 -53 -1531 -51
rect -1565 -119 -1531 -91
rect -1565 -125 -1531 -119
rect -1565 -187 -1531 -163
rect -1565 -197 -1531 -187
rect -1565 -255 -1531 -235
rect -1565 -269 -1531 -255
rect -1565 -323 -1531 -307
rect -1565 -341 -1531 -323
rect -1565 -391 -1531 -379
rect -1565 -413 -1531 -391
rect -1565 -459 -1531 -451
rect -1565 -485 -1531 -459
rect -1307 459 -1273 485
rect -1307 451 -1273 459
rect -1307 391 -1273 413
rect -1307 379 -1273 391
rect -1307 323 -1273 341
rect -1307 307 -1273 323
rect -1307 255 -1273 269
rect -1307 235 -1273 255
rect -1307 187 -1273 197
rect -1307 163 -1273 187
rect -1307 119 -1273 125
rect -1307 91 -1273 119
rect -1307 51 -1273 53
rect -1307 19 -1273 51
rect -1307 -51 -1273 -19
rect -1307 -53 -1273 -51
rect -1307 -119 -1273 -91
rect -1307 -125 -1273 -119
rect -1307 -187 -1273 -163
rect -1307 -197 -1273 -187
rect -1307 -255 -1273 -235
rect -1307 -269 -1273 -255
rect -1307 -323 -1273 -307
rect -1307 -341 -1273 -323
rect -1307 -391 -1273 -379
rect -1307 -413 -1273 -391
rect -1307 -459 -1273 -451
rect -1307 -485 -1273 -459
rect -1049 459 -1015 485
rect -1049 451 -1015 459
rect -1049 391 -1015 413
rect -1049 379 -1015 391
rect -1049 323 -1015 341
rect -1049 307 -1015 323
rect -1049 255 -1015 269
rect -1049 235 -1015 255
rect -1049 187 -1015 197
rect -1049 163 -1015 187
rect -1049 119 -1015 125
rect -1049 91 -1015 119
rect -1049 51 -1015 53
rect -1049 19 -1015 51
rect -1049 -51 -1015 -19
rect -1049 -53 -1015 -51
rect -1049 -119 -1015 -91
rect -1049 -125 -1015 -119
rect -1049 -187 -1015 -163
rect -1049 -197 -1015 -187
rect -1049 -255 -1015 -235
rect -1049 -269 -1015 -255
rect -1049 -323 -1015 -307
rect -1049 -341 -1015 -323
rect -1049 -391 -1015 -379
rect -1049 -413 -1015 -391
rect -1049 -459 -1015 -451
rect -1049 -485 -1015 -459
rect -791 459 -757 485
rect -791 451 -757 459
rect -791 391 -757 413
rect -791 379 -757 391
rect -791 323 -757 341
rect -791 307 -757 323
rect -791 255 -757 269
rect -791 235 -757 255
rect -791 187 -757 197
rect -791 163 -757 187
rect -791 119 -757 125
rect -791 91 -757 119
rect -791 51 -757 53
rect -791 19 -757 51
rect -791 -51 -757 -19
rect -791 -53 -757 -51
rect -791 -119 -757 -91
rect -791 -125 -757 -119
rect -791 -187 -757 -163
rect -791 -197 -757 -187
rect -791 -255 -757 -235
rect -791 -269 -757 -255
rect -791 -323 -757 -307
rect -791 -341 -757 -323
rect -791 -391 -757 -379
rect -791 -413 -757 -391
rect -791 -459 -757 -451
rect -791 -485 -757 -459
rect -533 459 -499 485
rect -533 451 -499 459
rect -533 391 -499 413
rect -533 379 -499 391
rect -533 323 -499 341
rect -533 307 -499 323
rect -533 255 -499 269
rect -533 235 -499 255
rect -533 187 -499 197
rect -533 163 -499 187
rect -533 119 -499 125
rect -533 91 -499 119
rect -533 51 -499 53
rect -533 19 -499 51
rect -533 -51 -499 -19
rect -533 -53 -499 -51
rect -533 -119 -499 -91
rect -533 -125 -499 -119
rect -533 -187 -499 -163
rect -533 -197 -499 -187
rect -533 -255 -499 -235
rect -533 -269 -499 -255
rect -533 -323 -499 -307
rect -533 -341 -499 -323
rect -533 -391 -499 -379
rect -533 -413 -499 -391
rect -533 -459 -499 -451
rect -533 -485 -499 -459
rect -275 459 -241 485
rect -275 451 -241 459
rect -275 391 -241 413
rect -275 379 -241 391
rect -275 323 -241 341
rect -275 307 -241 323
rect -275 255 -241 269
rect -275 235 -241 255
rect -275 187 -241 197
rect -275 163 -241 187
rect -275 119 -241 125
rect -275 91 -241 119
rect -275 51 -241 53
rect -275 19 -241 51
rect -275 -51 -241 -19
rect -275 -53 -241 -51
rect -275 -119 -241 -91
rect -275 -125 -241 -119
rect -275 -187 -241 -163
rect -275 -197 -241 -187
rect -275 -255 -241 -235
rect -275 -269 -241 -255
rect -275 -323 -241 -307
rect -275 -341 -241 -323
rect -275 -391 -241 -379
rect -275 -413 -241 -391
rect -275 -459 -241 -451
rect -275 -485 -241 -459
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect 241 459 275 485
rect 241 451 275 459
rect 241 391 275 413
rect 241 379 275 391
rect 241 323 275 341
rect 241 307 275 323
rect 241 255 275 269
rect 241 235 275 255
rect 241 187 275 197
rect 241 163 275 187
rect 241 119 275 125
rect 241 91 275 119
rect 241 51 275 53
rect 241 19 275 51
rect 241 -51 275 -19
rect 241 -53 275 -51
rect 241 -119 275 -91
rect 241 -125 275 -119
rect 241 -187 275 -163
rect 241 -197 275 -187
rect 241 -255 275 -235
rect 241 -269 275 -255
rect 241 -323 275 -307
rect 241 -341 275 -323
rect 241 -391 275 -379
rect 241 -413 275 -391
rect 241 -459 275 -451
rect 241 -485 275 -459
rect 499 459 533 485
rect 499 451 533 459
rect 499 391 533 413
rect 499 379 533 391
rect 499 323 533 341
rect 499 307 533 323
rect 499 255 533 269
rect 499 235 533 255
rect 499 187 533 197
rect 499 163 533 187
rect 499 119 533 125
rect 499 91 533 119
rect 499 51 533 53
rect 499 19 533 51
rect 499 -51 533 -19
rect 499 -53 533 -51
rect 499 -119 533 -91
rect 499 -125 533 -119
rect 499 -187 533 -163
rect 499 -197 533 -187
rect 499 -255 533 -235
rect 499 -269 533 -255
rect 499 -323 533 -307
rect 499 -341 533 -323
rect 499 -391 533 -379
rect 499 -413 533 -391
rect 499 -459 533 -451
rect 499 -485 533 -459
rect 757 459 791 485
rect 757 451 791 459
rect 757 391 791 413
rect 757 379 791 391
rect 757 323 791 341
rect 757 307 791 323
rect 757 255 791 269
rect 757 235 791 255
rect 757 187 791 197
rect 757 163 791 187
rect 757 119 791 125
rect 757 91 791 119
rect 757 51 791 53
rect 757 19 791 51
rect 757 -51 791 -19
rect 757 -53 791 -51
rect 757 -119 791 -91
rect 757 -125 791 -119
rect 757 -187 791 -163
rect 757 -197 791 -187
rect 757 -255 791 -235
rect 757 -269 791 -255
rect 757 -323 791 -307
rect 757 -341 791 -323
rect 757 -391 791 -379
rect 757 -413 791 -391
rect 757 -459 791 -451
rect 757 -485 791 -459
rect 1015 459 1049 485
rect 1015 451 1049 459
rect 1015 391 1049 413
rect 1015 379 1049 391
rect 1015 323 1049 341
rect 1015 307 1049 323
rect 1015 255 1049 269
rect 1015 235 1049 255
rect 1015 187 1049 197
rect 1015 163 1049 187
rect 1015 119 1049 125
rect 1015 91 1049 119
rect 1015 51 1049 53
rect 1015 19 1049 51
rect 1015 -51 1049 -19
rect 1015 -53 1049 -51
rect 1015 -119 1049 -91
rect 1015 -125 1049 -119
rect 1015 -187 1049 -163
rect 1015 -197 1049 -187
rect 1015 -255 1049 -235
rect 1015 -269 1049 -255
rect 1015 -323 1049 -307
rect 1015 -341 1049 -323
rect 1015 -391 1049 -379
rect 1015 -413 1049 -391
rect 1015 -459 1049 -451
rect 1015 -485 1049 -459
rect 1273 459 1307 485
rect 1273 451 1307 459
rect 1273 391 1307 413
rect 1273 379 1307 391
rect 1273 323 1307 341
rect 1273 307 1307 323
rect 1273 255 1307 269
rect 1273 235 1307 255
rect 1273 187 1307 197
rect 1273 163 1307 187
rect 1273 119 1307 125
rect 1273 91 1307 119
rect 1273 51 1307 53
rect 1273 19 1307 51
rect 1273 -51 1307 -19
rect 1273 -53 1307 -51
rect 1273 -119 1307 -91
rect 1273 -125 1307 -119
rect 1273 -187 1307 -163
rect 1273 -197 1307 -187
rect 1273 -255 1307 -235
rect 1273 -269 1307 -255
rect 1273 -323 1307 -307
rect 1273 -341 1307 -323
rect 1273 -391 1307 -379
rect 1273 -413 1307 -391
rect 1273 -459 1307 -451
rect 1273 -485 1307 -459
rect 1531 459 1565 485
rect 1531 451 1565 459
rect 1531 391 1565 413
rect 1531 379 1565 391
rect 1531 323 1565 341
rect 1531 307 1565 323
rect 1531 255 1565 269
rect 1531 235 1565 255
rect 1531 187 1565 197
rect 1531 163 1565 187
rect 1531 119 1565 125
rect 1531 91 1565 119
rect 1531 51 1565 53
rect 1531 19 1565 51
rect 1531 -51 1565 -19
rect 1531 -53 1565 -51
rect 1531 -119 1565 -91
rect 1531 -125 1565 -119
rect 1531 -187 1565 -163
rect 1531 -197 1565 -187
rect 1531 -255 1565 -235
rect 1531 -269 1565 -255
rect 1531 -323 1565 -307
rect 1531 -341 1565 -323
rect 1531 -391 1565 -379
rect 1531 -413 1565 -391
rect 1531 -459 1565 -451
rect 1531 -485 1565 -459
rect 1789 459 1823 485
rect 1789 451 1823 459
rect 1789 391 1823 413
rect 1789 379 1823 391
rect 1789 323 1823 341
rect 1789 307 1823 323
rect 1789 255 1823 269
rect 1789 235 1823 255
rect 1789 187 1823 197
rect 1789 163 1823 187
rect 1789 119 1823 125
rect 1789 91 1823 119
rect 1789 51 1823 53
rect 1789 19 1823 51
rect 1789 -51 1823 -19
rect 1789 -53 1823 -51
rect 1789 -119 1823 -91
rect 1789 -125 1823 -119
rect 1789 -187 1823 -163
rect 1789 -197 1823 -187
rect 1789 -255 1823 -235
rect 1789 -269 1823 -255
rect 1789 -323 1823 -307
rect 1789 -341 1823 -323
rect 1789 -391 1823 -379
rect 1789 -413 1823 -391
rect 1789 -459 1823 -451
rect 1789 -485 1823 -459
rect 2047 459 2081 485
rect 2047 451 2081 459
rect 2047 391 2081 413
rect 2047 379 2081 391
rect 2047 323 2081 341
rect 2047 307 2081 323
rect 2047 255 2081 269
rect 2047 235 2081 255
rect 2047 187 2081 197
rect 2047 163 2081 187
rect 2047 119 2081 125
rect 2047 91 2081 119
rect 2047 51 2081 53
rect 2047 19 2081 51
rect 2047 -51 2081 -19
rect 2047 -53 2081 -51
rect 2047 -119 2081 -91
rect 2047 -125 2081 -119
rect 2047 -187 2081 -163
rect 2047 -197 2081 -187
rect 2047 -255 2081 -235
rect 2047 -269 2081 -255
rect 2047 -323 2081 -307
rect 2047 -341 2081 -323
rect 2047 -391 2081 -379
rect 2047 -413 2081 -391
rect 2047 -459 2081 -451
rect 2047 -485 2081 -459
rect 2305 459 2339 485
rect 2305 451 2339 459
rect 2305 391 2339 413
rect 2305 379 2339 391
rect 2305 323 2339 341
rect 2305 307 2339 323
rect 2305 255 2339 269
rect 2305 235 2339 255
rect 2305 187 2339 197
rect 2305 163 2339 187
rect 2305 119 2339 125
rect 2305 91 2339 119
rect 2305 51 2339 53
rect 2305 19 2339 51
rect 2305 -51 2339 -19
rect 2305 -53 2339 -51
rect 2305 -119 2339 -91
rect 2305 -125 2339 -119
rect 2305 -187 2339 -163
rect 2305 -197 2339 -187
rect 2305 -255 2339 -235
rect 2305 -269 2339 -255
rect 2305 -323 2339 -307
rect 2305 -341 2339 -323
rect 2305 -391 2339 -379
rect 2305 -413 2339 -391
rect 2305 -459 2339 -451
rect 2305 -485 2339 -459
rect 2563 459 2597 485
rect 2563 451 2597 459
rect 2563 391 2597 413
rect 2563 379 2597 391
rect 2563 323 2597 341
rect 2563 307 2597 323
rect 2563 255 2597 269
rect 2563 235 2597 255
rect 2563 187 2597 197
rect 2563 163 2597 187
rect 2563 119 2597 125
rect 2563 91 2597 119
rect 2563 51 2597 53
rect 2563 19 2597 51
rect 2563 -51 2597 -19
rect 2563 -53 2597 -51
rect 2563 -119 2597 -91
rect 2563 -125 2597 -119
rect 2563 -187 2597 -163
rect 2563 -197 2597 -187
rect 2563 -255 2597 -235
rect 2563 -269 2597 -255
rect 2563 -323 2597 -307
rect 2563 -341 2597 -323
rect 2563 -391 2597 -379
rect 2563 -413 2597 -391
rect 2563 -459 2597 -451
rect 2563 -485 2597 -459
rect -2425 -1017 -2391 -983
rect -2225 -1017 -2191 -983
rect -2025 -1017 -1991 -983
rect -1825 -1017 -1791 -983
rect -1625 -1017 -1591 -983
rect -1425 -1017 -1391 -983
rect -1225 -1017 -1191 -983
rect -1025 -1017 -991 -983
rect -825 -1017 -791 -983
rect -625 -1017 -591 -983
rect -425 -1017 -391 -983
rect -225 -1017 -191 -983
rect -25 -1017 9 -983
rect 175 -1017 209 -983
rect 375 -1017 409 -983
rect 575 -1017 609 -983
rect 775 -1017 809 -983
rect 975 -1017 1009 -983
rect 1175 -1017 1209 -983
rect 1375 -1017 1409 -983
rect 1575 -1017 1609 -983
rect 1775 -1017 1809 -983
rect 1975 -1017 2009 -983
rect 2175 -1017 2209 -983
rect 2375 -1017 2409 -983
<< metal1 >>
rect -2706 897 2608 940
rect -2706 863 -2425 897
rect -2391 863 -2225 897
rect -2191 863 -2025 897
rect -1991 863 -1825 897
rect -1791 863 -1625 897
rect -1591 863 -1425 897
rect -1391 863 -1225 897
rect -1191 863 -1025 897
rect -991 863 -825 897
rect -791 863 -625 897
rect -591 863 -425 897
rect -391 863 -225 897
rect -191 863 -25 897
rect 9 863 175 897
rect 209 863 375 897
rect 409 863 575 897
rect 609 863 775 897
rect 809 863 975 897
rect 1009 863 1175 897
rect 1209 863 1375 897
rect 1409 863 1575 897
rect 1609 863 1775 897
rect 1809 863 1975 897
rect 2009 863 2175 897
rect 2209 863 2375 897
rect 2409 863 2608 897
rect -2706 820 2608 863
rect -2603 485 -2557 500
rect -2603 451 -2597 485
rect -2563 451 -2557 485
rect -2603 413 -2557 451
rect -2603 379 -2597 413
rect -2563 379 -2557 413
rect -2603 341 -2557 379
rect -2603 307 -2597 341
rect -2563 307 -2557 341
rect -2603 269 -2557 307
rect -2603 235 -2597 269
rect -2563 235 -2557 269
rect -2603 197 -2557 235
rect -2603 163 -2597 197
rect -2563 163 -2557 197
rect -2603 125 -2557 163
rect -2603 91 -2597 125
rect -2563 91 -2557 125
rect -2603 53 -2557 91
rect -2603 19 -2597 53
rect -2563 19 -2557 53
rect -2603 -19 -2557 19
rect -2603 -53 -2597 -19
rect -2563 -53 -2557 -19
rect -2603 -91 -2557 -53
rect -2603 -125 -2597 -91
rect -2563 -125 -2557 -91
rect -2603 -163 -2557 -125
rect -2603 -197 -2597 -163
rect -2563 -197 -2557 -163
rect -2603 -235 -2557 -197
rect -2603 -269 -2597 -235
rect -2563 -269 -2557 -235
rect -2603 -307 -2557 -269
rect -2603 -341 -2597 -307
rect -2563 -341 -2557 -307
rect -2603 -379 -2557 -341
rect -2603 -413 -2597 -379
rect -2563 -413 -2557 -379
rect -2603 -451 -2557 -413
rect -2603 -485 -2597 -451
rect -2563 -485 -2557 -451
rect -2603 -500 -2557 -485
rect -2345 485 -2299 500
rect -2345 451 -2339 485
rect -2305 451 -2299 485
rect -2345 413 -2299 451
rect -2345 379 -2339 413
rect -2305 379 -2299 413
rect -2345 341 -2299 379
rect -2345 307 -2339 341
rect -2305 307 -2299 341
rect -2345 269 -2299 307
rect -2345 235 -2339 269
rect -2305 235 -2299 269
rect -2345 197 -2299 235
rect -2345 163 -2339 197
rect -2305 163 -2299 197
rect -2345 125 -2299 163
rect -2345 91 -2339 125
rect -2305 91 -2299 125
rect -2345 53 -2299 91
rect -2345 19 -2339 53
rect -2305 19 -2299 53
rect -2345 -19 -2299 19
rect -2345 -53 -2339 -19
rect -2305 -53 -2299 -19
rect -2345 -91 -2299 -53
rect -2345 -125 -2339 -91
rect -2305 -125 -2299 -91
rect -2345 -163 -2299 -125
rect -2345 -197 -2339 -163
rect -2305 -197 -2299 -163
rect -2345 -235 -2299 -197
rect -2345 -269 -2339 -235
rect -2305 -269 -2299 -235
rect -2345 -307 -2299 -269
rect -2345 -341 -2339 -307
rect -2305 -341 -2299 -307
rect -2345 -379 -2299 -341
rect -2345 -413 -2339 -379
rect -2305 -413 -2299 -379
rect -2345 -451 -2299 -413
rect -2345 -485 -2339 -451
rect -2305 -485 -2299 -451
rect -2345 -500 -2299 -485
rect -2087 485 -2041 500
rect -2087 451 -2081 485
rect -2047 451 -2041 485
rect -2087 413 -2041 451
rect -2087 379 -2081 413
rect -2047 379 -2041 413
rect -2087 341 -2041 379
rect -2087 307 -2081 341
rect -2047 307 -2041 341
rect -2087 269 -2041 307
rect -2087 235 -2081 269
rect -2047 235 -2041 269
rect -2087 197 -2041 235
rect -2087 163 -2081 197
rect -2047 163 -2041 197
rect -2087 125 -2041 163
rect -2087 91 -2081 125
rect -2047 91 -2041 125
rect -2087 53 -2041 91
rect -2087 19 -2081 53
rect -2047 19 -2041 53
rect -2087 -19 -2041 19
rect -2087 -53 -2081 -19
rect -2047 -53 -2041 -19
rect -2087 -91 -2041 -53
rect -2087 -125 -2081 -91
rect -2047 -125 -2041 -91
rect -2087 -163 -2041 -125
rect -2087 -197 -2081 -163
rect -2047 -197 -2041 -163
rect -2087 -235 -2041 -197
rect -2087 -269 -2081 -235
rect -2047 -269 -2041 -235
rect -2087 -307 -2041 -269
rect -2087 -341 -2081 -307
rect -2047 -341 -2041 -307
rect -2087 -379 -2041 -341
rect -2087 -413 -2081 -379
rect -2047 -413 -2041 -379
rect -2087 -451 -2041 -413
rect -2087 -485 -2081 -451
rect -2047 -485 -2041 -451
rect -2087 -500 -2041 -485
rect -1829 485 -1783 500
rect -1829 451 -1823 485
rect -1789 451 -1783 485
rect -1829 413 -1783 451
rect -1829 379 -1823 413
rect -1789 379 -1783 413
rect -1829 341 -1783 379
rect -1829 307 -1823 341
rect -1789 307 -1783 341
rect -1829 269 -1783 307
rect -1829 235 -1823 269
rect -1789 235 -1783 269
rect -1829 197 -1783 235
rect -1829 163 -1823 197
rect -1789 163 -1783 197
rect -1829 125 -1783 163
rect -1829 91 -1823 125
rect -1789 91 -1783 125
rect -1829 53 -1783 91
rect -1829 19 -1823 53
rect -1789 19 -1783 53
rect -1829 -19 -1783 19
rect -1829 -53 -1823 -19
rect -1789 -53 -1783 -19
rect -1829 -91 -1783 -53
rect -1829 -125 -1823 -91
rect -1789 -125 -1783 -91
rect -1829 -163 -1783 -125
rect -1829 -197 -1823 -163
rect -1789 -197 -1783 -163
rect -1829 -235 -1783 -197
rect -1829 -269 -1823 -235
rect -1789 -269 -1783 -235
rect -1829 -307 -1783 -269
rect -1829 -341 -1823 -307
rect -1789 -341 -1783 -307
rect -1829 -379 -1783 -341
rect -1829 -413 -1823 -379
rect -1789 -413 -1783 -379
rect -1829 -451 -1783 -413
rect -1829 -485 -1823 -451
rect -1789 -485 -1783 -451
rect -1829 -500 -1783 -485
rect -1571 485 -1525 500
rect -1571 451 -1565 485
rect -1531 451 -1525 485
rect -1571 413 -1525 451
rect -1571 379 -1565 413
rect -1531 379 -1525 413
rect -1571 341 -1525 379
rect -1571 307 -1565 341
rect -1531 307 -1525 341
rect -1571 269 -1525 307
rect -1571 235 -1565 269
rect -1531 235 -1525 269
rect -1571 197 -1525 235
rect -1571 163 -1565 197
rect -1531 163 -1525 197
rect -1571 125 -1525 163
rect -1571 91 -1565 125
rect -1531 91 -1525 125
rect -1571 53 -1525 91
rect -1571 19 -1565 53
rect -1531 19 -1525 53
rect -1571 -19 -1525 19
rect -1571 -53 -1565 -19
rect -1531 -53 -1525 -19
rect -1571 -91 -1525 -53
rect -1571 -125 -1565 -91
rect -1531 -125 -1525 -91
rect -1571 -163 -1525 -125
rect -1571 -197 -1565 -163
rect -1531 -197 -1525 -163
rect -1571 -235 -1525 -197
rect -1571 -269 -1565 -235
rect -1531 -269 -1525 -235
rect -1571 -307 -1525 -269
rect -1571 -341 -1565 -307
rect -1531 -341 -1525 -307
rect -1571 -379 -1525 -341
rect -1571 -413 -1565 -379
rect -1531 -413 -1525 -379
rect -1571 -451 -1525 -413
rect -1571 -485 -1565 -451
rect -1531 -485 -1525 -451
rect -1571 -500 -1525 -485
rect -1313 485 -1267 500
rect -1313 451 -1307 485
rect -1273 451 -1267 485
rect -1313 413 -1267 451
rect -1313 379 -1307 413
rect -1273 379 -1267 413
rect -1313 341 -1267 379
rect -1313 307 -1307 341
rect -1273 307 -1267 341
rect -1313 269 -1267 307
rect -1313 235 -1307 269
rect -1273 235 -1267 269
rect -1313 197 -1267 235
rect -1313 163 -1307 197
rect -1273 163 -1267 197
rect -1313 125 -1267 163
rect -1313 91 -1307 125
rect -1273 91 -1267 125
rect -1313 53 -1267 91
rect -1313 19 -1307 53
rect -1273 19 -1267 53
rect -1313 -19 -1267 19
rect -1313 -53 -1307 -19
rect -1273 -53 -1267 -19
rect -1313 -91 -1267 -53
rect -1313 -125 -1307 -91
rect -1273 -125 -1267 -91
rect -1313 -163 -1267 -125
rect -1313 -197 -1307 -163
rect -1273 -197 -1267 -163
rect -1313 -235 -1267 -197
rect -1313 -269 -1307 -235
rect -1273 -269 -1267 -235
rect -1313 -307 -1267 -269
rect -1313 -341 -1307 -307
rect -1273 -341 -1267 -307
rect -1313 -379 -1267 -341
rect -1313 -413 -1307 -379
rect -1273 -413 -1267 -379
rect -1313 -451 -1267 -413
rect -1313 -485 -1307 -451
rect -1273 -485 -1267 -451
rect -1313 -500 -1267 -485
rect -1055 485 -1009 500
rect -1055 451 -1049 485
rect -1015 451 -1009 485
rect -1055 413 -1009 451
rect -1055 379 -1049 413
rect -1015 379 -1009 413
rect -1055 341 -1009 379
rect -1055 307 -1049 341
rect -1015 307 -1009 341
rect -1055 269 -1009 307
rect -1055 235 -1049 269
rect -1015 235 -1009 269
rect -1055 197 -1009 235
rect -1055 163 -1049 197
rect -1015 163 -1009 197
rect -1055 125 -1009 163
rect -1055 91 -1049 125
rect -1015 91 -1009 125
rect -1055 53 -1009 91
rect -1055 19 -1049 53
rect -1015 19 -1009 53
rect -1055 -19 -1009 19
rect -1055 -53 -1049 -19
rect -1015 -53 -1009 -19
rect -1055 -91 -1009 -53
rect -1055 -125 -1049 -91
rect -1015 -125 -1009 -91
rect -1055 -163 -1009 -125
rect -1055 -197 -1049 -163
rect -1015 -197 -1009 -163
rect -1055 -235 -1009 -197
rect -1055 -269 -1049 -235
rect -1015 -269 -1009 -235
rect -1055 -307 -1009 -269
rect -1055 -341 -1049 -307
rect -1015 -341 -1009 -307
rect -1055 -379 -1009 -341
rect -1055 -413 -1049 -379
rect -1015 -413 -1009 -379
rect -1055 -451 -1009 -413
rect -1055 -485 -1049 -451
rect -1015 -485 -1009 -451
rect -1055 -500 -1009 -485
rect -797 485 -751 500
rect -797 451 -791 485
rect -757 451 -751 485
rect -797 413 -751 451
rect -797 379 -791 413
rect -757 379 -751 413
rect -797 341 -751 379
rect -797 307 -791 341
rect -757 307 -751 341
rect -797 269 -751 307
rect -797 235 -791 269
rect -757 235 -751 269
rect -797 197 -751 235
rect -797 163 -791 197
rect -757 163 -751 197
rect -797 125 -751 163
rect -797 91 -791 125
rect -757 91 -751 125
rect -797 53 -751 91
rect -797 19 -791 53
rect -757 19 -751 53
rect -797 -19 -751 19
rect -797 -53 -791 -19
rect -757 -53 -751 -19
rect -797 -91 -751 -53
rect -797 -125 -791 -91
rect -757 -125 -751 -91
rect -797 -163 -751 -125
rect -797 -197 -791 -163
rect -757 -197 -751 -163
rect -797 -235 -751 -197
rect -797 -269 -791 -235
rect -757 -269 -751 -235
rect -797 -307 -751 -269
rect -797 -341 -791 -307
rect -757 -341 -751 -307
rect -797 -379 -751 -341
rect -797 -413 -791 -379
rect -757 -413 -751 -379
rect -797 -451 -751 -413
rect -797 -485 -791 -451
rect -757 -485 -751 -451
rect -797 -500 -751 -485
rect -539 485 -493 500
rect -539 451 -533 485
rect -499 451 -493 485
rect -539 413 -493 451
rect -539 379 -533 413
rect -499 379 -493 413
rect -539 341 -493 379
rect -539 307 -533 341
rect -499 307 -493 341
rect -539 269 -493 307
rect -539 235 -533 269
rect -499 235 -493 269
rect -539 197 -493 235
rect -539 163 -533 197
rect -499 163 -493 197
rect -539 125 -493 163
rect -539 91 -533 125
rect -499 91 -493 125
rect -539 53 -493 91
rect -539 19 -533 53
rect -499 19 -493 53
rect -539 -19 -493 19
rect -539 -53 -533 -19
rect -499 -53 -493 -19
rect -539 -91 -493 -53
rect -539 -125 -533 -91
rect -499 -125 -493 -91
rect -539 -163 -493 -125
rect -539 -197 -533 -163
rect -499 -197 -493 -163
rect -539 -235 -493 -197
rect -539 -269 -533 -235
rect -499 -269 -493 -235
rect -539 -307 -493 -269
rect -539 -341 -533 -307
rect -499 -341 -493 -307
rect -539 -379 -493 -341
rect -539 -413 -533 -379
rect -499 -413 -493 -379
rect -539 -451 -493 -413
rect -539 -485 -533 -451
rect -499 -485 -493 -451
rect -539 -500 -493 -485
rect -281 485 -235 500
rect -281 451 -275 485
rect -241 451 -235 485
rect -281 413 -235 451
rect -281 379 -275 413
rect -241 379 -235 413
rect -281 341 -235 379
rect -281 307 -275 341
rect -241 307 -235 341
rect -281 269 -235 307
rect -281 235 -275 269
rect -241 235 -235 269
rect -281 197 -235 235
rect -281 163 -275 197
rect -241 163 -235 197
rect -281 125 -235 163
rect -281 91 -275 125
rect -241 91 -235 125
rect -281 53 -235 91
rect -281 19 -275 53
rect -241 19 -235 53
rect -281 -19 -235 19
rect -281 -53 -275 -19
rect -241 -53 -235 -19
rect -281 -91 -235 -53
rect -281 -125 -275 -91
rect -241 -125 -235 -91
rect -281 -163 -235 -125
rect -281 -197 -275 -163
rect -241 -197 -235 -163
rect -281 -235 -235 -197
rect -281 -269 -275 -235
rect -241 -269 -235 -235
rect -281 -307 -235 -269
rect -281 -341 -275 -307
rect -241 -341 -235 -307
rect -281 -379 -235 -341
rect -281 -413 -275 -379
rect -241 -413 -235 -379
rect -281 -451 -235 -413
rect -281 -485 -275 -451
rect -241 -485 -235 -451
rect -281 -500 -235 -485
rect -23 485 23 500
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -500 23 -485
rect 235 485 281 500
rect 235 451 241 485
rect 275 451 281 485
rect 235 413 281 451
rect 235 379 241 413
rect 275 379 281 413
rect 235 341 281 379
rect 235 307 241 341
rect 275 307 281 341
rect 235 269 281 307
rect 235 235 241 269
rect 275 235 281 269
rect 235 197 281 235
rect 235 163 241 197
rect 275 163 281 197
rect 235 125 281 163
rect 235 91 241 125
rect 275 91 281 125
rect 235 53 281 91
rect 235 19 241 53
rect 275 19 281 53
rect 235 -19 281 19
rect 235 -53 241 -19
rect 275 -53 281 -19
rect 235 -91 281 -53
rect 235 -125 241 -91
rect 275 -125 281 -91
rect 235 -163 281 -125
rect 235 -197 241 -163
rect 275 -197 281 -163
rect 235 -235 281 -197
rect 235 -269 241 -235
rect 275 -269 281 -235
rect 235 -307 281 -269
rect 235 -341 241 -307
rect 275 -341 281 -307
rect 235 -379 281 -341
rect 235 -413 241 -379
rect 275 -413 281 -379
rect 235 -451 281 -413
rect 235 -485 241 -451
rect 275 -485 281 -451
rect 235 -500 281 -485
rect 493 485 539 500
rect 493 451 499 485
rect 533 451 539 485
rect 493 413 539 451
rect 493 379 499 413
rect 533 379 539 413
rect 493 341 539 379
rect 493 307 499 341
rect 533 307 539 341
rect 493 269 539 307
rect 493 235 499 269
rect 533 235 539 269
rect 493 197 539 235
rect 493 163 499 197
rect 533 163 539 197
rect 493 125 539 163
rect 493 91 499 125
rect 533 91 539 125
rect 493 53 539 91
rect 493 19 499 53
rect 533 19 539 53
rect 493 -19 539 19
rect 493 -53 499 -19
rect 533 -53 539 -19
rect 493 -91 539 -53
rect 493 -125 499 -91
rect 533 -125 539 -91
rect 493 -163 539 -125
rect 493 -197 499 -163
rect 533 -197 539 -163
rect 493 -235 539 -197
rect 493 -269 499 -235
rect 533 -269 539 -235
rect 493 -307 539 -269
rect 493 -341 499 -307
rect 533 -341 539 -307
rect 493 -379 539 -341
rect 493 -413 499 -379
rect 533 -413 539 -379
rect 493 -451 539 -413
rect 493 -485 499 -451
rect 533 -485 539 -451
rect 493 -500 539 -485
rect 751 485 797 500
rect 751 451 757 485
rect 791 451 797 485
rect 751 413 797 451
rect 751 379 757 413
rect 791 379 797 413
rect 751 341 797 379
rect 751 307 757 341
rect 791 307 797 341
rect 751 269 797 307
rect 751 235 757 269
rect 791 235 797 269
rect 751 197 797 235
rect 751 163 757 197
rect 791 163 797 197
rect 751 125 797 163
rect 751 91 757 125
rect 791 91 797 125
rect 751 53 797 91
rect 751 19 757 53
rect 791 19 797 53
rect 751 -19 797 19
rect 751 -53 757 -19
rect 791 -53 797 -19
rect 751 -91 797 -53
rect 751 -125 757 -91
rect 791 -125 797 -91
rect 751 -163 797 -125
rect 751 -197 757 -163
rect 791 -197 797 -163
rect 751 -235 797 -197
rect 751 -269 757 -235
rect 791 -269 797 -235
rect 751 -307 797 -269
rect 751 -341 757 -307
rect 791 -341 797 -307
rect 751 -379 797 -341
rect 751 -413 757 -379
rect 791 -413 797 -379
rect 751 -451 797 -413
rect 751 -485 757 -451
rect 791 -485 797 -451
rect 751 -500 797 -485
rect 1009 485 1055 500
rect 1009 451 1015 485
rect 1049 451 1055 485
rect 1009 413 1055 451
rect 1009 379 1015 413
rect 1049 379 1055 413
rect 1009 341 1055 379
rect 1009 307 1015 341
rect 1049 307 1055 341
rect 1009 269 1055 307
rect 1009 235 1015 269
rect 1049 235 1055 269
rect 1009 197 1055 235
rect 1009 163 1015 197
rect 1049 163 1055 197
rect 1009 125 1055 163
rect 1009 91 1015 125
rect 1049 91 1055 125
rect 1009 53 1055 91
rect 1009 19 1015 53
rect 1049 19 1055 53
rect 1009 -19 1055 19
rect 1009 -53 1015 -19
rect 1049 -53 1055 -19
rect 1009 -91 1055 -53
rect 1009 -125 1015 -91
rect 1049 -125 1055 -91
rect 1009 -163 1055 -125
rect 1009 -197 1015 -163
rect 1049 -197 1055 -163
rect 1009 -235 1055 -197
rect 1009 -269 1015 -235
rect 1049 -269 1055 -235
rect 1009 -307 1055 -269
rect 1009 -341 1015 -307
rect 1049 -341 1055 -307
rect 1009 -379 1055 -341
rect 1009 -413 1015 -379
rect 1049 -413 1055 -379
rect 1009 -451 1055 -413
rect 1009 -485 1015 -451
rect 1049 -485 1055 -451
rect 1009 -500 1055 -485
rect 1267 485 1313 500
rect 1267 451 1273 485
rect 1307 451 1313 485
rect 1267 413 1313 451
rect 1267 379 1273 413
rect 1307 379 1313 413
rect 1267 341 1313 379
rect 1267 307 1273 341
rect 1307 307 1313 341
rect 1267 269 1313 307
rect 1267 235 1273 269
rect 1307 235 1313 269
rect 1267 197 1313 235
rect 1267 163 1273 197
rect 1307 163 1313 197
rect 1267 125 1313 163
rect 1267 91 1273 125
rect 1307 91 1313 125
rect 1267 53 1313 91
rect 1267 19 1273 53
rect 1307 19 1313 53
rect 1267 -19 1313 19
rect 1267 -53 1273 -19
rect 1307 -53 1313 -19
rect 1267 -91 1313 -53
rect 1267 -125 1273 -91
rect 1307 -125 1313 -91
rect 1267 -163 1313 -125
rect 1267 -197 1273 -163
rect 1307 -197 1313 -163
rect 1267 -235 1313 -197
rect 1267 -269 1273 -235
rect 1307 -269 1313 -235
rect 1267 -307 1313 -269
rect 1267 -341 1273 -307
rect 1307 -341 1313 -307
rect 1267 -379 1313 -341
rect 1267 -413 1273 -379
rect 1307 -413 1313 -379
rect 1267 -451 1313 -413
rect 1267 -485 1273 -451
rect 1307 -485 1313 -451
rect 1267 -500 1313 -485
rect 1525 485 1571 500
rect 1525 451 1531 485
rect 1565 451 1571 485
rect 1525 413 1571 451
rect 1525 379 1531 413
rect 1565 379 1571 413
rect 1525 341 1571 379
rect 1525 307 1531 341
rect 1565 307 1571 341
rect 1525 269 1571 307
rect 1525 235 1531 269
rect 1565 235 1571 269
rect 1525 197 1571 235
rect 1525 163 1531 197
rect 1565 163 1571 197
rect 1525 125 1571 163
rect 1525 91 1531 125
rect 1565 91 1571 125
rect 1525 53 1571 91
rect 1525 19 1531 53
rect 1565 19 1571 53
rect 1525 -19 1571 19
rect 1525 -53 1531 -19
rect 1565 -53 1571 -19
rect 1525 -91 1571 -53
rect 1525 -125 1531 -91
rect 1565 -125 1571 -91
rect 1525 -163 1571 -125
rect 1525 -197 1531 -163
rect 1565 -197 1571 -163
rect 1525 -235 1571 -197
rect 1525 -269 1531 -235
rect 1565 -269 1571 -235
rect 1525 -307 1571 -269
rect 1525 -341 1531 -307
rect 1565 -341 1571 -307
rect 1525 -379 1571 -341
rect 1525 -413 1531 -379
rect 1565 -413 1571 -379
rect 1525 -451 1571 -413
rect 1525 -485 1531 -451
rect 1565 -485 1571 -451
rect 1525 -500 1571 -485
rect 1783 485 1829 500
rect 1783 451 1789 485
rect 1823 451 1829 485
rect 1783 413 1829 451
rect 1783 379 1789 413
rect 1823 379 1829 413
rect 1783 341 1829 379
rect 1783 307 1789 341
rect 1823 307 1829 341
rect 1783 269 1829 307
rect 1783 235 1789 269
rect 1823 235 1829 269
rect 1783 197 1829 235
rect 1783 163 1789 197
rect 1823 163 1829 197
rect 1783 125 1829 163
rect 1783 91 1789 125
rect 1823 91 1829 125
rect 1783 53 1829 91
rect 1783 19 1789 53
rect 1823 19 1829 53
rect 1783 -19 1829 19
rect 1783 -53 1789 -19
rect 1823 -53 1829 -19
rect 1783 -91 1829 -53
rect 1783 -125 1789 -91
rect 1823 -125 1829 -91
rect 1783 -163 1829 -125
rect 1783 -197 1789 -163
rect 1823 -197 1829 -163
rect 1783 -235 1829 -197
rect 1783 -269 1789 -235
rect 1823 -269 1829 -235
rect 1783 -307 1829 -269
rect 1783 -341 1789 -307
rect 1823 -341 1829 -307
rect 1783 -379 1829 -341
rect 1783 -413 1789 -379
rect 1823 -413 1829 -379
rect 1783 -451 1829 -413
rect 1783 -485 1789 -451
rect 1823 -485 1829 -451
rect 1783 -500 1829 -485
rect 2041 485 2087 500
rect 2041 451 2047 485
rect 2081 451 2087 485
rect 2041 413 2087 451
rect 2041 379 2047 413
rect 2081 379 2087 413
rect 2041 341 2087 379
rect 2041 307 2047 341
rect 2081 307 2087 341
rect 2041 269 2087 307
rect 2041 235 2047 269
rect 2081 235 2087 269
rect 2041 197 2087 235
rect 2041 163 2047 197
rect 2081 163 2087 197
rect 2041 125 2087 163
rect 2041 91 2047 125
rect 2081 91 2087 125
rect 2041 53 2087 91
rect 2041 19 2047 53
rect 2081 19 2087 53
rect 2041 -19 2087 19
rect 2041 -53 2047 -19
rect 2081 -53 2087 -19
rect 2041 -91 2087 -53
rect 2041 -125 2047 -91
rect 2081 -125 2087 -91
rect 2041 -163 2087 -125
rect 2041 -197 2047 -163
rect 2081 -197 2087 -163
rect 2041 -235 2087 -197
rect 2041 -269 2047 -235
rect 2081 -269 2087 -235
rect 2041 -307 2087 -269
rect 2041 -341 2047 -307
rect 2081 -341 2087 -307
rect 2041 -379 2087 -341
rect 2041 -413 2047 -379
rect 2081 -413 2087 -379
rect 2041 -451 2087 -413
rect 2041 -485 2047 -451
rect 2081 -485 2087 -451
rect 2041 -500 2087 -485
rect 2299 485 2345 500
rect 2299 451 2305 485
rect 2339 451 2345 485
rect 2299 413 2345 451
rect 2299 379 2305 413
rect 2339 379 2345 413
rect 2299 341 2345 379
rect 2299 307 2305 341
rect 2339 307 2345 341
rect 2299 269 2345 307
rect 2299 235 2305 269
rect 2339 235 2345 269
rect 2299 197 2345 235
rect 2299 163 2305 197
rect 2339 163 2345 197
rect 2299 125 2345 163
rect 2299 91 2305 125
rect 2339 91 2345 125
rect 2299 53 2345 91
rect 2299 19 2305 53
rect 2339 19 2345 53
rect 2299 -19 2345 19
rect 2299 -53 2305 -19
rect 2339 -53 2345 -19
rect 2299 -91 2345 -53
rect 2299 -125 2305 -91
rect 2339 -125 2345 -91
rect 2299 -163 2345 -125
rect 2299 -197 2305 -163
rect 2339 -197 2345 -163
rect 2299 -235 2345 -197
rect 2299 -269 2305 -235
rect 2339 -269 2345 -235
rect 2299 -307 2345 -269
rect 2299 -341 2305 -307
rect 2339 -341 2345 -307
rect 2299 -379 2345 -341
rect 2299 -413 2305 -379
rect 2339 -413 2345 -379
rect 2299 -451 2345 -413
rect 2299 -485 2305 -451
rect 2339 -485 2345 -451
rect 2299 -500 2345 -485
rect 2557 485 2603 500
rect 2557 451 2563 485
rect 2597 451 2603 485
rect 2557 413 2603 451
rect 2557 379 2563 413
rect 2597 379 2603 413
rect 2557 341 2603 379
rect 2557 307 2563 341
rect 2597 307 2603 341
rect 2557 269 2603 307
rect 2557 235 2563 269
rect 2597 235 2603 269
rect 2557 197 2603 235
rect 2557 163 2563 197
rect 2597 163 2603 197
rect 2557 125 2603 163
rect 2557 91 2563 125
rect 2597 91 2603 125
rect 2557 53 2603 91
rect 2557 19 2563 53
rect 2597 19 2603 53
rect 2557 -19 2603 19
rect 2557 -53 2563 -19
rect 2597 -53 2603 -19
rect 2557 -91 2603 -53
rect 2557 -125 2563 -91
rect 2597 -125 2603 -91
rect 2557 -163 2603 -125
rect 2557 -197 2563 -163
rect 2597 -197 2603 -163
rect 2557 -235 2603 -197
rect 2557 -269 2563 -235
rect 2597 -269 2603 -235
rect 2557 -307 2603 -269
rect 2557 -341 2563 -307
rect 2597 -341 2603 -307
rect 2557 -379 2603 -341
rect 2557 -413 2563 -379
rect 2597 -413 2603 -379
rect 2557 -451 2603 -413
rect 2557 -485 2563 -451
rect 2597 -485 2603 -451
rect 2557 -500 2603 -485
rect -2706 -983 2608 -940
rect -2706 -1017 -2425 -983
rect -2391 -1017 -2225 -983
rect -2191 -1017 -2025 -983
rect -1991 -1017 -1825 -983
rect -1791 -1017 -1625 -983
rect -1591 -1017 -1425 -983
rect -1391 -1017 -1225 -983
rect -1191 -1017 -1025 -983
rect -991 -1017 -825 -983
rect -791 -1017 -625 -983
rect -591 -1017 -425 -983
rect -391 -1017 -225 -983
rect -191 -1017 -25 -983
rect 9 -1017 175 -983
rect 209 -1017 375 -983
rect 409 -1017 575 -983
rect 609 -1017 775 -983
rect 809 -1017 975 -983
rect 1009 -1017 1175 -983
rect 1209 -1017 1375 -983
rect 1409 -1017 1575 -983
rect 1609 -1017 1775 -983
rect 1809 -1017 1975 -983
rect 2009 -1017 2175 -983
rect 2209 -1017 2375 -983
rect 2409 -1017 2608 -983
rect -2706 -1060 2608 -1017
<< labels >>
flabel metal1 s -2608 850 -2548 910 1 FreeSans 1000 0 0 0 VPWR
port 1 nsew
flabel metal1 s -2608 -1030 -2548 -970 1 FreeSans 1000 0 0 0 VGND
port 2 nsew
flabel locali s 2548 690 2608 750 1 FreeSans 1000 0 0 0 SOURCE
port 3 nsew
flabel locali s 2548 -630 2608 -570 1 FreeSans 1000 0 0 0 DRAIN
port 4 nsew
flabel locali s 2548 -796 2608 -736 1 FreeSans 1000 0 0 0 GATE
port 5 nsew
<< end >>
