magic
tech sky130A
timestamp 1655322987
<< metal3 >>
rect -90 76 90 90
rect -90 -76 -76 76
rect 76 -76 90 76
rect -90 -90 90 -76
<< via3 >>
rect -76 -76 76 76
<< metal4 >>
rect -90 76 90 90
rect -90 -76 -76 76
rect 76 -76 90 76
rect -90 -90 90 -76
<< end >>
