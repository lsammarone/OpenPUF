magic
tech sky130A
timestamp 1656715967
<< metal3 >>
rect -519 76 519 90
rect -519 -76 -516 76
rect 516 -76 519 76
rect -519 -90 519 -76
<< via3 >>
rect -516 -76 516 76
<< metal4 >>
rect -519 76 519 90
rect -519 -76 -516 76
rect 516 -76 519 76
rect -519 -90 519 -76
<< properties >>
string GDS_END 9357394
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/design_merged.gds
string GDS_START 9350606
<< end >>
