magic
tech sky130A
timestamp 1656729169
<< metal1 >>
rect -331 13 331 16
rect -331 -13 -317 13
rect -291 -13 -285 13
rect -259 -13 -253 13
rect -227 -13 -221 13
rect -195 -13 -189 13
rect -163 -13 -157 13
rect -131 -13 -125 13
rect -99 -13 -93 13
rect -67 -13 -61 13
rect -35 -13 -29 13
rect -3 -13 3 13
rect 29 -13 35 13
rect 61 -13 67 13
rect 93 -13 99 13
rect 125 -13 131 13
rect 157 -13 163 13
rect 189 -13 195 13
rect 221 -13 227 13
rect 253 -13 259 13
rect 285 -13 291 13
rect 317 -13 331 13
rect -331 -16 331 -13
<< via1 >>
rect -317 -13 -291 13
rect -285 -13 -259 13
rect -253 -13 -227 13
rect -221 -13 -195 13
rect -189 -13 -163 13
rect -157 -13 -131 13
rect -125 -13 -99 13
rect -93 -13 -67 13
rect -61 -13 -35 13
rect -29 -13 -3 13
rect 3 -13 29 13
rect 35 -13 61 13
rect 67 -13 93 13
rect 99 -13 125 13
rect 131 -13 157 13
rect 163 -13 189 13
rect 195 -13 221 13
rect 227 -13 253 13
rect 259 -13 285 13
rect 291 -13 317 13
<< metal2 >>
rect -331 13 331 16
rect -331 -13 -317 13
rect -291 -13 -285 13
rect -259 -13 -253 13
rect -227 -13 -221 13
rect -195 -13 -189 13
rect -163 -13 -157 13
rect -131 -13 -125 13
rect -99 -13 -93 13
rect -67 -13 -61 13
rect -35 -13 -29 13
rect -3 -13 3 13
rect 29 -13 35 13
rect 61 -13 67 13
rect 93 -13 99 13
rect 125 -13 131 13
rect 157 -13 163 13
rect 189 -13 195 13
rect 221 -13 227 13
rect 253 -13 259 13
rect 285 -13 291 13
rect 317 -13 331 13
rect -331 -16 331 -13
<< properties >>
string GDS_END 9361262
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/merge/design_merged.gds
string GDS_START 9359850
<< end >>
