magic
tech sky130A
magscale 1 2
timestamp 1655322987
<< metal3 >>
rect -1139 152 1138 180
rect -1139 -152 -1112 152
rect 1112 -152 1138 152
rect -1139 -180 1138 -152
<< via3 >>
rect -1112 -152 1112 152
<< metal4 >>
rect -1139 152 1138 180
rect -1139 -152 -1112 152
rect 1112 -152 1138 152
rect -1139 -180 1138 -152
<< end >>
