magic
tech sky130A
magscale 1 2
timestamp 1483428465
<< checkpaint >>
rect -1429 -1440 1429 1440
<< metal3 >>
rect -169 152 169 180
rect -169 -152 -152 152
rect 152 -152 169 152
rect -169 -180 169 -152
<< via3 >>
rect -152 -152 152 152
<< metal4 >>
rect -169 152 169 180
rect -169 -152 -152 152
rect 152 -152 169 152
rect -169 -180 169 -152
<< end >>
