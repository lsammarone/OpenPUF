magic
tech sky130A
magscale 1 2
timestamp 1654825959
<< nwell >>
rect 575170 493276 580556 493654
rect 575169 492152 580556 493276
rect 574448 404400 579834 404778
rect 574447 403276 579834 404400
rect 496808 399925 498454 400022
rect 493048 390125 494694 390222
rect 493048 362516 494695 390125
rect 496808 372316 498455 399925
rect 500568 392281 502214 392378
rect 500568 386656 502215 392281
rect 500801 386655 502215 386656
rect 500568 385617 502214 385714
rect 500568 379992 502215 385617
rect 523128 390125 524774 390222
rect 500801 379991 502215 379992
rect 504328 377483 505974 377580
rect 511848 377483 513494 377580
rect 504328 374606 505975 377483
rect 511848 374606 513495 377483
rect 504561 374605 505975 374606
rect 512081 374605 513495 374606
rect 497041 372315 498455 372316
rect 493281 362515 494695 362516
rect 523128 362516 524775 390125
rect 523361 362515 524775 362516
rect 574644 358972 580030 359350
rect 574643 357848 580030 358972
rect 575092 312804 580478 313182
rect 575091 311680 580478 312804
<< pwell >>
rect 560650 491970 565964 493466
rect 565000 491940 565964 491970
rect 504658 402809 505998 402962
rect 504658 401775 504811 402809
rect 505845 401775 505998 402809
rect 560592 402828 565906 404324
rect 560592 402798 561556 402828
rect 504658 401622 505998 401775
rect 497322 400294 498174 400862
rect 498522 400830 498694 400922
rect 493992 392568 494224 393236
rect 493562 390494 494414 391062
rect 494762 391030 494934 391122
rect 505272 399722 505504 400390
rect 505272 396978 505504 397646
rect 512792 396880 513024 397548
rect 505272 393946 505504 394614
rect 509032 394136 509264 394804
rect 512792 394136 513024 394804
rect 505272 390902 505504 391570
rect 509032 391104 509264 391772
rect 512792 391392 513024 392060
rect 516552 391000 516784 391668
rect 504842 385330 505694 389562
rect 506042 389530 506214 389622
rect 506112 388390 506214 388562
rect 506112 387090 506214 387262
rect 512792 386198 513024 386866
rect 516122 385330 516974 389562
rect 517322 389530 517494 389622
rect 520312 389530 520544 390198
rect 517392 388390 517494 388562
rect 517392 387090 517494 387262
rect 520312 386198 520544 386866
rect 520312 383454 520544 384122
rect 520312 380220 520544 380888
rect 501082 373472 501934 377704
rect 502282 377672 502454 377764
rect 502352 376532 502454 376704
rect 502352 375232 502454 375404
rect 516552 376006 516784 376674
rect 520312 376006 520544 376674
rect 516552 373262 516784 373930
rect 520312 373262 520544 373930
rect 500898 373017 502238 373170
rect 497138 371841 498478 371994
rect 497138 370807 497291 371841
rect 498325 370807 498478 371841
rect 497138 370501 498478 370807
rect 497138 369467 497291 370501
rect 498325 369467 498478 370501
rect 497138 369161 498478 369467
rect 497138 368127 497291 369161
rect 498325 368127 498478 369161
rect 497138 367821 498478 368127
rect 497138 366787 497291 367821
rect 498325 366787 498478 367821
rect 497138 366481 498478 366787
rect 497138 365447 497291 366481
rect 498325 365447 498478 366481
rect 497138 365141 498478 365447
rect 497138 364107 497291 365141
rect 498325 364107 498478 365141
rect 497138 363801 498478 364107
rect 497138 362767 497291 363801
rect 498325 362767 498478 363801
rect 497138 362614 498478 362767
rect 500898 371983 501051 373017
rect 502085 371983 502238 373017
rect 500898 371677 502238 371983
rect 500898 370643 501051 371677
rect 502085 370643 502238 371677
rect 500898 370337 502238 370643
rect 500898 369303 501051 370337
rect 502085 369303 502238 370337
rect 500898 368997 502238 369303
rect 500898 367963 501051 368997
rect 502085 367963 502238 368997
rect 500898 367657 502238 367963
rect 500898 366623 501051 367657
rect 502085 366623 502238 367657
rect 500898 366317 502238 366623
rect 500898 365283 501051 366317
rect 502085 365283 502238 366317
rect 500898 364977 502238 365283
rect 500898 363943 501051 364977
rect 502085 363943 502238 364977
rect 500898 363637 502238 363943
rect 500898 362603 501051 363637
rect 502085 362603 502238 363637
rect 500898 362450 502238 362603
rect 504658 373017 505998 373170
rect 504658 371983 504811 373017
rect 505845 371983 505998 373017
rect 504658 371677 505998 371983
rect 504658 370643 504811 371677
rect 505845 370643 505998 371677
rect 504658 370337 505998 370643
rect 504658 369303 504811 370337
rect 505845 369303 505998 370337
rect 504658 368997 505998 369303
rect 504658 367963 504811 368997
rect 505845 367963 505998 368997
rect 504658 367657 505998 367963
rect 504658 366623 504811 367657
rect 505845 366623 505998 367657
rect 504658 366317 505998 366623
rect 504658 365283 504811 366317
rect 505845 365283 505998 366317
rect 504658 364977 505998 365283
rect 504658 363943 504811 364977
rect 505845 363943 505998 364977
rect 504658 363637 505998 363943
rect 504658 362603 504811 363637
rect 505845 362603 505998 363637
rect 504658 362450 505998 362603
rect 508418 373017 509758 373170
rect 508418 371983 508571 373017
rect 509605 371983 509758 373017
rect 508418 371677 509758 371983
rect 508418 370643 508571 371677
rect 509605 370643 509758 371677
rect 508418 370337 509758 370643
rect 508418 369303 508571 370337
rect 509605 369303 509758 370337
rect 508418 368997 509758 369303
rect 508418 367963 508571 368997
rect 509605 367963 509758 368997
rect 508418 367657 509758 367963
rect 508418 366623 508571 367657
rect 509605 366623 509758 367657
rect 508418 366317 509758 366623
rect 508418 365283 508571 366317
rect 509605 365283 509758 366317
rect 508418 364977 509758 365283
rect 508418 363943 508571 364977
rect 509605 363943 509758 364977
rect 508418 363637 509758 363943
rect 508418 362603 508571 363637
rect 509605 362603 509758 363637
rect 508418 362450 509758 362603
rect 512178 373017 513518 373170
rect 512178 371983 512331 373017
rect 513365 371983 513518 373017
rect 512178 371677 513518 371983
rect 512178 370643 512331 371677
rect 513365 370643 513518 371677
rect 512178 370337 513518 370643
rect 516552 370518 516784 371186
rect 512178 369303 512331 370337
rect 513365 369303 513518 370337
rect 512178 368997 513518 369303
rect 512178 367963 512331 368997
rect 513365 367963 513518 368997
rect 512178 367657 513518 367963
rect 516552 367774 516784 368442
rect 512178 366623 512331 367657
rect 513365 366623 513518 367657
rect 512178 366317 513518 366623
rect 512178 365283 512331 366317
rect 513365 365283 513518 366317
rect 512178 364977 513518 365283
rect 516552 365030 516784 365698
rect 520312 365030 520544 365698
rect 512178 363943 512331 364977
rect 513365 363943 513518 364977
rect 512178 363637 513518 363943
rect 512178 362603 512331 363637
rect 513365 362603 513518 363637
rect 512178 362450 513518 362603
rect 527832 369538 528064 370206
rect 531592 369636 531824 370304
rect 535352 368852 535584 369520
rect 527832 366794 528064 367462
rect 531592 366892 531824 367560
rect 535352 366108 535584 366776
rect 527832 364050 528064 364718
rect 531592 364148 531824 364816
rect 535352 363364 535584 364032
rect 560542 357510 565856 359006
rect 564892 357480 565856 357510
rect 560404 311202 565718 312698
rect 564754 311172 565718 311202
<< nbase >>
rect 504811 401775 505845 402809
rect 497291 370807 498325 371841
rect 497291 369467 498325 370501
rect 497291 368127 498325 369161
rect 497291 366787 498325 367821
rect 497291 365447 498325 366481
rect 497291 364107 498325 365141
rect 497291 362767 498325 363801
rect 501051 371983 502085 373017
rect 501051 370643 502085 371677
rect 501051 369303 502085 370337
rect 501051 367963 502085 368997
rect 501051 366623 502085 367657
rect 501051 365283 502085 366317
rect 501051 363943 502085 364977
rect 501051 362603 502085 363637
rect 504811 371983 505845 373017
rect 504811 370643 505845 371677
rect 504811 369303 505845 370337
rect 504811 367963 505845 368997
rect 504811 366623 505845 367657
rect 504811 365283 505845 366317
rect 504811 363943 505845 364977
rect 504811 362603 505845 363637
rect 508571 371983 509605 373017
rect 508571 370643 509605 371677
rect 508571 369303 509605 370337
rect 508571 367963 509605 368997
rect 508571 366623 509605 367657
rect 508571 365283 509605 366317
rect 508571 363943 509605 364977
rect 508571 362603 509605 363637
rect 512331 371983 513365 373017
rect 512331 370643 513365 371677
rect 512331 369303 513365 370337
rect 512331 367963 513365 368997
rect 512331 366623 513365 367657
rect 512331 365283 513365 366317
rect 512331 363943 513365 364977
rect 512331 362603 513365 363637
<< pmoslvt >>
rect 575263 492214 575463 493214
rect 575521 492214 575721 493214
rect 575779 492214 575979 493214
rect 576037 492214 576237 493214
rect 576295 492214 576495 493214
rect 576553 492214 576753 493214
rect 576811 492214 577011 493214
rect 577069 492214 577269 493214
rect 577327 492214 577527 493214
rect 577585 492214 577785 493214
rect 577843 492214 578043 493214
rect 578101 492214 578301 493214
rect 578359 492214 578559 493214
rect 578617 492214 578817 493214
rect 578875 492214 579075 493214
rect 579133 492214 579333 493214
rect 579391 492214 579591 493214
rect 579649 492214 579849 493214
rect 579907 492214 580107 493214
rect 580165 492214 580365 493214
rect 574541 403338 574741 404338
rect 574799 403338 574999 404338
rect 575057 403338 575257 404338
rect 575315 403338 575515 404338
rect 575573 403338 575773 404338
rect 575831 403338 576031 404338
rect 576089 403338 576289 404338
rect 576347 403338 576547 404338
rect 576605 403338 576805 404338
rect 576863 403338 577063 404338
rect 577121 403338 577321 404338
rect 577379 403338 577579 404338
rect 577637 403338 577837 404338
rect 577895 403338 578095 404338
rect 578153 403338 578353 404338
rect 578411 403338 578611 404338
rect 578669 403338 578869 404338
rect 578927 403338 579127 404338
rect 579185 403338 579385 404338
rect 579443 403338 579643 404338
rect 497103 399431 498393 399831
rect 497103 398973 498393 399373
rect 497103 398515 498393 398915
rect 497103 398057 498393 398457
rect 497103 397599 498393 397999
rect 497103 397141 498393 397541
rect 497103 396683 498393 397083
rect 497103 396225 498393 396625
rect 497103 395767 498393 396167
rect 497103 395309 498393 395709
rect 497103 394851 498393 395251
rect 497103 394393 498393 394793
rect 497103 393935 498393 394335
rect 497103 393477 498393 393877
rect 497103 393019 498393 393419
rect 497103 392561 498393 392961
rect 497103 392103 498393 392503
rect 497103 391645 498393 392045
rect 500863 391787 502153 392187
rect 497103 391187 498393 391587
rect 500863 391329 502153 391729
rect 497103 390729 498393 391129
rect 497103 390271 498393 390671
rect 500863 390871 502153 391271
rect 493343 389631 494633 390031
rect 493343 389173 494633 389573
rect 497103 389813 498393 390213
rect 500863 390413 502153 390813
rect 497103 389355 498393 389755
rect 500863 389955 502153 390355
rect 500863 389497 502153 389897
rect 493343 388715 494633 389115
rect 497103 388897 498393 389297
rect 500863 389039 502153 389439
rect 493343 388257 494633 388657
rect 497103 388439 498393 388839
rect 500863 388581 502153 388981
rect 493343 387799 494633 388199
rect 497103 387981 498393 388381
rect 500863 388123 502153 388523
rect 493343 387341 494633 387741
rect 497103 387523 498393 387923
rect 523423 389631 524713 390031
rect 523423 389173 524713 389573
rect 523423 388715 524713 389115
rect 493343 386883 494633 387283
rect 497103 387065 498393 387465
rect 500863 387665 502153 388065
rect 523423 388257 524713 388657
rect 493343 386425 494633 386825
rect 497103 386607 498393 387007
rect 500863 387207 502153 387607
rect 493343 385967 494633 386367
rect 497103 386149 498393 386549
rect 500863 386749 502153 387149
rect 493343 385509 494633 385909
rect 497103 385691 498393 386091
rect 493343 385051 494633 385451
rect 497103 385233 498393 385633
rect 493343 384593 494633 384993
rect 497103 384775 498393 385175
rect 500863 385123 502153 385523
rect 523423 387799 524713 388199
rect 523423 387341 524713 387741
rect 523423 386883 524713 387283
rect 523423 386425 524713 386825
rect 523423 385967 524713 386367
rect 523423 385509 524713 385909
rect 493343 384135 494633 384535
rect 497103 384317 498393 384717
rect 500863 384665 502153 385065
rect 523423 385051 524713 385451
rect 493343 383677 494633 384077
rect 497103 383859 498393 384259
rect 500863 384207 502153 384607
rect 493343 383219 494633 383619
rect 497103 383401 498393 383801
rect 500863 383749 502153 384149
rect 493343 382761 494633 383161
rect 497103 382943 498393 383343
rect 500863 383291 502153 383691
rect 493343 382303 494633 382703
rect 497103 382485 498393 382885
rect 500863 382833 502153 383233
rect 493343 381845 494633 382245
rect 497103 382027 498393 382427
rect 500863 382375 502153 382775
rect 523423 384593 524713 384993
rect 523423 384135 524713 384535
rect 523423 383677 524713 384077
rect 523423 383219 524713 383619
rect 523423 382761 524713 383161
rect 493343 381387 494633 381787
rect 497103 381569 498393 381969
rect 500863 381917 502153 382317
rect 523423 382303 524713 382703
rect 493343 380929 494633 381329
rect 497103 381111 498393 381511
rect 500863 381459 502153 381859
rect 523423 381845 524713 382245
rect 493343 380471 494633 380871
rect 493343 380013 494633 380413
rect 497103 380653 498393 381053
rect 500863 381001 502153 381401
rect 497103 380195 498393 380595
rect 500863 380543 502153 380943
rect 493343 379555 494633 379955
rect 497103 379737 498393 380137
rect 500863 380085 502153 380485
rect 493343 379097 494633 379497
rect 497103 379279 498393 379679
rect 523423 381387 524713 381787
rect 523423 380929 524713 381329
rect 523423 380471 524713 380871
rect 523423 380013 524713 380413
rect 523423 379555 524713 379955
rect 493343 378639 494633 379039
rect 497103 378821 498393 379221
rect 523423 379097 524713 379497
rect 493343 378181 494633 378581
rect 497103 378363 498393 378763
rect 523423 378639 524713 379039
rect 493343 377723 494633 378123
rect 493343 377265 494633 377665
rect 497103 377905 498393 378305
rect 523423 378181 524713 378581
rect 493343 376807 494633 377207
rect 497103 377447 498393 377847
rect 523423 377723 524713 378123
rect 493343 376349 494633 376749
rect 497103 376989 498393 377389
rect 497103 376531 498393 376931
rect 504623 376989 505913 377389
rect 493343 375891 494633 376291
rect 497103 376073 498393 376473
rect 504623 376531 505913 376931
rect 512143 376989 513433 377389
rect 512143 376531 513433 376931
rect 493343 375433 494633 375833
rect 497103 375615 498393 376015
rect 504623 376073 505913 376473
rect 512143 376073 513433 376473
rect 493343 374975 494633 375375
rect 497103 375157 498393 375557
rect 504623 375615 505913 376015
rect 493343 374517 494633 374917
rect 493343 374059 494633 374459
rect 497103 374699 498393 375099
rect 504623 375157 505913 375557
rect 512143 375615 513433 376015
rect 493343 373601 494633 374001
rect 497103 374241 498393 374641
rect 493343 373143 494633 373543
rect 497103 373783 498393 374183
rect 504623 374699 505913 375099
rect 512143 375157 513433 375557
rect 512143 374699 513433 375099
rect 523423 377265 524713 377665
rect 523423 376807 524713 377207
rect 523423 376349 524713 376749
rect 523423 375891 524713 376291
rect 523423 375433 524713 375833
rect 523423 374975 524713 375375
rect 497103 373325 498393 373725
rect 493343 372685 494633 373085
rect 497103 372867 498393 373267
rect 493343 372227 494633 372627
rect 497103 372409 498393 372809
rect 493343 371769 494633 372169
rect 493343 371311 494633 371711
rect 493343 370853 494633 371253
rect 493343 370395 494633 370795
rect 493343 369937 494633 370337
rect 493343 369479 494633 369879
rect 493343 369021 494633 369421
rect 493343 368563 494633 368963
rect 493343 368105 494633 368505
rect 493343 367647 494633 368047
rect 493343 367189 494633 367589
rect 493343 366731 494633 367131
rect 493343 366273 494633 366673
rect 493343 365815 494633 366215
rect 493343 365357 494633 365757
rect 493343 364899 494633 365299
rect 493343 364441 494633 364841
rect 493343 363983 494633 364383
rect 493343 363525 494633 363925
rect 493343 363067 494633 363467
rect 493343 362609 494633 363009
rect 523423 374517 524713 374917
rect 523423 374059 524713 374459
rect 523423 373601 524713 374001
rect 523423 373143 524713 373543
rect 523423 372685 524713 373085
rect 523423 372227 524713 372627
rect 523423 371769 524713 372169
rect 523423 371311 524713 371711
rect 523423 370853 524713 371253
rect 523423 370395 524713 370795
rect 523423 369937 524713 370337
rect 523423 369479 524713 369879
rect 523423 369021 524713 369421
rect 523423 368563 524713 368963
rect 523423 368105 524713 368505
rect 523423 367647 524713 368047
rect 523423 367189 524713 367589
rect 523423 366731 524713 367131
rect 523423 366273 524713 366673
rect 523423 365815 524713 366215
rect 523423 365357 524713 365757
rect 523423 364899 524713 365299
rect 523423 364441 524713 364841
rect 523423 363983 524713 364383
rect 523423 363525 524713 363925
rect 523423 363067 524713 363467
rect 523423 362609 524713 363009
rect 574737 357910 574937 358910
rect 574995 357910 575195 358910
rect 575253 357910 575453 358910
rect 575511 357910 575711 358910
rect 575769 357910 575969 358910
rect 576027 357910 576227 358910
rect 576285 357910 576485 358910
rect 576543 357910 576743 358910
rect 576801 357910 577001 358910
rect 577059 357910 577259 358910
rect 577317 357910 577517 358910
rect 577575 357910 577775 358910
rect 577833 357910 578033 358910
rect 578091 357910 578291 358910
rect 578349 357910 578549 358910
rect 578607 357910 578807 358910
rect 578865 357910 579065 358910
rect 579123 357910 579323 358910
rect 579381 357910 579581 358910
rect 579639 357910 579839 358910
rect 575185 311742 575385 312742
rect 575443 311742 575643 312742
rect 575701 311742 575901 312742
rect 575959 311742 576159 312742
rect 576217 311742 576417 312742
rect 576475 311742 576675 312742
rect 576733 311742 576933 312742
rect 576991 311742 577191 312742
rect 577249 311742 577449 312742
rect 577507 311742 577707 312742
rect 577765 311742 577965 312742
rect 578023 311742 578223 312742
rect 578281 311742 578481 312742
rect 578539 311742 578739 312742
rect 578797 311742 578997 312742
rect 579055 311742 579255 312742
rect 579313 311742 579513 312742
rect 579571 311742 579771 312742
rect 579829 311742 580029 312742
rect 580087 311742 580287 312742
<< nmoslvt >>
rect 560707 492440 560907 493440
rect 560965 492440 561165 493440
rect 561223 492440 561423 493440
rect 561481 492440 561681 493440
rect 561739 492440 561939 493440
rect 561997 492440 562197 493440
rect 562255 492440 562455 493440
rect 562513 492440 562713 493440
rect 562771 492440 562971 493440
rect 563029 492440 563229 493440
rect 563287 492440 563487 493440
rect 563545 492440 563745 493440
rect 563803 492440 564003 493440
rect 564061 492440 564261 493440
rect 564319 492440 564519 493440
rect 564577 492440 564777 493440
rect 564835 492440 565035 493440
rect 565093 492440 565293 493440
rect 565351 492440 565551 493440
rect 565609 492440 565809 493440
rect 560747 403298 560947 404298
rect 561005 403298 561205 404298
rect 561263 403298 561463 404298
rect 561521 403298 561721 404298
rect 561779 403298 561979 404298
rect 562037 403298 562237 404298
rect 562295 403298 562495 404298
rect 562553 403298 562753 404298
rect 562811 403298 563011 404298
rect 563069 403298 563269 404298
rect 563327 403298 563527 404298
rect 563585 403298 563785 404298
rect 563843 403298 564043 404298
rect 564101 403298 564301 404298
rect 564359 403298 564559 404298
rect 564617 403298 564817 404298
rect 564875 403298 565075 404298
rect 565133 403298 565333 404298
rect 565391 403298 565591 404298
rect 565649 403298 565849 404298
rect 497348 400378 498148 400778
rect 493588 390578 494388 390978
rect 504868 389078 505668 389478
rect 504868 388620 505668 389020
rect 516148 389078 516948 389478
rect 504868 388162 505668 388562
rect 516148 388620 516948 389020
rect 516148 388162 516948 388562
rect 504868 387704 505668 388104
rect 504868 387246 505668 387646
rect 504868 386788 505668 387188
rect 504868 386330 505668 386730
rect 504868 385872 505668 386272
rect 504868 385414 505668 385814
rect 516148 387704 516948 388104
rect 516148 387246 516948 387646
rect 516148 386788 516948 387188
rect 516148 386330 516948 386730
rect 516148 385872 516948 386272
rect 516148 385414 516948 385814
rect 501108 377220 501908 377620
rect 501108 376762 501908 377162
rect 501108 376304 501908 376704
rect 501108 375846 501908 376246
rect 501108 375388 501908 375788
rect 501108 374930 501908 375330
rect 501108 374472 501908 374872
rect 501108 374014 501908 374414
rect 501108 373556 501908 373956
rect 560599 357980 560799 358980
rect 560857 357980 561057 358980
rect 561115 357980 561315 358980
rect 561373 357980 561573 358980
rect 561631 357980 561831 358980
rect 561889 357980 562089 358980
rect 562147 357980 562347 358980
rect 562405 357980 562605 358980
rect 562663 357980 562863 358980
rect 562921 357980 563121 358980
rect 563179 357980 563379 358980
rect 563437 357980 563637 358980
rect 563695 357980 563895 358980
rect 563953 357980 564153 358980
rect 564211 357980 564411 358980
rect 564469 357980 564669 358980
rect 564727 357980 564927 358980
rect 564985 357980 565185 358980
rect 565243 357980 565443 358980
rect 565501 357980 565701 358980
rect 560461 311672 560661 312672
rect 560719 311672 560919 312672
rect 560977 311672 561177 312672
rect 561235 311672 561435 312672
rect 561493 311672 561693 312672
rect 561751 311672 561951 312672
rect 562009 311672 562209 312672
rect 562267 311672 562467 312672
rect 562525 311672 562725 312672
rect 562783 311672 562983 312672
rect 563041 311672 563241 312672
rect 563299 311672 563499 312672
rect 563557 311672 563757 312672
rect 563815 311672 564015 312672
rect 564073 311672 564273 312672
rect 564331 311672 564531 312672
rect 564589 311672 564789 312672
rect 564847 311672 565047 312672
rect 565105 311672 565305 312672
rect 565363 311672 565563 312672
<< ndiff >>
rect 560649 493428 560707 493440
rect 560649 492452 560661 493428
rect 560695 492452 560707 493428
rect 560649 492440 560707 492452
rect 560907 493428 560965 493440
rect 560907 492452 560919 493428
rect 560953 492452 560965 493428
rect 560907 492440 560965 492452
rect 561165 493428 561223 493440
rect 561165 492452 561177 493428
rect 561211 492452 561223 493428
rect 561165 492440 561223 492452
rect 561423 493428 561481 493440
rect 561423 492452 561435 493428
rect 561469 492452 561481 493428
rect 561423 492440 561481 492452
rect 561681 493428 561739 493440
rect 561681 492452 561693 493428
rect 561727 492452 561739 493428
rect 561681 492440 561739 492452
rect 561939 493428 561997 493440
rect 561939 492452 561951 493428
rect 561985 492452 561997 493428
rect 561939 492440 561997 492452
rect 562197 493428 562255 493440
rect 562197 492452 562209 493428
rect 562243 492452 562255 493428
rect 562197 492440 562255 492452
rect 562455 493428 562513 493440
rect 562455 492452 562467 493428
rect 562501 492452 562513 493428
rect 562455 492440 562513 492452
rect 562713 493428 562771 493440
rect 562713 492452 562725 493428
rect 562759 492452 562771 493428
rect 562713 492440 562771 492452
rect 562971 493428 563029 493440
rect 562971 492452 562983 493428
rect 563017 492452 563029 493428
rect 562971 492440 563029 492452
rect 563229 493428 563287 493440
rect 563229 492452 563241 493428
rect 563275 492452 563287 493428
rect 563229 492440 563287 492452
rect 563487 493428 563545 493440
rect 563487 492452 563499 493428
rect 563533 492452 563545 493428
rect 563487 492440 563545 492452
rect 563745 493428 563803 493440
rect 563745 492452 563757 493428
rect 563791 492452 563803 493428
rect 563745 492440 563803 492452
rect 564003 493428 564061 493440
rect 564003 492452 564015 493428
rect 564049 492452 564061 493428
rect 564003 492440 564061 492452
rect 564261 493428 564319 493440
rect 564261 492452 564273 493428
rect 564307 492452 564319 493428
rect 564261 492440 564319 492452
rect 564519 493428 564577 493440
rect 564519 492452 564531 493428
rect 564565 492452 564577 493428
rect 564519 492440 564577 492452
rect 564777 493428 564835 493440
rect 564777 492452 564789 493428
rect 564823 492452 564835 493428
rect 564777 492440 564835 492452
rect 565035 493428 565093 493440
rect 565035 492452 565047 493428
rect 565081 492452 565093 493428
rect 565035 492440 565093 492452
rect 565293 493428 565351 493440
rect 565293 492452 565305 493428
rect 565339 492452 565351 493428
rect 565293 492440 565351 492452
rect 565551 493428 565609 493440
rect 565551 492452 565563 493428
rect 565597 492452 565609 493428
rect 565551 492440 565609 492452
rect 565809 493428 565867 493440
rect 565809 492452 565821 493428
rect 565855 492452 565867 493428
rect 565809 492440 565867 492452
rect 560689 404286 560747 404298
rect 560689 403310 560701 404286
rect 560735 403310 560747 404286
rect 560689 403298 560747 403310
rect 560947 404286 561005 404298
rect 560947 403310 560959 404286
rect 560993 403310 561005 404286
rect 560947 403298 561005 403310
rect 561205 404286 561263 404298
rect 561205 403310 561217 404286
rect 561251 403310 561263 404286
rect 561205 403298 561263 403310
rect 561463 404286 561521 404298
rect 561463 403310 561475 404286
rect 561509 403310 561521 404286
rect 561463 403298 561521 403310
rect 561721 404286 561779 404298
rect 561721 403310 561733 404286
rect 561767 403310 561779 404286
rect 561721 403298 561779 403310
rect 561979 404286 562037 404298
rect 561979 403310 561991 404286
rect 562025 403310 562037 404286
rect 561979 403298 562037 403310
rect 562237 404286 562295 404298
rect 562237 403310 562249 404286
rect 562283 403310 562295 404286
rect 562237 403298 562295 403310
rect 562495 404286 562553 404298
rect 562495 403310 562507 404286
rect 562541 403310 562553 404286
rect 562495 403298 562553 403310
rect 562753 404286 562811 404298
rect 562753 403310 562765 404286
rect 562799 403310 562811 404286
rect 562753 403298 562811 403310
rect 563011 404286 563069 404298
rect 563011 403310 563023 404286
rect 563057 403310 563069 404286
rect 563011 403298 563069 403310
rect 563269 404286 563327 404298
rect 563269 403310 563281 404286
rect 563315 403310 563327 404286
rect 563269 403298 563327 403310
rect 563527 404286 563585 404298
rect 563527 403310 563539 404286
rect 563573 403310 563585 404286
rect 563527 403298 563585 403310
rect 563785 404286 563843 404298
rect 563785 403310 563797 404286
rect 563831 403310 563843 404286
rect 563785 403298 563843 403310
rect 564043 404286 564101 404298
rect 564043 403310 564055 404286
rect 564089 403310 564101 404286
rect 564043 403298 564101 403310
rect 564301 404286 564359 404298
rect 564301 403310 564313 404286
rect 564347 403310 564359 404286
rect 564301 403298 564359 403310
rect 564559 404286 564617 404298
rect 564559 403310 564571 404286
rect 564605 403310 564617 404286
rect 564559 403298 564617 403310
rect 564817 404286 564875 404298
rect 564817 403310 564829 404286
rect 564863 403310 564875 404286
rect 564817 403298 564875 403310
rect 565075 404286 565133 404298
rect 565075 403310 565087 404286
rect 565121 403310 565133 404286
rect 565075 403298 565133 403310
rect 565333 404286 565391 404298
rect 565333 403310 565345 404286
rect 565379 403310 565391 404286
rect 565333 403298 565391 403310
rect 565591 404286 565649 404298
rect 565591 403310 565603 404286
rect 565637 403310 565649 404286
rect 565591 403298 565649 403310
rect 565849 404286 565907 404298
rect 565849 403310 565861 404286
rect 565895 403310 565907 404286
rect 565849 403298 565907 403310
rect 497348 400824 498148 400836
rect 497348 400790 497391 400824
rect 497425 400790 497459 400824
rect 497493 400790 497527 400824
rect 497561 400790 497595 400824
rect 497629 400790 497663 400824
rect 497697 400790 497731 400824
rect 497765 400790 497799 400824
rect 497833 400790 497867 400824
rect 497901 400790 497935 400824
rect 497969 400790 498003 400824
rect 498037 400790 498071 400824
rect 498105 400790 498148 400824
rect 497348 400778 498148 400790
rect 497348 400366 498148 400378
rect 497348 400332 497391 400366
rect 497425 400332 497459 400366
rect 497493 400332 497527 400366
rect 497561 400332 497595 400366
rect 497629 400332 497663 400366
rect 497697 400332 497731 400366
rect 497765 400332 497799 400366
rect 497833 400332 497867 400366
rect 497901 400332 497935 400366
rect 497969 400332 498003 400366
rect 498037 400332 498071 400366
rect 498105 400332 498148 400366
rect 497348 400320 498148 400332
rect 493588 391024 494388 391036
rect 493588 390990 493631 391024
rect 493665 390990 493699 391024
rect 493733 390990 493767 391024
rect 493801 390990 493835 391024
rect 493869 390990 493903 391024
rect 493937 390990 493971 391024
rect 494005 390990 494039 391024
rect 494073 390990 494107 391024
rect 494141 390990 494175 391024
rect 494209 390990 494243 391024
rect 494277 390990 494311 391024
rect 494345 390990 494388 391024
rect 493588 390978 494388 390990
rect 493588 390566 494388 390578
rect 493588 390532 493631 390566
rect 493665 390532 493699 390566
rect 493733 390532 493767 390566
rect 493801 390532 493835 390566
rect 493869 390532 493903 390566
rect 493937 390532 493971 390566
rect 494005 390532 494039 390566
rect 494073 390532 494107 390566
rect 494141 390532 494175 390566
rect 494209 390532 494243 390566
rect 494277 390532 494311 390566
rect 494345 390532 494388 390566
rect 493588 390520 494388 390532
rect 504868 389524 505668 389536
rect 504868 389490 504911 389524
rect 504945 389490 504979 389524
rect 505013 389490 505047 389524
rect 505081 389490 505115 389524
rect 505149 389490 505183 389524
rect 505217 389490 505251 389524
rect 505285 389490 505319 389524
rect 505353 389490 505387 389524
rect 505421 389490 505455 389524
rect 505489 389490 505523 389524
rect 505557 389490 505591 389524
rect 505625 389490 505668 389524
rect 504868 389478 505668 389490
rect 516148 389524 516948 389536
rect 516148 389490 516191 389524
rect 516225 389490 516259 389524
rect 516293 389490 516327 389524
rect 516361 389490 516395 389524
rect 516429 389490 516463 389524
rect 516497 389490 516531 389524
rect 516565 389490 516599 389524
rect 516633 389490 516667 389524
rect 516701 389490 516735 389524
rect 516769 389490 516803 389524
rect 516837 389490 516871 389524
rect 516905 389490 516948 389524
rect 516148 389478 516948 389490
rect 504868 389066 505668 389078
rect 504868 389032 504911 389066
rect 504945 389032 504979 389066
rect 505013 389032 505047 389066
rect 505081 389032 505115 389066
rect 505149 389032 505183 389066
rect 505217 389032 505251 389066
rect 505285 389032 505319 389066
rect 505353 389032 505387 389066
rect 505421 389032 505455 389066
rect 505489 389032 505523 389066
rect 505557 389032 505591 389066
rect 505625 389032 505668 389066
rect 504868 389020 505668 389032
rect 516148 389066 516948 389078
rect 516148 389032 516191 389066
rect 516225 389032 516259 389066
rect 516293 389032 516327 389066
rect 516361 389032 516395 389066
rect 516429 389032 516463 389066
rect 516497 389032 516531 389066
rect 516565 389032 516599 389066
rect 516633 389032 516667 389066
rect 516701 389032 516735 389066
rect 516769 389032 516803 389066
rect 516837 389032 516871 389066
rect 516905 389032 516948 389066
rect 516148 389020 516948 389032
rect 504868 388608 505668 388620
rect 504868 388574 504911 388608
rect 504945 388574 504979 388608
rect 505013 388574 505047 388608
rect 505081 388574 505115 388608
rect 505149 388574 505183 388608
rect 505217 388574 505251 388608
rect 505285 388574 505319 388608
rect 505353 388574 505387 388608
rect 505421 388574 505455 388608
rect 505489 388574 505523 388608
rect 505557 388574 505591 388608
rect 505625 388574 505668 388608
rect 504868 388562 505668 388574
rect 516148 388608 516948 388620
rect 516148 388574 516191 388608
rect 516225 388574 516259 388608
rect 516293 388574 516327 388608
rect 516361 388574 516395 388608
rect 516429 388574 516463 388608
rect 516497 388574 516531 388608
rect 516565 388574 516599 388608
rect 516633 388574 516667 388608
rect 516701 388574 516735 388608
rect 516769 388574 516803 388608
rect 516837 388574 516871 388608
rect 516905 388574 516948 388608
rect 516148 388562 516948 388574
rect 504868 388150 505668 388162
rect 504868 388116 504911 388150
rect 504945 388116 504979 388150
rect 505013 388116 505047 388150
rect 505081 388116 505115 388150
rect 505149 388116 505183 388150
rect 505217 388116 505251 388150
rect 505285 388116 505319 388150
rect 505353 388116 505387 388150
rect 505421 388116 505455 388150
rect 505489 388116 505523 388150
rect 505557 388116 505591 388150
rect 505625 388116 505668 388150
rect 504868 388104 505668 388116
rect 516148 388150 516948 388162
rect 516148 388116 516191 388150
rect 516225 388116 516259 388150
rect 516293 388116 516327 388150
rect 516361 388116 516395 388150
rect 516429 388116 516463 388150
rect 516497 388116 516531 388150
rect 516565 388116 516599 388150
rect 516633 388116 516667 388150
rect 516701 388116 516735 388150
rect 516769 388116 516803 388150
rect 516837 388116 516871 388150
rect 516905 388116 516948 388150
rect 516148 388104 516948 388116
rect 504868 387692 505668 387704
rect 504868 387658 504911 387692
rect 504945 387658 504979 387692
rect 505013 387658 505047 387692
rect 505081 387658 505115 387692
rect 505149 387658 505183 387692
rect 505217 387658 505251 387692
rect 505285 387658 505319 387692
rect 505353 387658 505387 387692
rect 505421 387658 505455 387692
rect 505489 387658 505523 387692
rect 505557 387658 505591 387692
rect 505625 387658 505668 387692
rect 504868 387646 505668 387658
rect 504868 387234 505668 387246
rect 504868 387200 504911 387234
rect 504945 387200 504979 387234
rect 505013 387200 505047 387234
rect 505081 387200 505115 387234
rect 505149 387200 505183 387234
rect 505217 387200 505251 387234
rect 505285 387200 505319 387234
rect 505353 387200 505387 387234
rect 505421 387200 505455 387234
rect 505489 387200 505523 387234
rect 505557 387200 505591 387234
rect 505625 387200 505668 387234
rect 504868 387188 505668 387200
rect 504868 386776 505668 386788
rect 504868 386742 504911 386776
rect 504945 386742 504979 386776
rect 505013 386742 505047 386776
rect 505081 386742 505115 386776
rect 505149 386742 505183 386776
rect 505217 386742 505251 386776
rect 505285 386742 505319 386776
rect 505353 386742 505387 386776
rect 505421 386742 505455 386776
rect 505489 386742 505523 386776
rect 505557 386742 505591 386776
rect 505625 386742 505668 386776
rect 504868 386730 505668 386742
rect 504868 386318 505668 386330
rect 504868 386284 504911 386318
rect 504945 386284 504979 386318
rect 505013 386284 505047 386318
rect 505081 386284 505115 386318
rect 505149 386284 505183 386318
rect 505217 386284 505251 386318
rect 505285 386284 505319 386318
rect 505353 386284 505387 386318
rect 505421 386284 505455 386318
rect 505489 386284 505523 386318
rect 505557 386284 505591 386318
rect 505625 386284 505668 386318
rect 504868 386272 505668 386284
rect 504868 385860 505668 385872
rect 504868 385826 504911 385860
rect 504945 385826 504979 385860
rect 505013 385826 505047 385860
rect 505081 385826 505115 385860
rect 505149 385826 505183 385860
rect 505217 385826 505251 385860
rect 505285 385826 505319 385860
rect 505353 385826 505387 385860
rect 505421 385826 505455 385860
rect 505489 385826 505523 385860
rect 505557 385826 505591 385860
rect 505625 385826 505668 385860
rect 504868 385814 505668 385826
rect 504868 385402 505668 385414
rect 504868 385368 504911 385402
rect 504945 385368 504979 385402
rect 505013 385368 505047 385402
rect 505081 385368 505115 385402
rect 505149 385368 505183 385402
rect 505217 385368 505251 385402
rect 505285 385368 505319 385402
rect 505353 385368 505387 385402
rect 505421 385368 505455 385402
rect 505489 385368 505523 385402
rect 505557 385368 505591 385402
rect 505625 385368 505668 385402
rect 504868 385356 505668 385368
rect 516148 387692 516948 387704
rect 516148 387658 516191 387692
rect 516225 387658 516259 387692
rect 516293 387658 516327 387692
rect 516361 387658 516395 387692
rect 516429 387658 516463 387692
rect 516497 387658 516531 387692
rect 516565 387658 516599 387692
rect 516633 387658 516667 387692
rect 516701 387658 516735 387692
rect 516769 387658 516803 387692
rect 516837 387658 516871 387692
rect 516905 387658 516948 387692
rect 516148 387646 516948 387658
rect 516148 387234 516948 387246
rect 516148 387200 516191 387234
rect 516225 387200 516259 387234
rect 516293 387200 516327 387234
rect 516361 387200 516395 387234
rect 516429 387200 516463 387234
rect 516497 387200 516531 387234
rect 516565 387200 516599 387234
rect 516633 387200 516667 387234
rect 516701 387200 516735 387234
rect 516769 387200 516803 387234
rect 516837 387200 516871 387234
rect 516905 387200 516948 387234
rect 516148 387188 516948 387200
rect 516148 386776 516948 386788
rect 516148 386742 516191 386776
rect 516225 386742 516259 386776
rect 516293 386742 516327 386776
rect 516361 386742 516395 386776
rect 516429 386742 516463 386776
rect 516497 386742 516531 386776
rect 516565 386742 516599 386776
rect 516633 386742 516667 386776
rect 516701 386742 516735 386776
rect 516769 386742 516803 386776
rect 516837 386742 516871 386776
rect 516905 386742 516948 386776
rect 516148 386730 516948 386742
rect 516148 386318 516948 386330
rect 516148 386284 516191 386318
rect 516225 386284 516259 386318
rect 516293 386284 516327 386318
rect 516361 386284 516395 386318
rect 516429 386284 516463 386318
rect 516497 386284 516531 386318
rect 516565 386284 516599 386318
rect 516633 386284 516667 386318
rect 516701 386284 516735 386318
rect 516769 386284 516803 386318
rect 516837 386284 516871 386318
rect 516905 386284 516948 386318
rect 516148 386272 516948 386284
rect 516148 385860 516948 385872
rect 516148 385826 516191 385860
rect 516225 385826 516259 385860
rect 516293 385826 516327 385860
rect 516361 385826 516395 385860
rect 516429 385826 516463 385860
rect 516497 385826 516531 385860
rect 516565 385826 516599 385860
rect 516633 385826 516667 385860
rect 516701 385826 516735 385860
rect 516769 385826 516803 385860
rect 516837 385826 516871 385860
rect 516905 385826 516948 385860
rect 516148 385814 516948 385826
rect 516148 385402 516948 385414
rect 516148 385368 516191 385402
rect 516225 385368 516259 385402
rect 516293 385368 516327 385402
rect 516361 385368 516395 385402
rect 516429 385368 516463 385402
rect 516497 385368 516531 385402
rect 516565 385368 516599 385402
rect 516633 385368 516667 385402
rect 516701 385368 516735 385402
rect 516769 385368 516803 385402
rect 516837 385368 516871 385402
rect 516905 385368 516948 385402
rect 516148 385356 516948 385368
rect 501108 377666 501908 377678
rect 501108 377632 501151 377666
rect 501185 377632 501219 377666
rect 501253 377632 501287 377666
rect 501321 377632 501355 377666
rect 501389 377632 501423 377666
rect 501457 377632 501491 377666
rect 501525 377632 501559 377666
rect 501593 377632 501627 377666
rect 501661 377632 501695 377666
rect 501729 377632 501763 377666
rect 501797 377632 501831 377666
rect 501865 377632 501908 377666
rect 501108 377620 501908 377632
rect 501108 377208 501908 377220
rect 501108 377174 501151 377208
rect 501185 377174 501219 377208
rect 501253 377174 501287 377208
rect 501321 377174 501355 377208
rect 501389 377174 501423 377208
rect 501457 377174 501491 377208
rect 501525 377174 501559 377208
rect 501593 377174 501627 377208
rect 501661 377174 501695 377208
rect 501729 377174 501763 377208
rect 501797 377174 501831 377208
rect 501865 377174 501908 377208
rect 501108 377162 501908 377174
rect 501108 376750 501908 376762
rect 501108 376716 501151 376750
rect 501185 376716 501219 376750
rect 501253 376716 501287 376750
rect 501321 376716 501355 376750
rect 501389 376716 501423 376750
rect 501457 376716 501491 376750
rect 501525 376716 501559 376750
rect 501593 376716 501627 376750
rect 501661 376716 501695 376750
rect 501729 376716 501763 376750
rect 501797 376716 501831 376750
rect 501865 376716 501908 376750
rect 501108 376704 501908 376716
rect 501108 376292 501908 376304
rect 501108 376258 501151 376292
rect 501185 376258 501219 376292
rect 501253 376258 501287 376292
rect 501321 376258 501355 376292
rect 501389 376258 501423 376292
rect 501457 376258 501491 376292
rect 501525 376258 501559 376292
rect 501593 376258 501627 376292
rect 501661 376258 501695 376292
rect 501729 376258 501763 376292
rect 501797 376258 501831 376292
rect 501865 376258 501908 376292
rect 501108 376246 501908 376258
rect 501108 375834 501908 375846
rect 501108 375800 501151 375834
rect 501185 375800 501219 375834
rect 501253 375800 501287 375834
rect 501321 375800 501355 375834
rect 501389 375800 501423 375834
rect 501457 375800 501491 375834
rect 501525 375800 501559 375834
rect 501593 375800 501627 375834
rect 501661 375800 501695 375834
rect 501729 375800 501763 375834
rect 501797 375800 501831 375834
rect 501865 375800 501908 375834
rect 501108 375788 501908 375800
rect 501108 375376 501908 375388
rect 501108 375342 501151 375376
rect 501185 375342 501219 375376
rect 501253 375342 501287 375376
rect 501321 375342 501355 375376
rect 501389 375342 501423 375376
rect 501457 375342 501491 375376
rect 501525 375342 501559 375376
rect 501593 375342 501627 375376
rect 501661 375342 501695 375376
rect 501729 375342 501763 375376
rect 501797 375342 501831 375376
rect 501865 375342 501908 375376
rect 501108 375330 501908 375342
rect 501108 374918 501908 374930
rect 501108 374884 501151 374918
rect 501185 374884 501219 374918
rect 501253 374884 501287 374918
rect 501321 374884 501355 374918
rect 501389 374884 501423 374918
rect 501457 374884 501491 374918
rect 501525 374884 501559 374918
rect 501593 374884 501627 374918
rect 501661 374884 501695 374918
rect 501729 374884 501763 374918
rect 501797 374884 501831 374918
rect 501865 374884 501908 374918
rect 501108 374872 501908 374884
rect 501108 374460 501908 374472
rect 501108 374426 501151 374460
rect 501185 374426 501219 374460
rect 501253 374426 501287 374460
rect 501321 374426 501355 374460
rect 501389 374426 501423 374460
rect 501457 374426 501491 374460
rect 501525 374426 501559 374460
rect 501593 374426 501627 374460
rect 501661 374426 501695 374460
rect 501729 374426 501763 374460
rect 501797 374426 501831 374460
rect 501865 374426 501908 374460
rect 501108 374414 501908 374426
rect 501108 374002 501908 374014
rect 501108 373968 501151 374002
rect 501185 373968 501219 374002
rect 501253 373968 501287 374002
rect 501321 373968 501355 374002
rect 501389 373968 501423 374002
rect 501457 373968 501491 374002
rect 501525 373968 501559 374002
rect 501593 373968 501627 374002
rect 501661 373968 501695 374002
rect 501729 373968 501763 374002
rect 501797 373968 501831 374002
rect 501865 373968 501908 374002
rect 501108 373956 501908 373968
rect 501108 373544 501908 373556
rect 501108 373510 501151 373544
rect 501185 373510 501219 373544
rect 501253 373510 501287 373544
rect 501321 373510 501355 373544
rect 501389 373510 501423 373544
rect 501457 373510 501491 373544
rect 501525 373510 501559 373544
rect 501593 373510 501627 373544
rect 501661 373510 501695 373544
rect 501729 373510 501763 373544
rect 501797 373510 501831 373544
rect 501865 373510 501908 373544
rect 501108 373498 501908 373510
rect 560541 358968 560599 358980
rect 560541 357992 560553 358968
rect 560587 357992 560599 358968
rect 560541 357980 560599 357992
rect 560799 358968 560857 358980
rect 560799 357992 560811 358968
rect 560845 357992 560857 358968
rect 560799 357980 560857 357992
rect 561057 358968 561115 358980
rect 561057 357992 561069 358968
rect 561103 357992 561115 358968
rect 561057 357980 561115 357992
rect 561315 358968 561373 358980
rect 561315 357992 561327 358968
rect 561361 357992 561373 358968
rect 561315 357980 561373 357992
rect 561573 358968 561631 358980
rect 561573 357992 561585 358968
rect 561619 357992 561631 358968
rect 561573 357980 561631 357992
rect 561831 358968 561889 358980
rect 561831 357992 561843 358968
rect 561877 357992 561889 358968
rect 561831 357980 561889 357992
rect 562089 358968 562147 358980
rect 562089 357992 562101 358968
rect 562135 357992 562147 358968
rect 562089 357980 562147 357992
rect 562347 358968 562405 358980
rect 562347 357992 562359 358968
rect 562393 357992 562405 358968
rect 562347 357980 562405 357992
rect 562605 358968 562663 358980
rect 562605 357992 562617 358968
rect 562651 357992 562663 358968
rect 562605 357980 562663 357992
rect 562863 358968 562921 358980
rect 562863 357992 562875 358968
rect 562909 357992 562921 358968
rect 562863 357980 562921 357992
rect 563121 358968 563179 358980
rect 563121 357992 563133 358968
rect 563167 357992 563179 358968
rect 563121 357980 563179 357992
rect 563379 358968 563437 358980
rect 563379 357992 563391 358968
rect 563425 357992 563437 358968
rect 563379 357980 563437 357992
rect 563637 358968 563695 358980
rect 563637 357992 563649 358968
rect 563683 357992 563695 358968
rect 563637 357980 563695 357992
rect 563895 358968 563953 358980
rect 563895 357992 563907 358968
rect 563941 357992 563953 358968
rect 563895 357980 563953 357992
rect 564153 358968 564211 358980
rect 564153 357992 564165 358968
rect 564199 357992 564211 358968
rect 564153 357980 564211 357992
rect 564411 358968 564469 358980
rect 564411 357992 564423 358968
rect 564457 357992 564469 358968
rect 564411 357980 564469 357992
rect 564669 358968 564727 358980
rect 564669 357992 564681 358968
rect 564715 357992 564727 358968
rect 564669 357980 564727 357992
rect 564927 358968 564985 358980
rect 564927 357992 564939 358968
rect 564973 357992 564985 358968
rect 564927 357980 564985 357992
rect 565185 358968 565243 358980
rect 565185 357992 565197 358968
rect 565231 357992 565243 358968
rect 565185 357980 565243 357992
rect 565443 358968 565501 358980
rect 565443 357992 565455 358968
rect 565489 357992 565501 358968
rect 565443 357980 565501 357992
rect 565701 358968 565759 358980
rect 565701 357992 565713 358968
rect 565747 357992 565759 358968
rect 565701 357980 565759 357992
rect 560403 312660 560461 312672
rect 560403 311684 560415 312660
rect 560449 311684 560461 312660
rect 560403 311672 560461 311684
rect 560661 312660 560719 312672
rect 560661 311684 560673 312660
rect 560707 311684 560719 312660
rect 560661 311672 560719 311684
rect 560919 312660 560977 312672
rect 560919 311684 560931 312660
rect 560965 311684 560977 312660
rect 560919 311672 560977 311684
rect 561177 312660 561235 312672
rect 561177 311684 561189 312660
rect 561223 311684 561235 312660
rect 561177 311672 561235 311684
rect 561435 312660 561493 312672
rect 561435 311684 561447 312660
rect 561481 311684 561493 312660
rect 561435 311672 561493 311684
rect 561693 312660 561751 312672
rect 561693 311684 561705 312660
rect 561739 311684 561751 312660
rect 561693 311672 561751 311684
rect 561951 312660 562009 312672
rect 561951 311684 561963 312660
rect 561997 311684 562009 312660
rect 561951 311672 562009 311684
rect 562209 312660 562267 312672
rect 562209 311684 562221 312660
rect 562255 311684 562267 312660
rect 562209 311672 562267 311684
rect 562467 312660 562525 312672
rect 562467 311684 562479 312660
rect 562513 311684 562525 312660
rect 562467 311672 562525 311684
rect 562725 312660 562783 312672
rect 562725 311684 562737 312660
rect 562771 311684 562783 312660
rect 562725 311672 562783 311684
rect 562983 312660 563041 312672
rect 562983 311684 562995 312660
rect 563029 311684 563041 312660
rect 562983 311672 563041 311684
rect 563241 312660 563299 312672
rect 563241 311684 563253 312660
rect 563287 311684 563299 312660
rect 563241 311672 563299 311684
rect 563499 312660 563557 312672
rect 563499 311684 563511 312660
rect 563545 311684 563557 312660
rect 563499 311672 563557 311684
rect 563757 312660 563815 312672
rect 563757 311684 563769 312660
rect 563803 311684 563815 312660
rect 563757 311672 563815 311684
rect 564015 312660 564073 312672
rect 564015 311684 564027 312660
rect 564061 311684 564073 312660
rect 564015 311672 564073 311684
rect 564273 312660 564331 312672
rect 564273 311684 564285 312660
rect 564319 311684 564331 312660
rect 564273 311672 564331 311684
rect 564531 312660 564589 312672
rect 564531 311684 564543 312660
rect 564577 311684 564589 312660
rect 564531 311672 564589 311684
rect 564789 312660 564847 312672
rect 564789 311684 564801 312660
rect 564835 311684 564847 312660
rect 564789 311672 564847 311684
rect 565047 312660 565105 312672
rect 565047 311684 565059 312660
rect 565093 311684 565105 312660
rect 565047 311672 565105 311684
rect 565305 312660 565363 312672
rect 565305 311684 565317 312660
rect 565351 311684 565363 312660
rect 565305 311672 565363 311684
rect 565563 312660 565621 312672
rect 565563 311684 565575 312660
rect 565609 311684 565621 312660
rect 565563 311672 565621 311684
<< pdiff >>
rect 575205 493202 575263 493214
rect 575205 492226 575217 493202
rect 575251 492226 575263 493202
rect 575205 492214 575263 492226
rect 575463 493202 575521 493214
rect 575463 492226 575475 493202
rect 575509 492226 575521 493202
rect 575463 492214 575521 492226
rect 575721 493202 575779 493214
rect 575721 492226 575733 493202
rect 575767 492226 575779 493202
rect 575721 492214 575779 492226
rect 575979 493202 576037 493214
rect 575979 492226 575991 493202
rect 576025 492226 576037 493202
rect 575979 492214 576037 492226
rect 576237 493202 576295 493214
rect 576237 492226 576249 493202
rect 576283 492226 576295 493202
rect 576237 492214 576295 492226
rect 576495 493202 576553 493214
rect 576495 492226 576507 493202
rect 576541 492226 576553 493202
rect 576495 492214 576553 492226
rect 576753 493202 576811 493214
rect 576753 492226 576765 493202
rect 576799 492226 576811 493202
rect 576753 492214 576811 492226
rect 577011 493202 577069 493214
rect 577011 492226 577023 493202
rect 577057 492226 577069 493202
rect 577011 492214 577069 492226
rect 577269 493202 577327 493214
rect 577269 492226 577281 493202
rect 577315 492226 577327 493202
rect 577269 492214 577327 492226
rect 577527 493202 577585 493214
rect 577527 492226 577539 493202
rect 577573 492226 577585 493202
rect 577527 492214 577585 492226
rect 577785 493202 577843 493214
rect 577785 492226 577797 493202
rect 577831 492226 577843 493202
rect 577785 492214 577843 492226
rect 578043 493202 578101 493214
rect 578043 492226 578055 493202
rect 578089 492226 578101 493202
rect 578043 492214 578101 492226
rect 578301 493202 578359 493214
rect 578301 492226 578313 493202
rect 578347 492226 578359 493202
rect 578301 492214 578359 492226
rect 578559 493202 578617 493214
rect 578559 492226 578571 493202
rect 578605 492226 578617 493202
rect 578559 492214 578617 492226
rect 578817 493202 578875 493214
rect 578817 492226 578829 493202
rect 578863 492226 578875 493202
rect 578817 492214 578875 492226
rect 579075 493202 579133 493214
rect 579075 492226 579087 493202
rect 579121 492226 579133 493202
rect 579075 492214 579133 492226
rect 579333 493202 579391 493214
rect 579333 492226 579345 493202
rect 579379 492226 579391 493202
rect 579333 492214 579391 492226
rect 579591 493202 579649 493214
rect 579591 492226 579603 493202
rect 579637 492226 579649 493202
rect 579591 492214 579649 492226
rect 579849 493202 579907 493214
rect 579849 492226 579861 493202
rect 579895 492226 579907 493202
rect 579849 492214 579907 492226
rect 580107 493202 580165 493214
rect 580107 492226 580119 493202
rect 580153 492226 580165 493202
rect 580107 492214 580165 492226
rect 580365 493202 580423 493214
rect 580365 492226 580377 493202
rect 580411 492226 580423 493202
rect 580365 492214 580423 492226
rect 574483 404326 574541 404338
rect 574483 403350 574495 404326
rect 574529 403350 574541 404326
rect 574483 403338 574541 403350
rect 574741 404326 574799 404338
rect 574741 403350 574753 404326
rect 574787 403350 574799 404326
rect 574741 403338 574799 403350
rect 574999 404326 575057 404338
rect 574999 403350 575011 404326
rect 575045 403350 575057 404326
rect 574999 403338 575057 403350
rect 575257 404326 575315 404338
rect 575257 403350 575269 404326
rect 575303 403350 575315 404326
rect 575257 403338 575315 403350
rect 575515 404326 575573 404338
rect 575515 403350 575527 404326
rect 575561 403350 575573 404326
rect 575515 403338 575573 403350
rect 575773 404326 575831 404338
rect 575773 403350 575785 404326
rect 575819 403350 575831 404326
rect 575773 403338 575831 403350
rect 576031 404326 576089 404338
rect 576031 403350 576043 404326
rect 576077 403350 576089 404326
rect 576031 403338 576089 403350
rect 576289 404326 576347 404338
rect 576289 403350 576301 404326
rect 576335 403350 576347 404326
rect 576289 403338 576347 403350
rect 576547 404326 576605 404338
rect 576547 403350 576559 404326
rect 576593 403350 576605 404326
rect 576547 403338 576605 403350
rect 576805 404326 576863 404338
rect 576805 403350 576817 404326
rect 576851 403350 576863 404326
rect 576805 403338 576863 403350
rect 577063 404326 577121 404338
rect 577063 403350 577075 404326
rect 577109 403350 577121 404326
rect 577063 403338 577121 403350
rect 577321 404326 577379 404338
rect 577321 403350 577333 404326
rect 577367 403350 577379 404326
rect 577321 403338 577379 403350
rect 577579 404326 577637 404338
rect 577579 403350 577591 404326
rect 577625 403350 577637 404326
rect 577579 403338 577637 403350
rect 577837 404326 577895 404338
rect 577837 403350 577849 404326
rect 577883 403350 577895 404326
rect 577837 403338 577895 403350
rect 578095 404326 578153 404338
rect 578095 403350 578107 404326
rect 578141 403350 578153 404326
rect 578095 403338 578153 403350
rect 578353 404326 578411 404338
rect 578353 403350 578365 404326
rect 578399 403350 578411 404326
rect 578353 403338 578411 403350
rect 578611 404326 578669 404338
rect 578611 403350 578623 404326
rect 578657 403350 578669 404326
rect 578611 403338 578669 403350
rect 578869 404326 578927 404338
rect 578869 403350 578881 404326
rect 578915 403350 578927 404326
rect 578869 403338 578927 403350
rect 579127 404326 579185 404338
rect 579127 403350 579139 404326
rect 579173 403350 579185 404326
rect 579127 403338 579185 403350
rect 579385 404326 579443 404338
rect 579385 403350 579397 404326
rect 579431 403350 579443 404326
rect 579385 403338 579443 403350
rect 579643 404326 579701 404338
rect 579643 403350 579655 404326
rect 579689 403350 579701 404326
rect 579643 403338 579701 403350
rect 504988 402578 505668 402632
rect 504988 402544 505040 402578
rect 505074 402544 505130 402578
rect 505164 402544 505220 402578
rect 505254 402544 505310 402578
rect 505344 402544 505400 402578
rect 505434 402544 505490 402578
rect 505524 402544 505580 402578
rect 505614 402544 505668 402578
rect 504988 402488 505668 402544
rect 504988 402454 505040 402488
rect 505074 402454 505130 402488
rect 505164 402454 505220 402488
rect 505254 402454 505310 402488
rect 505344 402454 505400 402488
rect 505434 402454 505490 402488
rect 505524 402454 505580 402488
rect 505614 402454 505668 402488
rect 504988 402398 505668 402454
rect 504988 402364 505040 402398
rect 505074 402364 505130 402398
rect 505164 402364 505220 402398
rect 505254 402364 505310 402398
rect 505344 402364 505400 402398
rect 505434 402364 505490 402398
rect 505524 402364 505580 402398
rect 505614 402364 505668 402398
rect 504988 402308 505668 402364
rect 504988 402274 505040 402308
rect 505074 402274 505130 402308
rect 505164 402274 505220 402308
rect 505254 402274 505310 402308
rect 505344 402274 505400 402308
rect 505434 402274 505490 402308
rect 505524 402274 505580 402308
rect 505614 402274 505668 402308
rect 504988 402218 505668 402274
rect 504988 402184 505040 402218
rect 505074 402184 505130 402218
rect 505164 402184 505220 402218
rect 505254 402184 505310 402218
rect 505344 402184 505400 402218
rect 505434 402184 505490 402218
rect 505524 402184 505580 402218
rect 505614 402184 505668 402218
rect 504988 402128 505668 402184
rect 504988 402094 505040 402128
rect 505074 402094 505130 402128
rect 505164 402094 505220 402128
rect 505254 402094 505310 402128
rect 505344 402094 505400 402128
rect 505434 402094 505490 402128
rect 505524 402094 505580 402128
rect 505614 402094 505668 402128
rect 504988 402038 505668 402094
rect 504988 402004 505040 402038
rect 505074 402004 505130 402038
rect 505164 402004 505220 402038
rect 505254 402004 505310 402038
rect 505344 402004 505400 402038
rect 505434 402004 505490 402038
rect 505524 402004 505580 402038
rect 505614 402004 505668 402038
rect 504988 401952 505668 402004
rect 497103 399877 498393 399889
rect 497103 399843 497119 399877
rect 497153 399843 497187 399877
rect 497221 399843 497255 399877
rect 497289 399843 497323 399877
rect 497357 399843 497391 399877
rect 497425 399843 497459 399877
rect 497493 399843 497527 399877
rect 497561 399843 497595 399877
rect 497629 399843 497663 399877
rect 497697 399843 497731 399877
rect 497765 399843 497799 399877
rect 497833 399843 497867 399877
rect 497901 399843 497935 399877
rect 497969 399843 498003 399877
rect 498037 399843 498071 399877
rect 498105 399843 498139 399877
rect 498173 399843 498207 399877
rect 498241 399843 498275 399877
rect 498309 399843 498343 399877
rect 498377 399843 498393 399877
rect 497103 399831 498393 399843
rect 497103 399419 498393 399431
rect 497103 399385 497119 399419
rect 497153 399385 497187 399419
rect 497221 399385 497255 399419
rect 497289 399385 497323 399419
rect 497357 399385 497391 399419
rect 497425 399385 497459 399419
rect 497493 399385 497527 399419
rect 497561 399385 497595 399419
rect 497629 399385 497663 399419
rect 497697 399385 497731 399419
rect 497765 399385 497799 399419
rect 497833 399385 497867 399419
rect 497901 399385 497935 399419
rect 497969 399385 498003 399419
rect 498037 399385 498071 399419
rect 498105 399385 498139 399419
rect 498173 399385 498207 399419
rect 498241 399385 498275 399419
rect 498309 399385 498343 399419
rect 498377 399385 498393 399419
rect 497103 399373 498393 399385
rect 497103 398961 498393 398973
rect 497103 398927 497119 398961
rect 497153 398927 497187 398961
rect 497221 398927 497255 398961
rect 497289 398927 497323 398961
rect 497357 398927 497391 398961
rect 497425 398927 497459 398961
rect 497493 398927 497527 398961
rect 497561 398927 497595 398961
rect 497629 398927 497663 398961
rect 497697 398927 497731 398961
rect 497765 398927 497799 398961
rect 497833 398927 497867 398961
rect 497901 398927 497935 398961
rect 497969 398927 498003 398961
rect 498037 398927 498071 398961
rect 498105 398927 498139 398961
rect 498173 398927 498207 398961
rect 498241 398927 498275 398961
rect 498309 398927 498343 398961
rect 498377 398927 498393 398961
rect 497103 398915 498393 398927
rect 497103 398503 498393 398515
rect 497103 398469 497119 398503
rect 497153 398469 497187 398503
rect 497221 398469 497255 398503
rect 497289 398469 497323 398503
rect 497357 398469 497391 398503
rect 497425 398469 497459 398503
rect 497493 398469 497527 398503
rect 497561 398469 497595 398503
rect 497629 398469 497663 398503
rect 497697 398469 497731 398503
rect 497765 398469 497799 398503
rect 497833 398469 497867 398503
rect 497901 398469 497935 398503
rect 497969 398469 498003 398503
rect 498037 398469 498071 398503
rect 498105 398469 498139 398503
rect 498173 398469 498207 398503
rect 498241 398469 498275 398503
rect 498309 398469 498343 398503
rect 498377 398469 498393 398503
rect 497103 398457 498393 398469
rect 497103 398045 498393 398057
rect 497103 398011 497119 398045
rect 497153 398011 497187 398045
rect 497221 398011 497255 398045
rect 497289 398011 497323 398045
rect 497357 398011 497391 398045
rect 497425 398011 497459 398045
rect 497493 398011 497527 398045
rect 497561 398011 497595 398045
rect 497629 398011 497663 398045
rect 497697 398011 497731 398045
rect 497765 398011 497799 398045
rect 497833 398011 497867 398045
rect 497901 398011 497935 398045
rect 497969 398011 498003 398045
rect 498037 398011 498071 398045
rect 498105 398011 498139 398045
rect 498173 398011 498207 398045
rect 498241 398011 498275 398045
rect 498309 398011 498343 398045
rect 498377 398011 498393 398045
rect 497103 397999 498393 398011
rect 497103 397587 498393 397599
rect 497103 397553 497119 397587
rect 497153 397553 497187 397587
rect 497221 397553 497255 397587
rect 497289 397553 497323 397587
rect 497357 397553 497391 397587
rect 497425 397553 497459 397587
rect 497493 397553 497527 397587
rect 497561 397553 497595 397587
rect 497629 397553 497663 397587
rect 497697 397553 497731 397587
rect 497765 397553 497799 397587
rect 497833 397553 497867 397587
rect 497901 397553 497935 397587
rect 497969 397553 498003 397587
rect 498037 397553 498071 397587
rect 498105 397553 498139 397587
rect 498173 397553 498207 397587
rect 498241 397553 498275 397587
rect 498309 397553 498343 397587
rect 498377 397553 498393 397587
rect 497103 397541 498393 397553
rect 497103 397129 498393 397141
rect 497103 397095 497119 397129
rect 497153 397095 497187 397129
rect 497221 397095 497255 397129
rect 497289 397095 497323 397129
rect 497357 397095 497391 397129
rect 497425 397095 497459 397129
rect 497493 397095 497527 397129
rect 497561 397095 497595 397129
rect 497629 397095 497663 397129
rect 497697 397095 497731 397129
rect 497765 397095 497799 397129
rect 497833 397095 497867 397129
rect 497901 397095 497935 397129
rect 497969 397095 498003 397129
rect 498037 397095 498071 397129
rect 498105 397095 498139 397129
rect 498173 397095 498207 397129
rect 498241 397095 498275 397129
rect 498309 397095 498343 397129
rect 498377 397095 498393 397129
rect 497103 397083 498393 397095
rect 497103 396671 498393 396683
rect 497103 396637 497119 396671
rect 497153 396637 497187 396671
rect 497221 396637 497255 396671
rect 497289 396637 497323 396671
rect 497357 396637 497391 396671
rect 497425 396637 497459 396671
rect 497493 396637 497527 396671
rect 497561 396637 497595 396671
rect 497629 396637 497663 396671
rect 497697 396637 497731 396671
rect 497765 396637 497799 396671
rect 497833 396637 497867 396671
rect 497901 396637 497935 396671
rect 497969 396637 498003 396671
rect 498037 396637 498071 396671
rect 498105 396637 498139 396671
rect 498173 396637 498207 396671
rect 498241 396637 498275 396671
rect 498309 396637 498343 396671
rect 498377 396637 498393 396671
rect 497103 396625 498393 396637
rect 497103 396213 498393 396225
rect 497103 396179 497119 396213
rect 497153 396179 497187 396213
rect 497221 396179 497255 396213
rect 497289 396179 497323 396213
rect 497357 396179 497391 396213
rect 497425 396179 497459 396213
rect 497493 396179 497527 396213
rect 497561 396179 497595 396213
rect 497629 396179 497663 396213
rect 497697 396179 497731 396213
rect 497765 396179 497799 396213
rect 497833 396179 497867 396213
rect 497901 396179 497935 396213
rect 497969 396179 498003 396213
rect 498037 396179 498071 396213
rect 498105 396179 498139 396213
rect 498173 396179 498207 396213
rect 498241 396179 498275 396213
rect 498309 396179 498343 396213
rect 498377 396179 498393 396213
rect 497103 396167 498393 396179
rect 497103 395755 498393 395767
rect 497103 395721 497119 395755
rect 497153 395721 497187 395755
rect 497221 395721 497255 395755
rect 497289 395721 497323 395755
rect 497357 395721 497391 395755
rect 497425 395721 497459 395755
rect 497493 395721 497527 395755
rect 497561 395721 497595 395755
rect 497629 395721 497663 395755
rect 497697 395721 497731 395755
rect 497765 395721 497799 395755
rect 497833 395721 497867 395755
rect 497901 395721 497935 395755
rect 497969 395721 498003 395755
rect 498037 395721 498071 395755
rect 498105 395721 498139 395755
rect 498173 395721 498207 395755
rect 498241 395721 498275 395755
rect 498309 395721 498343 395755
rect 498377 395721 498393 395755
rect 497103 395709 498393 395721
rect 497103 395297 498393 395309
rect 497103 395263 497119 395297
rect 497153 395263 497187 395297
rect 497221 395263 497255 395297
rect 497289 395263 497323 395297
rect 497357 395263 497391 395297
rect 497425 395263 497459 395297
rect 497493 395263 497527 395297
rect 497561 395263 497595 395297
rect 497629 395263 497663 395297
rect 497697 395263 497731 395297
rect 497765 395263 497799 395297
rect 497833 395263 497867 395297
rect 497901 395263 497935 395297
rect 497969 395263 498003 395297
rect 498037 395263 498071 395297
rect 498105 395263 498139 395297
rect 498173 395263 498207 395297
rect 498241 395263 498275 395297
rect 498309 395263 498343 395297
rect 498377 395263 498393 395297
rect 497103 395251 498393 395263
rect 497103 394839 498393 394851
rect 497103 394805 497119 394839
rect 497153 394805 497187 394839
rect 497221 394805 497255 394839
rect 497289 394805 497323 394839
rect 497357 394805 497391 394839
rect 497425 394805 497459 394839
rect 497493 394805 497527 394839
rect 497561 394805 497595 394839
rect 497629 394805 497663 394839
rect 497697 394805 497731 394839
rect 497765 394805 497799 394839
rect 497833 394805 497867 394839
rect 497901 394805 497935 394839
rect 497969 394805 498003 394839
rect 498037 394805 498071 394839
rect 498105 394805 498139 394839
rect 498173 394805 498207 394839
rect 498241 394805 498275 394839
rect 498309 394805 498343 394839
rect 498377 394805 498393 394839
rect 497103 394793 498393 394805
rect 497103 394381 498393 394393
rect 497103 394347 497119 394381
rect 497153 394347 497187 394381
rect 497221 394347 497255 394381
rect 497289 394347 497323 394381
rect 497357 394347 497391 394381
rect 497425 394347 497459 394381
rect 497493 394347 497527 394381
rect 497561 394347 497595 394381
rect 497629 394347 497663 394381
rect 497697 394347 497731 394381
rect 497765 394347 497799 394381
rect 497833 394347 497867 394381
rect 497901 394347 497935 394381
rect 497969 394347 498003 394381
rect 498037 394347 498071 394381
rect 498105 394347 498139 394381
rect 498173 394347 498207 394381
rect 498241 394347 498275 394381
rect 498309 394347 498343 394381
rect 498377 394347 498393 394381
rect 497103 394335 498393 394347
rect 497103 393923 498393 393935
rect 497103 393889 497119 393923
rect 497153 393889 497187 393923
rect 497221 393889 497255 393923
rect 497289 393889 497323 393923
rect 497357 393889 497391 393923
rect 497425 393889 497459 393923
rect 497493 393889 497527 393923
rect 497561 393889 497595 393923
rect 497629 393889 497663 393923
rect 497697 393889 497731 393923
rect 497765 393889 497799 393923
rect 497833 393889 497867 393923
rect 497901 393889 497935 393923
rect 497969 393889 498003 393923
rect 498037 393889 498071 393923
rect 498105 393889 498139 393923
rect 498173 393889 498207 393923
rect 498241 393889 498275 393923
rect 498309 393889 498343 393923
rect 498377 393889 498393 393923
rect 497103 393877 498393 393889
rect 497103 393465 498393 393477
rect 497103 393431 497119 393465
rect 497153 393431 497187 393465
rect 497221 393431 497255 393465
rect 497289 393431 497323 393465
rect 497357 393431 497391 393465
rect 497425 393431 497459 393465
rect 497493 393431 497527 393465
rect 497561 393431 497595 393465
rect 497629 393431 497663 393465
rect 497697 393431 497731 393465
rect 497765 393431 497799 393465
rect 497833 393431 497867 393465
rect 497901 393431 497935 393465
rect 497969 393431 498003 393465
rect 498037 393431 498071 393465
rect 498105 393431 498139 393465
rect 498173 393431 498207 393465
rect 498241 393431 498275 393465
rect 498309 393431 498343 393465
rect 498377 393431 498393 393465
rect 497103 393419 498393 393431
rect 497103 393007 498393 393019
rect 497103 392973 497119 393007
rect 497153 392973 497187 393007
rect 497221 392973 497255 393007
rect 497289 392973 497323 393007
rect 497357 392973 497391 393007
rect 497425 392973 497459 393007
rect 497493 392973 497527 393007
rect 497561 392973 497595 393007
rect 497629 392973 497663 393007
rect 497697 392973 497731 393007
rect 497765 392973 497799 393007
rect 497833 392973 497867 393007
rect 497901 392973 497935 393007
rect 497969 392973 498003 393007
rect 498037 392973 498071 393007
rect 498105 392973 498139 393007
rect 498173 392973 498207 393007
rect 498241 392973 498275 393007
rect 498309 392973 498343 393007
rect 498377 392973 498393 393007
rect 497103 392961 498393 392973
rect 497103 392549 498393 392561
rect 497103 392515 497119 392549
rect 497153 392515 497187 392549
rect 497221 392515 497255 392549
rect 497289 392515 497323 392549
rect 497357 392515 497391 392549
rect 497425 392515 497459 392549
rect 497493 392515 497527 392549
rect 497561 392515 497595 392549
rect 497629 392515 497663 392549
rect 497697 392515 497731 392549
rect 497765 392515 497799 392549
rect 497833 392515 497867 392549
rect 497901 392515 497935 392549
rect 497969 392515 498003 392549
rect 498037 392515 498071 392549
rect 498105 392515 498139 392549
rect 498173 392515 498207 392549
rect 498241 392515 498275 392549
rect 498309 392515 498343 392549
rect 498377 392515 498393 392549
rect 497103 392503 498393 392515
rect 500863 392233 502153 392245
rect 500863 392199 500879 392233
rect 500913 392199 500947 392233
rect 500981 392199 501015 392233
rect 501049 392199 501083 392233
rect 501117 392199 501151 392233
rect 501185 392199 501219 392233
rect 501253 392199 501287 392233
rect 501321 392199 501355 392233
rect 501389 392199 501423 392233
rect 501457 392199 501491 392233
rect 501525 392199 501559 392233
rect 501593 392199 501627 392233
rect 501661 392199 501695 392233
rect 501729 392199 501763 392233
rect 501797 392199 501831 392233
rect 501865 392199 501899 392233
rect 501933 392199 501967 392233
rect 502001 392199 502035 392233
rect 502069 392199 502103 392233
rect 502137 392199 502153 392233
rect 500863 392187 502153 392199
rect 497103 392091 498393 392103
rect 497103 392057 497119 392091
rect 497153 392057 497187 392091
rect 497221 392057 497255 392091
rect 497289 392057 497323 392091
rect 497357 392057 497391 392091
rect 497425 392057 497459 392091
rect 497493 392057 497527 392091
rect 497561 392057 497595 392091
rect 497629 392057 497663 392091
rect 497697 392057 497731 392091
rect 497765 392057 497799 392091
rect 497833 392057 497867 392091
rect 497901 392057 497935 392091
rect 497969 392057 498003 392091
rect 498037 392057 498071 392091
rect 498105 392057 498139 392091
rect 498173 392057 498207 392091
rect 498241 392057 498275 392091
rect 498309 392057 498343 392091
rect 498377 392057 498393 392091
rect 497103 392045 498393 392057
rect 500863 391775 502153 391787
rect 500863 391741 500879 391775
rect 500913 391741 500947 391775
rect 500981 391741 501015 391775
rect 501049 391741 501083 391775
rect 501117 391741 501151 391775
rect 501185 391741 501219 391775
rect 501253 391741 501287 391775
rect 501321 391741 501355 391775
rect 501389 391741 501423 391775
rect 501457 391741 501491 391775
rect 501525 391741 501559 391775
rect 501593 391741 501627 391775
rect 501661 391741 501695 391775
rect 501729 391741 501763 391775
rect 501797 391741 501831 391775
rect 501865 391741 501899 391775
rect 501933 391741 501967 391775
rect 502001 391741 502035 391775
rect 502069 391741 502103 391775
rect 502137 391741 502153 391775
rect 500863 391729 502153 391741
rect 497103 391633 498393 391645
rect 497103 391599 497119 391633
rect 497153 391599 497187 391633
rect 497221 391599 497255 391633
rect 497289 391599 497323 391633
rect 497357 391599 497391 391633
rect 497425 391599 497459 391633
rect 497493 391599 497527 391633
rect 497561 391599 497595 391633
rect 497629 391599 497663 391633
rect 497697 391599 497731 391633
rect 497765 391599 497799 391633
rect 497833 391599 497867 391633
rect 497901 391599 497935 391633
rect 497969 391599 498003 391633
rect 498037 391599 498071 391633
rect 498105 391599 498139 391633
rect 498173 391599 498207 391633
rect 498241 391599 498275 391633
rect 498309 391599 498343 391633
rect 498377 391599 498393 391633
rect 497103 391587 498393 391599
rect 497103 391175 498393 391187
rect 497103 391141 497119 391175
rect 497153 391141 497187 391175
rect 497221 391141 497255 391175
rect 497289 391141 497323 391175
rect 497357 391141 497391 391175
rect 497425 391141 497459 391175
rect 497493 391141 497527 391175
rect 497561 391141 497595 391175
rect 497629 391141 497663 391175
rect 497697 391141 497731 391175
rect 497765 391141 497799 391175
rect 497833 391141 497867 391175
rect 497901 391141 497935 391175
rect 497969 391141 498003 391175
rect 498037 391141 498071 391175
rect 498105 391141 498139 391175
rect 498173 391141 498207 391175
rect 498241 391141 498275 391175
rect 498309 391141 498343 391175
rect 498377 391141 498393 391175
rect 497103 391129 498393 391141
rect 500863 391317 502153 391329
rect 500863 391283 500879 391317
rect 500913 391283 500947 391317
rect 500981 391283 501015 391317
rect 501049 391283 501083 391317
rect 501117 391283 501151 391317
rect 501185 391283 501219 391317
rect 501253 391283 501287 391317
rect 501321 391283 501355 391317
rect 501389 391283 501423 391317
rect 501457 391283 501491 391317
rect 501525 391283 501559 391317
rect 501593 391283 501627 391317
rect 501661 391283 501695 391317
rect 501729 391283 501763 391317
rect 501797 391283 501831 391317
rect 501865 391283 501899 391317
rect 501933 391283 501967 391317
rect 502001 391283 502035 391317
rect 502069 391283 502103 391317
rect 502137 391283 502153 391317
rect 500863 391271 502153 391283
rect 497103 390717 498393 390729
rect 497103 390683 497119 390717
rect 497153 390683 497187 390717
rect 497221 390683 497255 390717
rect 497289 390683 497323 390717
rect 497357 390683 497391 390717
rect 497425 390683 497459 390717
rect 497493 390683 497527 390717
rect 497561 390683 497595 390717
rect 497629 390683 497663 390717
rect 497697 390683 497731 390717
rect 497765 390683 497799 390717
rect 497833 390683 497867 390717
rect 497901 390683 497935 390717
rect 497969 390683 498003 390717
rect 498037 390683 498071 390717
rect 498105 390683 498139 390717
rect 498173 390683 498207 390717
rect 498241 390683 498275 390717
rect 498309 390683 498343 390717
rect 498377 390683 498393 390717
rect 497103 390671 498393 390683
rect 500863 390859 502153 390871
rect 500863 390825 500879 390859
rect 500913 390825 500947 390859
rect 500981 390825 501015 390859
rect 501049 390825 501083 390859
rect 501117 390825 501151 390859
rect 501185 390825 501219 390859
rect 501253 390825 501287 390859
rect 501321 390825 501355 390859
rect 501389 390825 501423 390859
rect 501457 390825 501491 390859
rect 501525 390825 501559 390859
rect 501593 390825 501627 390859
rect 501661 390825 501695 390859
rect 501729 390825 501763 390859
rect 501797 390825 501831 390859
rect 501865 390825 501899 390859
rect 501933 390825 501967 390859
rect 502001 390825 502035 390859
rect 502069 390825 502103 390859
rect 502137 390825 502153 390859
rect 500863 390813 502153 390825
rect 497103 390259 498393 390271
rect 497103 390225 497119 390259
rect 497153 390225 497187 390259
rect 497221 390225 497255 390259
rect 497289 390225 497323 390259
rect 497357 390225 497391 390259
rect 497425 390225 497459 390259
rect 497493 390225 497527 390259
rect 497561 390225 497595 390259
rect 497629 390225 497663 390259
rect 497697 390225 497731 390259
rect 497765 390225 497799 390259
rect 497833 390225 497867 390259
rect 497901 390225 497935 390259
rect 497969 390225 498003 390259
rect 498037 390225 498071 390259
rect 498105 390225 498139 390259
rect 498173 390225 498207 390259
rect 498241 390225 498275 390259
rect 498309 390225 498343 390259
rect 498377 390225 498393 390259
rect 497103 390213 498393 390225
rect 493343 390077 494633 390089
rect 493343 390043 493359 390077
rect 493393 390043 493427 390077
rect 493461 390043 493495 390077
rect 493529 390043 493563 390077
rect 493597 390043 493631 390077
rect 493665 390043 493699 390077
rect 493733 390043 493767 390077
rect 493801 390043 493835 390077
rect 493869 390043 493903 390077
rect 493937 390043 493971 390077
rect 494005 390043 494039 390077
rect 494073 390043 494107 390077
rect 494141 390043 494175 390077
rect 494209 390043 494243 390077
rect 494277 390043 494311 390077
rect 494345 390043 494379 390077
rect 494413 390043 494447 390077
rect 494481 390043 494515 390077
rect 494549 390043 494583 390077
rect 494617 390043 494633 390077
rect 493343 390031 494633 390043
rect 493343 389619 494633 389631
rect 493343 389585 493359 389619
rect 493393 389585 493427 389619
rect 493461 389585 493495 389619
rect 493529 389585 493563 389619
rect 493597 389585 493631 389619
rect 493665 389585 493699 389619
rect 493733 389585 493767 389619
rect 493801 389585 493835 389619
rect 493869 389585 493903 389619
rect 493937 389585 493971 389619
rect 494005 389585 494039 389619
rect 494073 389585 494107 389619
rect 494141 389585 494175 389619
rect 494209 389585 494243 389619
rect 494277 389585 494311 389619
rect 494345 389585 494379 389619
rect 494413 389585 494447 389619
rect 494481 389585 494515 389619
rect 494549 389585 494583 389619
rect 494617 389585 494633 389619
rect 493343 389573 494633 389585
rect 500863 390401 502153 390413
rect 500863 390367 500879 390401
rect 500913 390367 500947 390401
rect 500981 390367 501015 390401
rect 501049 390367 501083 390401
rect 501117 390367 501151 390401
rect 501185 390367 501219 390401
rect 501253 390367 501287 390401
rect 501321 390367 501355 390401
rect 501389 390367 501423 390401
rect 501457 390367 501491 390401
rect 501525 390367 501559 390401
rect 501593 390367 501627 390401
rect 501661 390367 501695 390401
rect 501729 390367 501763 390401
rect 501797 390367 501831 390401
rect 501865 390367 501899 390401
rect 501933 390367 501967 390401
rect 502001 390367 502035 390401
rect 502069 390367 502103 390401
rect 502137 390367 502153 390401
rect 500863 390355 502153 390367
rect 497103 389801 498393 389813
rect 497103 389767 497119 389801
rect 497153 389767 497187 389801
rect 497221 389767 497255 389801
rect 497289 389767 497323 389801
rect 497357 389767 497391 389801
rect 497425 389767 497459 389801
rect 497493 389767 497527 389801
rect 497561 389767 497595 389801
rect 497629 389767 497663 389801
rect 497697 389767 497731 389801
rect 497765 389767 497799 389801
rect 497833 389767 497867 389801
rect 497901 389767 497935 389801
rect 497969 389767 498003 389801
rect 498037 389767 498071 389801
rect 498105 389767 498139 389801
rect 498173 389767 498207 389801
rect 498241 389767 498275 389801
rect 498309 389767 498343 389801
rect 498377 389767 498393 389801
rect 497103 389755 498393 389767
rect 500863 389943 502153 389955
rect 500863 389909 500879 389943
rect 500913 389909 500947 389943
rect 500981 389909 501015 389943
rect 501049 389909 501083 389943
rect 501117 389909 501151 389943
rect 501185 389909 501219 389943
rect 501253 389909 501287 389943
rect 501321 389909 501355 389943
rect 501389 389909 501423 389943
rect 501457 389909 501491 389943
rect 501525 389909 501559 389943
rect 501593 389909 501627 389943
rect 501661 389909 501695 389943
rect 501729 389909 501763 389943
rect 501797 389909 501831 389943
rect 501865 389909 501899 389943
rect 501933 389909 501967 389943
rect 502001 389909 502035 389943
rect 502069 389909 502103 389943
rect 502137 389909 502153 389943
rect 500863 389897 502153 389909
rect 493343 389161 494633 389173
rect 493343 389127 493359 389161
rect 493393 389127 493427 389161
rect 493461 389127 493495 389161
rect 493529 389127 493563 389161
rect 493597 389127 493631 389161
rect 493665 389127 493699 389161
rect 493733 389127 493767 389161
rect 493801 389127 493835 389161
rect 493869 389127 493903 389161
rect 493937 389127 493971 389161
rect 494005 389127 494039 389161
rect 494073 389127 494107 389161
rect 494141 389127 494175 389161
rect 494209 389127 494243 389161
rect 494277 389127 494311 389161
rect 494345 389127 494379 389161
rect 494413 389127 494447 389161
rect 494481 389127 494515 389161
rect 494549 389127 494583 389161
rect 494617 389127 494633 389161
rect 493343 389115 494633 389127
rect 497103 389343 498393 389355
rect 497103 389309 497119 389343
rect 497153 389309 497187 389343
rect 497221 389309 497255 389343
rect 497289 389309 497323 389343
rect 497357 389309 497391 389343
rect 497425 389309 497459 389343
rect 497493 389309 497527 389343
rect 497561 389309 497595 389343
rect 497629 389309 497663 389343
rect 497697 389309 497731 389343
rect 497765 389309 497799 389343
rect 497833 389309 497867 389343
rect 497901 389309 497935 389343
rect 497969 389309 498003 389343
rect 498037 389309 498071 389343
rect 498105 389309 498139 389343
rect 498173 389309 498207 389343
rect 498241 389309 498275 389343
rect 498309 389309 498343 389343
rect 498377 389309 498393 389343
rect 497103 389297 498393 389309
rect 500863 389485 502153 389497
rect 500863 389451 500879 389485
rect 500913 389451 500947 389485
rect 500981 389451 501015 389485
rect 501049 389451 501083 389485
rect 501117 389451 501151 389485
rect 501185 389451 501219 389485
rect 501253 389451 501287 389485
rect 501321 389451 501355 389485
rect 501389 389451 501423 389485
rect 501457 389451 501491 389485
rect 501525 389451 501559 389485
rect 501593 389451 501627 389485
rect 501661 389451 501695 389485
rect 501729 389451 501763 389485
rect 501797 389451 501831 389485
rect 501865 389451 501899 389485
rect 501933 389451 501967 389485
rect 502001 389451 502035 389485
rect 502069 389451 502103 389485
rect 502137 389451 502153 389485
rect 500863 389439 502153 389451
rect 500863 389027 502153 389039
rect 500863 388993 500879 389027
rect 500913 388993 500947 389027
rect 500981 388993 501015 389027
rect 501049 388993 501083 389027
rect 501117 388993 501151 389027
rect 501185 388993 501219 389027
rect 501253 388993 501287 389027
rect 501321 388993 501355 389027
rect 501389 388993 501423 389027
rect 501457 388993 501491 389027
rect 501525 388993 501559 389027
rect 501593 388993 501627 389027
rect 501661 388993 501695 389027
rect 501729 388993 501763 389027
rect 501797 388993 501831 389027
rect 501865 388993 501899 389027
rect 501933 388993 501967 389027
rect 502001 388993 502035 389027
rect 502069 388993 502103 389027
rect 502137 388993 502153 389027
rect 500863 388981 502153 388993
rect 497103 388885 498393 388897
rect 497103 388851 497119 388885
rect 497153 388851 497187 388885
rect 497221 388851 497255 388885
rect 497289 388851 497323 388885
rect 497357 388851 497391 388885
rect 497425 388851 497459 388885
rect 497493 388851 497527 388885
rect 497561 388851 497595 388885
rect 497629 388851 497663 388885
rect 497697 388851 497731 388885
rect 497765 388851 497799 388885
rect 497833 388851 497867 388885
rect 497901 388851 497935 388885
rect 497969 388851 498003 388885
rect 498037 388851 498071 388885
rect 498105 388851 498139 388885
rect 498173 388851 498207 388885
rect 498241 388851 498275 388885
rect 498309 388851 498343 388885
rect 498377 388851 498393 388885
rect 497103 388839 498393 388851
rect 493343 388703 494633 388715
rect 493343 388669 493359 388703
rect 493393 388669 493427 388703
rect 493461 388669 493495 388703
rect 493529 388669 493563 388703
rect 493597 388669 493631 388703
rect 493665 388669 493699 388703
rect 493733 388669 493767 388703
rect 493801 388669 493835 388703
rect 493869 388669 493903 388703
rect 493937 388669 493971 388703
rect 494005 388669 494039 388703
rect 494073 388669 494107 388703
rect 494141 388669 494175 388703
rect 494209 388669 494243 388703
rect 494277 388669 494311 388703
rect 494345 388669 494379 388703
rect 494413 388669 494447 388703
rect 494481 388669 494515 388703
rect 494549 388669 494583 388703
rect 494617 388669 494633 388703
rect 493343 388657 494633 388669
rect 500863 388569 502153 388581
rect 500863 388535 500879 388569
rect 500913 388535 500947 388569
rect 500981 388535 501015 388569
rect 501049 388535 501083 388569
rect 501117 388535 501151 388569
rect 501185 388535 501219 388569
rect 501253 388535 501287 388569
rect 501321 388535 501355 388569
rect 501389 388535 501423 388569
rect 501457 388535 501491 388569
rect 501525 388535 501559 388569
rect 501593 388535 501627 388569
rect 501661 388535 501695 388569
rect 501729 388535 501763 388569
rect 501797 388535 501831 388569
rect 501865 388535 501899 388569
rect 501933 388535 501967 388569
rect 502001 388535 502035 388569
rect 502069 388535 502103 388569
rect 502137 388535 502153 388569
rect 500863 388523 502153 388535
rect 497103 388427 498393 388439
rect 497103 388393 497119 388427
rect 497153 388393 497187 388427
rect 497221 388393 497255 388427
rect 497289 388393 497323 388427
rect 497357 388393 497391 388427
rect 497425 388393 497459 388427
rect 497493 388393 497527 388427
rect 497561 388393 497595 388427
rect 497629 388393 497663 388427
rect 497697 388393 497731 388427
rect 497765 388393 497799 388427
rect 497833 388393 497867 388427
rect 497901 388393 497935 388427
rect 497969 388393 498003 388427
rect 498037 388393 498071 388427
rect 498105 388393 498139 388427
rect 498173 388393 498207 388427
rect 498241 388393 498275 388427
rect 498309 388393 498343 388427
rect 498377 388393 498393 388427
rect 497103 388381 498393 388393
rect 493343 388245 494633 388257
rect 493343 388211 493359 388245
rect 493393 388211 493427 388245
rect 493461 388211 493495 388245
rect 493529 388211 493563 388245
rect 493597 388211 493631 388245
rect 493665 388211 493699 388245
rect 493733 388211 493767 388245
rect 493801 388211 493835 388245
rect 493869 388211 493903 388245
rect 493937 388211 493971 388245
rect 494005 388211 494039 388245
rect 494073 388211 494107 388245
rect 494141 388211 494175 388245
rect 494209 388211 494243 388245
rect 494277 388211 494311 388245
rect 494345 388211 494379 388245
rect 494413 388211 494447 388245
rect 494481 388211 494515 388245
rect 494549 388211 494583 388245
rect 494617 388211 494633 388245
rect 493343 388199 494633 388211
rect 497103 387969 498393 387981
rect 497103 387935 497119 387969
rect 497153 387935 497187 387969
rect 497221 387935 497255 387969
rect 497289 387935 497323 387969
rect 497357 387935 497391 387969
rect 497425 387935 497459 387969
rect 497493 387935 497527 387969
rect 497561 387935 497595 387969
rect 497629 387935 497663 387969
rect 497697 387935 497731 387969
rect 497765 387935 497799 387969
rect 497833 387935 497867 387969
rect 497901 387935 497935 387969
rect 497969 387935 498003 387969
rect 498037 387935 498071 387969
rect 498105 387935 498139 387969
rect 498173 387935 498207 387969
rect 498241 387935 498275 387969
rect 498309 387935 498343 387969
rect 498377 387935 498393 387969
rect 497103 387923 498393 387935
rect 493343 387787 494633 387799
rect 493343 387753 493359 387787
rect 493393 387753 493427 387787
rect 493461 387753 493495 387787
rect 493529 387753 493563 387787
rect 493597 387753 493631 387787
rect 493665 387753 493699 387787
rect 493733 387753 493767 387787
rect 493801 387753 493835 387787
rect 493869 387753 493903 387787
rect 493937 387753 493971 387787
rect 494005 387753 494039 387787
rect 494073 387753 494107 387787
rect 494141 387753 494175 387787
rect 494209 387753 494243 387787
rect 494277 387753 494311 387787
rect 494345 387753 494379 387787
rect 494413 387753 494447 387787
rect 494481 387753 494515 387787
rect 494549 387753 494583 387787
rect 494617 387753 494633 387787
rect 493343 387741 494633 387753
rect 500863 388111 502153 388123
rect 500863 388077 500879 388111
rect 500913 388077 500947 388111
rect 500981 388077 501015 388111
rect 501049 388077 501083 388111
rect 501117 388077 501151 388111
rect 501185 388077 501219 388111
rect 501253 388077 501287 388111
rect 501321 388077 501355 388111
rect 501389 388077 501423 388111
rect 501457 388077 501491 388111
rect 501525 388077 501559 388111
rect 501593 388077 501627 388111
rect 501661 388077 501695 388111
rect 501729 388077 501763 388111
rect 501797 388077 501831 388111
rect 501865 388077 501899 388111
rect 501933 388077 501967 388111
rect 502001 388077 502035 388111
rect 502069 388077 502103 388111
rect 502137 388077 502153 388111
rect 500863 388065 502153 388077
rect 523423 390077 524713 390089
rect 523423 390043 523439 390077
rect 523473 390043 523507 390077
rect 523541 390043 523575 390077
rect 523609 390043 523643 390077
rect 523677 390043 523711 390077
rect 523745 390043 523779 390077
rect 523813 390043 523847 390077
rect 523881 390043 523915 390077
rect 523949 390043 523983 390077
rect 524017 390043 524051 390077
rect 524085 390043 524119 390077
rect 524153 390043 524187 390077
rect 524221 390043 524255 390077
rect 524289 390043 524323 390077
rect 524357 390043 524391 390077
rect 524425 390043 524459 390077
rect 524493 390043 524527 390077
rect 524561 390043 524595 390077
rect 524629 390043 524663 390077
rect 524697 390043 524713 390077
rect 523423 390031 524713 390043
rect 523423 389619 524713 389631
rect 523423 389585 523439 389619
rect 523473 389585 523507 389619
rect 523541 389585 523575 389619
rect 523609 389585 523643 389619
rect 523677 389585 523711 389619
rect 523745 389585 523779 389619
rect 523813 389585 523847 389619
rect 523881 389585 523915 389619
rect 523949 389585 523983 389619
rect 524017 389585 524051 389619
rect 524085 389585 524119 389619
rect 524153 389585 524187 389619
rect 524221 389585 524255 389619
rect 524289 389585 524323 389619
rect 524357 389585 524391 389619
rect 524425 389585 524459 389619
rect 524493 389585 524527 389619
rect 524561 389585 524595 389619
rect 524629 389585 524663 389619
rect 524697 389585 524713 389619
rect 523423 389573 524713 389585
rect 523423 389161 524713 389173
rect 523423 389127 523439 389161
rect 523473 389127 523507 389161
rect 523541 389127 523575 389161
rect 523609 389127 523643 389161
rect 523677 389127 523711 389161
rect 523745 389127 523779 389161
rect 523813 389127 523847 389161
rect 523881 389127 523915 389161
rect 523949 389127 523983 389161
rect 524017 389127 524051 389161
rect 524085 389127 524119 389161
rect 524153 389127 524187 389161
rect 524221 389127 524255 389161
rect 524289 389127 524323 389161
rect 524357 389127 524391 389161
rect 524425 389127 524459 389161
rect 524493 389127 524527 389161
rect 524561 389127 524595 389161
rect 524629 389127 524663 389161
rect 524697 389127 524713 389161
rect 523423 389115 524713 389127
rect 523423 388703 524713 388715
rect 523423 388669 523439 388703
rect 523473 388669 523507 388703
rect 523541 388669 523575 388703
rect 523609 388669 523643 388703
rect 523677 388669 523711 388703
rect 523745 388669 523779 388703
rect 523813 388669 523847 388703
rect 523881 388669 523915 388703
rect 523949 388669 523983 388703
rect 524017 388669 524051 388703
rect 524085 388669 524119 388703
rect 524153 388669 524187 388703
rect 524221 388669 524255 388703
rect 524289 388669 524323 388703
rect 524357 388669 524391 388703
rect 524425 388669 524459 388703
rect 524493 388669 524527 388703
rect 524561 388669 524595 388703
rect 524629 388669 524663 388703
rect 524697 388669 524713 388703
rect 523423 388657 524713 388669
rect 493343 387329 494633 387341
rect 493343 387295 493359 387329
rect 493393 387295 493427 387329
rect 493461 387295 493495 387329
rect 493529 387295 493563 387329
rect 493597 387295 493631 387329
rect 493665 387295 493699 387329
rect 493733 387295 493767 387329
rect 493801 387295 493835 387329
rect 493869 387295 493903 387329
rect 493937 387295 493971 387329
rect 494005 387295 494039 387329
rect 494073 387295 494107 387329
rect 494141 387295 494175 387329
rect 494209 387295 494243 387329
rect 494277 387295 494311 387329
rect 494345 387295 494379 387329
rect 494413 387295 494447 387329
rect 494481 387295 494515 387329
rect 494549 387295 494583 387329
rect 494617 387295 494633 387329
rect 493343 387283 494633 387295
rect 497103 387511 498393 387523
rect 497103 387477 497119 387511
rect 497153 387477 497187 387511
rect 497221 387477 497255 387511
rect 497289 387477 497323 387511
rect 497357 387477 497391 387511
rect 497425 387477 497459 387511
rect 497493 387477 497527 387511
rect 497561 387477 497595 387511
rect 497629 387477 497663 387511
rect 497697 387477 497731 387511
rect 497765 387477 497799 387511
rect 497833 387477 497867 387511
rect 497901 387477 497935 387511
rect 497969 387477 498003 387511
rect 498037 387477 498071 387511
rect 498105 387477 498139 387511
rect 498173 387477 498207 387511
rect 498241 387477 498275 387511
rect 498309 387477 498343 387511
rect 498377 387477 498393 387511
rect 497103 387465 498393 387477
rect 523423 388245 524713 388257
rect 523423 388211 523439 388245
rect 523473 388211 523507 388245
rect 523541 388211 523575 388245
rect 523609 388211 523643 388245
rect 523677 388211 523711 388245
rect 523745 388211 523779 388245
rect 523813 388211 523847 388245
rect 523881 388211 523915 388245
rect 523949 388211 523983 388245
rect 524017 388211 524051 388245
rect 524085 388211 524119 388245
rect 524153 388211 524187 388245
rect 524221 388211 524255 388245
rect 524289 388211 524323 388245
rect 524357 388211 524391 388245
rect 524425 388211 524459 388245
rect 524493 388211 524527 388245
rect 524561 388211 524595 388245
rect 524629 388211 524663 388245
rect 524697 388211 524713 388245
rect 523423 388199 524713 388211
rect 500863 387653 502153 387665
rect 500863 387619 500879 387653
rect 500913 387619 500947 387653
rect 500981 387619 501015 387653
rect 501049 387619 501083 387653
rect 501117 387619 501151 387653
rect 501185 387619 501219 387653
rect 501253 387619 501287 387653
rect 501321 387619 501355 387653
rect 501389 387619 501423 387653
rect 501457 387619 501491 387653
rect 501525 387619 501559 387653
rect 501593 387619 501627 387653
rect 501661 387619 501695 387653
rect 501729 387619 501763 387653
rect 501797 387619 501831 387653
rect 501865 387619 501899 387653
rect 501933 387619 501967 387653
rect 502001 387619 502035 387653
rect 502069 387619 502103 387653
rect 502137 387619 502153 387653
rect 500863 387607 502153 387619
rect 493343 386871 494633 386883
rect 493343 386837 493359 386871
rect 493393 386837 493427 386871
rect 493461 386837 493495 386871
rect 493529 386837 493563 386871
rect 493597 386837 493631 386871
rect 493665 386837 493699 386871
rect 493733 386837 493767 386871
rect 493801 386837 493835 386871
rect 493869 386837 493903 386871
rect 493937 386837 493971 386871
rect 494005 386837 494039 386871
rect 494073 386837 494107 386871
rect 494141 386837 494175 386871
rect 494209 386837 494243 386871
rect 494277 386837 494311 386871
rect 494345 386837 494379 386871
rect 494413 386837 494447 386871
rect 494481 386837 494515 386871
rect 494549 386837 494583 386871
rect 494617 386837 494633 386871
rect 493343 386825 494633 386837
rect 497103 387053 498393 387065
rect 497103 387019 497119 387053
rect 497153 387019 497187 387053
rect 497221 387019 497255 387053
rect 497289 387019 497323 387053
rect 497357 387019 497391 387053
rect 497425 387019 497459 387053
rect 497493 387019 497527 387053
rect 497561 387019 497595 387053
rect 497629 387019 497663 387053
rect 497697 387019 497731 387053
rect 497765 387019 497799 387053
rect 497833 387019 497867 387053
rect 497901 387019 497935 387053
rect 497969 387019 498003 387053
rect 498037 387019 498071 387053
rect 498105 387019 498139 387053
rect 498173 387019 498207 387053
rect 498241 387019 498275 387053
rect 498309 387019 498343 387053
rect 498377 387019 498393 387053
rect 497103 387007 498393 387019
rect 500863 387195 502153 387207
rect 500863 387161 500879 387195
rect 500913 387161 500947 387195
rect 500981 387161 501015 387195
rect 501049 387161 501083 387195
rect 501117 387161 501151 387195
rect 501185 387161 501219 387195
rect 501253 387161 501287 387195
rect 501321 387161 501355 387195
rect 501389 387161 501423 387195
rect 501457 387161 501491 387195
rect 501525 387161 501559 387195
rect 501593 387161 501627 387195
rect 501661 387161 501695 387195
rect 501729 387161 501763 387195
rect 501797 387161 501831 387195
rect 501865 387161 501899 387195
rect 501933 387161 501967 387195
rect 502001 387161 502035 387195
rect 502069 387161 502103 387195
rect 502137 387161 502153 387195
rect 500863 387149 502153 387161
rect 493343 386413 494633 386425
rect 493343 386379 493359 386413
rect 493393 386379 493427 386413
rect 493461 386379 493495 386413
rect 493529 386379 493563 386413
rect 493597 386379 493631 386413
rect 493665 386379 493699 386413
rect 493733 386379 493767 386413
rect 493801 386379 493835 386413
rect 493869 386379 493903 386413
rect 493937 386379 493971 386413
rect 494005 386379 494039 386413
rect 494073 386379 494107 386413
rect 494141 386379 494175 386413
rect 494209 386379 494243 386413
rect 494277 386379 494311 386413
rect 494345 386379 494379 386413
rect 494413 386379 494447 386413
rect 494481 386379 494515 386413
rect 494549 386379 494583 386413
rect 494617 386379 494633 386413
rect 493343 386367 494633 386379
rect 497103 386595 498393 386607
rect 497103 386561 497119 386595
rect 497153 386561 497187 386595
rect 497221 386561 497255 386595
rect 497289 386561 497323 386595
rect 497357 386561 497391 386595
rect 497425 386561 497459 386595
rect 497493 386561 497527 386595
rect 497561 386561 497595 386595
rect 497629 386561 497663 386595
rect 497697 386561 497731 386595
rect 497765 386561 497799 386595
rect 497833 386561 497867 386595
rect 497901 386561 497935 386595
rect 497969 386561 498003 386595
rect 498037 386561 498071 386595
rect 498105 386561 498139 386595
rect 498173 386561 498207 386595
rect 498241 386561 498275 386595
rect 498309 386561 498343 386595
rect 498377 386561 498393 386595
rect 497103 386549 498393 386561
rect 500863 386737 502153 386749
rect 500863 386703 500879 386737
rect 500913 386703 500947 386737
rect 500981 386703 501015 386737
rect 501049 386703 501083 386737
rect 501117 386703 501151 386737
rect 501185 386703 501219 386737
rect 501253 386703 501287 386737
rect 501321 386703 501355 386737
rect 501389 386703 501423 386737
rect 501457 386703 501491 386737
rect 501525 386703 501559 386737
rect 501593 386703 501627 386737
rect 501661 386703 501695 386737
rect 501729 386703 501763 386737
rect 501797 386703 501831 386737
rect 501865 386703 501899 386737
rect 501933 386703 501967 386737
rect 502001 386703 502035 386737
rect 502069 386703 502103 386737
rect 502137 386703 502153 386737
rect 500863 386691 502153 386703
rect 493343 385955 494633 385967
rect 493343 385921 493359 385955
rect 493393 385921 493427 385955
rect 493461 385921 493495 385955
rect 493529 385921 493563 385955
rect 493597 385921 493631 385955
rect 493665 385921 493699 385955
rect 493733 385921 493767 385955
rect 493801 385921 493835 385955
rect 493869 385921 493903 385955
rect 493937 385921 493971 385955
rect 494005 385921 494039 385955
rect 494073 385921 494107 385955
rect 494141 385921 494175 385955
rect 494209 385921 494243 385955
rect 494277 385921 494311 385955
rect 494345 385921 494379 385955
rect 494413 385921 494447 385955
rect 494481 385921 494515 385955
rect 494549 385921 494583 385955
rect 494617 385921 494633 385955
rect 493343 385909 494633 385921
rect 497103 386137 498393 386149
rect 497103 386103 497119 386137
rect 497153 386103 497187 386137
rect 497221 386103 497255 386137
rect 497289 386103 497323 386137
rect 497357 386103 497391 386137
rect 497425 386103 497459 386137
rect 497493 386103 497527 386137
rect 497561 386103 497595 386137
rect 497629 386103 497663 386137
rect 497697 386103 497731 386137
rect 497765 386103 497799 386137
rect 497833 386103 497867 386137
rect 497901 386103 497935 386137
rect 497969 386103 498003 386137
rect 498037 386103 498071 386137
rect 498105 386103 498139 386137
rect 498173 386103 498207 386137
rect 498241 386103 498275 386137
rect 498309 386103 498343 386137
rect 498377 386103 498393 386137
rect 497103 386091 498393 386103
rect 497103 385679 498393 385691
rect 497103 385645 497119 385679
rect 497153 385645 497187 385679
rect 497221 385645 497255 385679
rect 497289 385645 497323 385679
rect 497357 385645 497391 385679
rect 497425 385645 497459 385679
rect 497493 385645 497527 385679
rect 497561 385645 497595 385679
rect 497629 385645 497663 385679
rect 497697 385645 497731 385679
rect 497765 385645 497799 385679
rect 497833 385645 497867 385679
rect 497901 385645 497935 385679
rect 497969 385645 498003 385679
rect 498037 385645 498071 385679
rect 498105 385645 498139 385679
rect 498173 385645 498207 385679
rect 498241 385645 498275 385679
rect 498309 385645 498343 385679
rect 498377 385645 498393 385679
rect 497103 385633 498393 385645
rect 493343 385497 494633 385509
rect 493343 385463 493359 385497
rect 493393 385463 493427 385497
rect 493461 385463 493495 385497
rect 493529 385463 493563 385497
rect 493597 385463 493631 385497
rect 493665 385463 493699 385497
rect 493733 385463 493767 385497
rect 493801 385463 493835 385497
rect 493869 385463 493903 385497
rect 493937 385463 493971 385497
rect 494005 385463 494039 385497
rect 494073 385463 494107 385497
rect 494141 385463 494175 385497
rect 494209 385463 494243 385497
rect 494277 385463 494311 385497
rect 494345 385463 494379 385497
rect 494413 385463 494447 385497
rect 494481 385463 494515 385497
rect 494549 385463 494583 385497
rect 494617 385463 494633 385497
rect 493343 385451 494633 385463
rect 500863 385569 502153 385581
rect 500863 385535 500879 385569
rect 500913 385535 500947 385569
rect 500981 385535 501015 385569
rect 501049 385535 501083 385569
rect 501117 385535 501151 385569
rect 501185 385535 501219 385569
rect 501253 385535 501287 385569
rect 501321 385535 501355 385569
rect 501389 385535 501423 385569
rect 501457 385535 501491 385569
rect 501525 385535 501559 385569
rect 501593 385535 501627 385569
rect 501661 385535 501695 385569
rect 501729 385535 501763 385569
rect 501797 385535 501831 385569
rect 501865 385535 501899 385569
rect 501933 385535 501967 385569
rect 502001 385535 502035 385569
rect 502069 385535 502103 385569
rect 502137 385535 502153 385569
rect 500863 385523 502153 385535
rect 497103 385221 498393 385233
rect 497103 385187 497119 385221
rect 497153 385187 497187 385221
rect 497221 385187 497255 385221
rect 497289 385187 497323 385221
rect 497357 385187 497391 385221
rect 497425 385187 497459 385221
rect 497493 385187 497527 385221
rect 497561 385187 497595 385221
rect 497629 385187 497663 385221
rect 497697 385187 497731 385221
rect 497765 385187 497799 385221
rect 497833 385187 497867 385221
rect 497901 385187 497935 385221
rect 497969 385187 498003 385221
rect 498037 385187 498071 385221
rect 498105 385187 498139 385221
rect 498173 385187 498207 385221
rect 498241 385187 498275 385221
rect 498309 385187 498343 385221
rect 498377 385187 498393 385221
rect 497103 385175 498393 385187
rect 493343 385039 494633 385051
rect 493343 385005 493359 385039
rect 493393 385005 493427 385039
rect 493461 385005 493495 385039
rect 493529 385005 493563 385039
rect 493597 385005 493631 385039
rect 493665 385005 493699 385039
rect 493733 385005 493767 385039
rect 493801 385005 493835 385039
rect 493869 385005 493903 385039
rect 493937 385005 493971 385039
rect 494005 385005 494039 385039
rect 494073 385005 494107 385039
rect 494141 385005 494175 385039
rect 494209 385005 494243 385039
rect 494277 385005 494311 385039
rect 494345 385005 494379 385039
rect 494413 385005 494447 385039
rect 494481 385005 494515 385039
rect 494549 385005 494583 385039
rect 494617 385005 494633 385039
rect 493343 384993 494633 385005
rect 523423 387787 524713 387799
rect 523423 387753 523439 387787
rect 523473 387753 523507 387787
rect 523541 387753 523575 387787
rect 523609 387753 523643 387787
rect 523677 387753 523711 387787
rect 523745 387753 523779 387787
rect 523813 387753 523847 387787
rect 523881 387753 523915 387787
rect 523949 387753 523983 387787
rect 524017 387753 524051 387787
rect 524085 387753 524119 387787
rect 524153 387753 524187 387787
rect 524221 387753 524255 387787
rect 524289 387753 524323 387787
rect 524357 387753 524391 387787
rect 524425 387753 524459 387787
rect 524493 387753 524527 387787
rect 524561 387753 524595 387787
rect 524629 387753 524663 387787
rect 524697 387753 524713 387787
rect 523423 387741 524713 387753
rect 523423 387329 524713 387341
rect 523423 387295 523439 387329
rect 523473 387295 523507 387329
rect 523541 387295 523575 387329
rect 523609 387295 523643 387329
rect 523677 387295 523711 387329
rect 523745 387295 523779 387329
rect 523813 387295 523847 387329
rect 523881 387295 523915 387329
rect 523949 387295 523983 387329
rect 524017 387295 524051 387329
rect 524085 387295 524119 387329
rect 524153 387295 524187 387329
rect 524221 387295 524255 387329
rect 524289 387295 524323 387329
rect 524357 387295 524391 387329
rect 524425 387295 524459 387329
rect 524493 387295 524527 387329
rect 524561 387295 524595 387329
rect 524629 387295 524663 387329
rect 524697 387295 524713 387329
rect 523423 387283 524713 387295
rect 523423 386871 524713 386883
rect 523423 386837 523439 386871
rect 523473 386837 523507 386871
rect 523541 386837 523575 386871
rect 523609 386837 523643 386871
rect 523677 386837 523711 386871
rect 523745 386837 523779 386871
rect 523813 386837 523847 386871
rect 523881 386837 523915 386871
rect 523949 386837 523983 386871
rect 524017 386837 524051 386871
rect 524085 386837 524119 386871
rect 524153 386837 524187 386871
rect 524221 386837 524255 386871
rect 524289 386837 524323 386871
rect 524357 386837 524391 386871
rect 524425 386837 524459 386871
rect 524493 386837 524527 386871
rect 524561 386837 524595 386871
rect 524629 386837 524663 386871
rect 524697 386837 524713 386871
rect 523423 386825 524713 386837
rect 523423 386413 524713 386425
rect 523423 386379 523439 386413
rect 523473 386379 523507 386413
rect 523541 386379 523575 386413
rect 523609 386379 523643 386413
rect 523677 386379 523711 386413
rect 523745 386379 523779 386413
rect 523813 386379 523847 386413
rect 523881 386379 523915 386413
rect 523949 386379 523983 386413
rect 524017 386379 524051 386413
rect 524085 386379 524119 386413
rect 524153 386379 524187 386413
rect 524221 386379 524255 386413
rect 524289 386379 524323 386413
rect 524357 386379 524391 386413
rect 524425 386379 524459 386413
rect 524493 386379 524527 386413
rect 524561 386379 524595 386413
rect 524629 386379 524663 386413
rect 524697 386379 524713 386413
rect 523423 386367 524713 386379
rect 523423 385955 524713 385967
rect 523423 385921 523439 385955
rect 523473 385921 523507 385955
rect 523541 385921 523575 385955
rect 523609 385921 523643 385955
rect 523677 385921 523711 385955
rect 523745 385921 523779 385955
rect 523813 385921 523847 385955
rect 523881 385921 523915 385955
rect 523949 385921 523983 385955
rect 524017 385921 524051 385955
rect 524085 385921 524119 385955
rect 524153 385921 524187 385955
rect 524221 385921 524255 385955
rect 524289 385921 524323 385955
rect 524357 385921 524391 385955
rect 524425 385921 524459 385955
rect 524493 385921 524527 385955
rect 524561 385921 524595 385955
rect 524629 385921 524663 385955
rect 524697 385921 524713 385955
rect 523423 385909 524713 385921
rect 523423 385497 524713 385509
rect 523423 385463 523439 385497
rect 523473 385463 523507 385497
rect 523541 385463 523575 385497
rect 523609 385463 523643 385497
rect 523677 385463 523711 385497
rect 523745 385463 523779 385497
rect 523813 385463 523847 385497
rect 523881 385463 523915 385497
rect 523949 385463 523983 385497
rect 524017 385463 524051 385497
rect 524085 385463 524119 385497
rect 524153 385463 524187 385497
rect 524221 385463 524255 385497
rect 524289 385463 524323 385497
rect 524357 385463 524391 385497
rect 524425 385463 524459 385497
rect 524493 385463 524527 385497
rect 524561 385463 524595 385497
rect 524629 385463 524663 385497
rect 524697 385463 524713 385497
rect 523423 385451 524713 385463
rect 500863 385111 502153 385123
rect 500863 385077 500879 385111
rect 500913 385077 500947 385111
rect 500981 385077 501015 385111
rect 501049 385077 501083 385111
rect 501117 385077 501151 385111
rect 501185 385077 501219 385111
rect 501253 385077 501287 385111
rect 501321 385077 501355 385111
rect 501389 385077 501423 385111
rect 501457 385077 501491 385111
rect 501525 385077 501559 385111
rect 501593 385077 501627 385111
rect 501661 385077 501695 385111
rect 501729 385077 501763 385111
rect 501797 385077 501831 385111
rect 501865 385077 501899 385111
rect 501933 385077 501967 385111
rect 502001 385077 502035 385111
rect 502069 385077 502103 385111
rect 502137 385077 502153 385111
rect 500863 385065 502153 385077
rect 497103 384763 498393 384775
rect 497103 384729 497119 384763
rect 497153 384729 497187 384763
rect 497221 384729 497255 384763
rect 497289 384729 497323 384763
rect 497357 384729 497391 384763
rect 497425 384729 497459 384763
rect 497493 384729 497527 384763
rect 497561 384729 497595 384763
rect 497629 384729 497663 384763
rect 497697 384729 497731 384763
rect 497765 384729 497799 384763
rect 497833 384729 497867 384763
rect 497901 384729 497935 384763
rect 497969 384729 498003 384763
rect 498037 384729 498071 384763
rect 498105 384729 498139 384763
rect 498173 384729 498207 384763
rect 498241 384729 498275 384763
rect 498309 384729 498343 384763
rect 498377 384729 498393 384763
rect 497103 384717 498393 384729
rect 493343 384581 494633 384593
rect 493343 384547 493359 384581
rect 493393 384547 493427 384581
rect 493461 384547 493495 384581
rect 493529 384547 493563 384581
rect 493597 384547 493631 384581
rect 493665 384547 493699 384581
rect 493733 384547 493767 384581
rect 493801 384547 493835 384581
rect 493869 384547 493903 384581
rect 493937 384547 493971 384581
rect 494005 384547 494039 384581
rect 494073 384547 494107 384581
rect 494141 384547 494175 384581
rect 494209 384547 494243 384581
rect 494277 384547 494311 384581
rect 494345 384547 494379 384581
rect 494413 384547 494447 384581
rect 494481 384547 494515 384581
rect 494549 384547 494583 384581
rect 494617 384547 494633 384581
rect 493343 384535 494633 384547
rect 523423 385039 524713 385051
rect 500863 384653 502153 384665
rect 500863 384619 500879 384653
rect 500913 384619 500947 384653
rect 500981 384619 501015 384653
rect 501049 384619 501083 384653
rect 501117 384619 501151 384653
rect 501185 384619 501219 384653
rect 501253 384619 501287 384653
rect 501321 384619 501355 384653
rect 501389 384619 501423 384653
rect 501457 384619 501491 384653
rect 501525 384619 501559 384653
rect 501593 384619 501627 384653
rect 501661 384619 501695 384653
rect 501729 384619 501763 384653
rect 501797 384619 501831 384653
rect 501865 384619 501899 384653
rect 501933 384619 501967 384653
rect 502001 384619 502035 384653
rect 502069 384619 502103 384653
rect 502137 384619 502153 384653
rect 493343 384123 494633 384135
rect 493343 384089 493359 384123
rect 493393 384089 493427 384123
rect 493461 384089 493495 384123
rect 493529 384089 493563 384123
rect 493597 384089 493631 384123
rect 493665 384089 493699 384123
rect 493733 384089 493767 384123
rect 493801 384089 493835 384123
rect 493869 384089 493903 384123
rect 493937 384089 493971 384123
rect 494005 384089 494039 384123
rect 494073 384089 494107 384123
rect 494141 384089 494175 384123
rect 494209 384089 494243 384123
rect 494277 384089 494311 384123
rect 494345 384089 494379 384123
rect 494413 384089 494447 384123
rect 494481 384089 494515 384123
rect 494549 384089 494583 384123
rect 494617 384089 494633 384123
rect 493343 384077 494633 384089
rect 497103 384305 498393 384317
rect 497103 384271 497119 384305
rect 497153 384271 497187 384305
rect 497221 384271 497255 384305
rect 497289 384271 497323 384305
rect 497357 384271 497391 384305
rect 497425 384271 497459 384305
rect 497493 384271 497527 384305
rect 497561 384271 497595 384305
rect 497629 384271 497663 384305
rect 497697 384271 497731 384305
rect 497765 384271 497799 384305
rect 497833 384271 497867 384305
rect 497901 384271 497935 384305
rect 497969 384271 498003 384305
rect 498037 384271 498071 384305
rect 498105 384271 498139 384305
rect 498173 384271 498207 384305
rect 498241 384271 498275 384305
rect 498309 384271 498343 384305
rect 498377 384271 498393 384305
rect 497103 384259 498393 384271
rect 500863 384607 502153 384619
rect 500863 384195 502153 384207
rect 500863 384161 500879 384195
rect 500913 384161 500947 384195
rect 500981 384161 501015 384195
rect 501049 384161 501083 384195
rect 501117 384161 501151 384195
rect 501185 384161 501219 384195
rect 501253 384161 501287 384195
rect 501321 384161 501355 384195
rect 501389 384161 501423 384195
rect 501457 384161 501491 384195
rect 501525 384161 501559 384195
rect 501593 384161 501627 384195
rect 501661 384161 501695 384195
rect 501729 384161 501763 384195
rect 501797 384161 501831 384195
rect 501865 384161 501899 384195
rect 501933 384161 501967 384195
rect 502001 384161 502035 384195
rect 502069 384161 502103 384195
rect 502137 384161 502153 384195
rect 500863 384149 502153 384161
rect 493343 383665 494633 383677
rect 493343 383631 493359 383665
rect 493393 383631 493427 383665
rect 493461 383631 493495 383665
rect 493529 383631 493563 383665
rect 493597 383631 493631 383665
rect 493665 383631 493699 383665
rect 493733 383631 493767 383665
rect 493801 383631 493835 383665
rect 493869 383631 493903 383665
rect 493937 383631 493971 383665
rect 494005 383631 494039 383665
rect 494073 383631 494107 383665
rect 494141 383631 494175 383665
rect 494209 383631 494243 383665
rect 494277 383631 494311 383665
rect 494345 383631 494379 383665
rect 494413 383631 494447 383665
rect 494481 383631 494515 383665
rect 494549 383631 494583 383665
rect 494617 383631 494633 383665
rect 493343 383619 494633 383631
rect 497103 383847 498393 383859
rect 497103 383813 497119 383847
rect 497153 383813 497187 383847
rect 497221 383813 497255 383847
rect 497289 383813 497323 383847
rect 497357 383813 497391 383847
rect 497425 383813 497459 383847
rect 497493 383813 497527 383847
rect 497561 383813 497595 383847
rect 497629 383813 497663 383847
rect 497697 383813 497731 383847
rect 497765 383813 497799 383847
rect 497833 383813 497867 383847
rect 497901 383813 497935 383847
rect 497969 383813 498003 383847
rect 498037 383813 498071 383847
rect 498105 383813 498139 383847
rect 498173 383813 498207 383847
rect 498241 383813 498275 383847
rect 498309 383813 498343 383847
rect 498377 383813 498393 383847
rect 497103 383801 498393 383813
rect 500863 383737 502153 383749
rect 500863 383703 500879 383737
rect 500913 383703 500947 383737
rect 500981 383703 501015 383737
rect 501049 383703 501083 383737
rect 501117 383703 501151 383737
rect 501185 383703 501219 383737
rect 501253 383703 501287 383737
rect 501321 383703 501355 383737
rect 501389 383703 501423 383737
rect 501457 383703 501491 383737
rect 501525 383703 501559 383737
rect 501593 383703 501627 383737
rect 501661 383703 501695 383737
rect 501729 383703 501763 383737
rect 501797 383703 501831 383737
rect 501865 383703 501899 383737
rect 501933 383703 501967 383737
rect 502001 383703 502035 383737
rect 502069 383703 502103 383737
rect 502137 383703 502153 383737
rect 500863 383691 502153 383703
rect 493343 383207 494633 383219
rect 493343 383173 493359 383207
rect 493393 383173 493427 383207
rect 493461 383173 493495 383207
rect 493529 383173 493563 383207
rect 493597 383173 493631 383207
rect 493665 383173 493699 383207
rect 493733 383173 493767 383207
rect 493801 383173 493835 383207
rect 493869 383173 493903 383207
rect 493937 383173 493971 383207
rect 494005 383173 494039 383207
rect 494073 383173 494107 383207
rect 494141 383173 494175 383207
rect 494209 383173 494243 383207
rect 494277 383173 494311 383207
rect 494345 383173 494379 383207
rect 494413 383173 494447 383207
rect 494481 383173 494515 383207
rect 494549 383173 494583 383207
rect 494617 383173 494633 383207
rect 493343 383161 494633 383173
rect 497103 383389 498393 383401
rect 497103 383355 497119 383389
rect 497153 383355 497187 383389
rect 497221 383355 497255 383389
rect 497289 383355 497323 383389
rect 497357 383355 497391 383389
rect 497425 383355 497459 383389
rect 497493 383355 497527 383389
rect 497561 383355 497595 383389
rect 497629 383355 497663 383389
rect 497697 383355 497731 383389
rect 497765 383355 497799 383389
rect 497833 383355 497867 383389
rect 497901 383355 497935 383389
rect 497969 383355 498003 383389
rect 498037 383355 498071 383389
rect 498105 383355 498139 383389
rect 498173 383355 498207 383389
rect 498241 383355 498275 383389
rect 498309 383355 498343 383389
rect 498377 383355 498393 383389
rect 497103 383343 498393 383355
rect 500863 383279 502153 383291
rect 500863 383245 500879 383279
rect 500913 383245 500947 383279
rect 500981 383245 501015 383279
rect 501049 383245 501083 383279
rect 501117 383245 501151 383279
rect 501185 383245 501219 383279
rect 501253 383245 501287 383279
rect 501321 383245 501355 383279
rect 501389 383245 501423 383279
rect 501457 383245 501491 383279
rect 501525 383245 501559 383279
rect 501593 383245 501627 383279
rect 501661 383245 501695 383279
rect 501729 383245 501763 383279
rect 501797 383245 501831 383279
rect 501865 383245 501899 383279
rect 501933 383245 501967 383279
rect 502001 383245 502035 383279
rect 502069 383245 502103 383279
rect 502137 383245 502153 383279
rect 500863 383233 502153 383245
rect 493343 382749 494633 382761
rect 493343 382715 493359 382749
rect 493393 382715 493427 382749
rect 493461 382715 493495 382749
rect 493529 382715 493563 382749
rect 493597 382715 493631 382749
rect 493665 382715 493699 382749
rect 493733 382715 493767 382749
rect 493801 382715 493835 382749
rect 493869 382715 493903 382749
rect 493937 382715 493971 382749
rect 494005 382715 494039 382749
rect 494073 382715 494107 382749
rect 494141 382715 494175 382749
rect 494209 382715 494243 382749
rect 494277 382715 494311 382749
rect 494345 382715 494379 382749
rect 494413 382715 494447 382749
rect 494481 382715 494515 382749
rect 494549 382715 494583 382749
rect 494617 382715 494633 382749
rect 493343 382703 494633 382715
rect 497103 382931 498393 382943
rect 497103 382897 497119 382931
rect 497153 382897 497187 382931
rect 497221 382897 497255 382931
rect 497289 382897 497323 382931
rect 497357 382897 497391 382931
rect 497425 382897 497459 382931
rect 497493 382897 497527 382931
rect 497561 382897 497595 382931
rect 497629 382897 497663 382931
rect 497697 382897 497731 382931
rect 497765 382897 497799 382931
rect 497833 382897 497867 382931
rect 497901 382897 497935 382931
rect 497969 382897 498003 382931
rect 498037 382897 498071 382931
rect 498105 382897 498139 382931
rect 498173 382897 498207 382931
rect 498241 382897 498275 382931
rect 498309 382897 498343 382931
rect 498377 382897 498393 382931
rect 497103 382885 498393 382897
rect 500863 382821 502153 382833
rect 500863 382787 500879 382821
rect 500913 382787 500947 382821
rect 500981 382787 501015 382821
rect 501049 382787 501083 382821
rect 501117 382787 501151 382821
rect 501185 382787 501219 382821
rect 501253 382787 501287 382821
rect 501321 382787 501355 382821
rect 501389 382787 501423 382821
rect 501457 382787 501491 382821
rect 501525 382787 501559 382821
rect 501593 382787 501627 382821
rect 501661 382787 501695 382821
rect 501729 382787 501763 382821
rect 501797 382787 501831 382821
rect 501865 382787 501899 382821
rect 501933 382787 501967 382821
rect 502001 382787 502035 382821
rect 502069 382787 502103 382821
rect 502137 382787 502153 382821
rect 500863 382775 502153 382787
rect 497103 382473 498393 382485
rect 497103 382439 497119 382473
rect 497153 382439 497187 382473
rect 497221 382439 497255 382473
rect 497289 382439 497323 382473
rect 497357 382439 497391 382473
rect 497425 382439 497459 382473
rect 497493 382439 497527 382473
rect 497561 382439 497595 382473
rect 497629 382439 497663 382473
rect 497697 382439 497731 382473
rect 497765 382439 497799 382473
rect 497833 382439 497867 382473
rect 497901 382439 497935 382473
rect 497969 382439 498003 382473
rect 498037 382439 498071 382473
rect 498105 382439 498139 382473
rect 498173 382439 498207 382473
rect 498241 382439 498275 382473
rect 498309 382439 498343 382473
rect 498377 382439 498393 382473
rect 497103 382427 498393 382439
rect 493343 382291 494633 382303
rect 493343 382257 493359 382291
rect 493393 382257 493427 382291
rect 493461 382257 493495 382291
rect 493529 382257 493563 382291
rect 493597 382257 493631 382291
rect 493665 382257 493699 382291
rect 493733 382257 493767 382291
rect 493801 382257 493835 382291
rect 493869 382257 493903 382291
rect 493937 382257 493971 382291
rect 494005 382257 494039 382291
rect 494073 382257 494107 382291
rect 494141 382257 494175 382291
rect 494209 382257 494243 382291
rect 494277 382257 494311 382291
rect 494345 382257 494379 382291
rect 494413 382257 494447 382291
rect 494481 382257 494515 382291
rect 494549 382257 494583 382291
rect 494617 382257 494633 382291
rect 493343 382245 494633 382257
rect 523423 385005 523439 385039
rect 523473 385005 523507 385039
rect 523541 385005 523575 385039
rect 523609 385005 523643 385039
rect 523677 385005 523711 385039
rect 523745 385005 523779 385039
rect 523813 385005 523847 385039
rect 523881 385005 523915 385039
rect 523949 385005 523983 385039
rect 524017 385005 524051 385039
rect 524085 385005 524119 385039
rect 524153 385005 524187 385039
rect 524221 385005 524255 385039
rect 524289 385005 524323 385039
rect 524357 385005 524391 385039
rect 524425 385005 524459 385039
rect 524493 385005 524527 385039
rect 524561 385005 524595 385039
rect 524629 385005 524663 385039
rect 524697 385005 524713 385039
rect 523423 384993 524713 385005
rect 523423 384581 524713 384593
rect 523423 384547 523439 384581
rect 523473 384547 523507 384581
rect 523541 384547 523575 384581
rect 523609 384547 523643 384581
rect 523677 384547 523711 384581
rect 523745 384547 523779 384581
rect 523813 384547 523847 384581
rect 523881 384547 523915 384581
rect 523949 384547 523983 384581
rect 524017 384547 524051 384581
rect 524085 384547 524119 384581
rect 524153 384547 524187 384581
rect 524221 384547 524255 384581
rect 524289 384547 524323 384581
rect 524357 384547 524391 384581
rect 524425 384547 524459 384581
rect 524493 384547 524527 384581
rect 524561 384547 524595 384581
rect 524629 384547 524663 384581
rect 524697 384547 524713 384581
rect 523423 384535 524713 384547
rect 523423 384123 524713 384135
rect 523423 384089 523439 384123
rect 523473 384089 523507 384123
rect 523541 384089 523575 384123
rect 523609 384089 523643 384123
rect 523677 384089 523711 384123
rect 523745 384089 523779 384123
rect 523813 384089 523847 384123
rect 523881 384089 523915 384123
rect 523949 384089 523983 384123
rect 524017 384089 524051 384123
rect 524085 384089 524119 384123
rect 524153 384089 524187 384123
rect 524221 384089 524255 384123
rect 524289 384089 524323 384123
rect 524357 384089 524391 384123
rect 524425 384089 524459 384123
rect 524493 384089 524527 384123
rect 524561 384089 524595 384123
rect 524629 384089 524663 384123
rect 524697 384089 524713 384123
rect 523423 384077 524713 384089
rect 523423 383665 524713 383677
rect 523423 383631 523439 383665
rect 523473 383631 523507 383665
rect 523541 383631 523575 383665
rect 523609 383631 523643 383665
rect 523677 383631 523711 383665
rect 523745 383631 523779 383665
rect 523813 383631 523847 383665
rect 523881 383631 523915 383665
rect 523949 383631 523983 383665
rect 524017 383631 524051 383665
rect 524085 383631 524119 383665
rect 524153 383631 524187 383665
rect 524221 383631 524255 383665
rect 524289 383631 524323 383665
rect 524357 383631 524391 383665
rect 524425 383631 524459 383665
rect 524493 383631 524527 383665
rect 524561 383631 524595 383665
rect 524629 383631 524663 383665
rect 524697 383631 524713 383665
rect 523423 383619 524713 383631
rect 523423 383207 524713 383219
rect 523423 383173 523439 383207
rect 523473 383173 523507 383207
rect 523541 383173 523575 383207
rect 523609 383173 523643 383207
rect 523677 383173 523711 383207
rect 523745 383173 523779 383207
rect 523813 383173 523847 383207
rect 523881 383173 523915 383207
rect 523949 383173 523983 383207
rect 524017 383173 524051 383207
rect 524085 383173 524119 383207
rect 524153 383173 524187 383207
rect 524221 383173 524255 383207
rect 524289 383173 524323 383207
rect 524357 383173 524391 383207
rect 524425 383173 524459 383207
rect 524493 383173 524527 383207
rect 524561 383173 524595 383207
rect 524629 383173 524663 383207
rect 524697 383173 524713 383207
rect 523423 383161 524713 383173
rect 523423 382749 524713 382761
rect 523423 382715 523439 382749
rect 523473 382715 523507 382749
rect 523541 382715 523575 382749
rect 523609 382715 523643 382749
rect 523677 382715 523711 382749
rect 523745 382715 523779 382749
rect 523813 382715 523847 382749
rect 523881 382715 523915 382749
rect 523949 382715 523983 382749
rect 524017 382715 524051 382749
rect 524085 382715 524119 382749
rect 524153 382715 524187 382749
rect 524221 382715 524255 382749
rect 524289 382715 524323 382749
rect 524357 382715 524391 382749
rect 524425 382715 524459 382749
rect 524493 382715 524527 382749
rect 524561 382715 524595 382749
rect 524629 382715 524663 382749
rect 524697 382715 524713 382749
rect 523423 382703 524713 382715
rect 500863 382363 502153 382375
rect 500863 382329 500879 382363
rect 500913 382329 500947 382363
rect 500981 382329 501015 382363
rect 501049 382329 501083 382363
rect 501117 382329 501151 382363
rect 501185 382329 501219 382363
rect 501253 382329 501287 382363
rect 501321 382329 501355 382363
rect 501389 382329 501423 382363
rect 501457 382329 501491 382363
rect 501525 382329 501559 382363
rect 501593 382329 501627 382363
rect 501661 382329 501695 382363
rect 501729 382329 501763 382363
rect 501797 382329 501831 382363
rect 501865 382329 501899 382363
rect 501933 382329 501967 382363
rect 502001 382329 502035 382363
rect 502069 382329 502103 382363
rect 502137 382329 502153 382363
rect 500863 382317 502153 382329
rect 493343 381833 494633 381845
rect 493343 381799 493359 381833
rect 493393 381799 493427 381833
rect 493461 381799 493495 381833
rect 493529 381799 493563 381833
rect 493597 381799 493631 381833
rect 493665 381799 493699 381833
rect 493733 381799 493767 381833
rect 493801 381799 493835 381833
rect 493869 381799 493903 381833
rect 493937 381799 493971 381833
rect 494005 381799 494039 381833
rect 494073 381799 494107 381833
rect 494141 381799 494175 381833
rect 494209 381799 494243 381833
rect 494277 381799 494311 381833
rect 494345 381799 494379 381833
rect 494413 381799 494447 381833
rect 494481 381799 494515 381833
rect 494549 381799 494583 381833
rect 494617 381799 494633 381833
rect 493343 381787 494633 381799
rect 497103 382015 498393 382027
rect 497103 381981 497119 382015
rect 497153 381981 497187 382015
rect 497221 381981 497255 382015
rect 497289 381981 497323 382015
rect 497357 381981 497391 382015
rect 497425 381981 497459 382015
rect 497493 381981 497527 382015
rect 497561 381981 497595 382015
rect 497629 381981 497663 382015
rect 497697 381981 497731 382015
rect 497765 381981 497799 382015
rect 497833 381981 497867 382015
rect 497901 381981 497935 382015
rect 497969 381981 498003 382015
rect 498037 381981 498071 382015
rect 498105 381981 498139 382015
rect 498173 381981 498207 382015
rect 498241 381981 498275 382015
rect 498309 381981 498343 382015
rect 498377 381981 498393 382015
rect 497103 381969 498393 381981
rect 523423 382291 524713 382303
rect 523423 382257 523439 382291
rect 523473 382257 523507 382291
rect 523541 382257 523575 382291
rect 523609 382257 523643 382291
rect 523677 382257 523711 382291
rect 523745 382257 523779 382291
rect 523813 382257 523847 382291
rect 523881 382257 523915 382291
rect 523949 382257 523983 382291
rect 524017 382257 524051 382291
rect 524085 382257 524119 382291
rect 524153 382257 524187 382291
rect 524221 382257 524255 382291
rect 524289 382257 524323 382291
rect 524357 382257 524391 382291
rect 524425 382257 524459 382291
rect 524493 382257 524527 382291
rect 524561 382257 524595 382291
rect 524629 382257 524663 382291
rect 524697 382257 524713 382291
rect 523423 382245 524713 382257
rect 500863 381905 502153 381917
rect 500863 381871 500879 381905
rect 500913 381871 500947 381905
rect 500981 381871 501015 381905
rect 501049 381871 501083 381905
rect 501117 381871 501151 381905
rect 501185 381871 501219 381905
rect 501253 381871 501287 381905
rect 501321 381871 501355 381905
rect 501389 381871 501423 381905
rect 501457 381871 501491 381905
rect 501525 381871 501559 381905
rect 501593 381871 501627 381905
rect 501661 381871 501695 381905
rect 501729 381871 501763 381905
rect 501797 381871 501831 381905
rect 501865 381871 501899 381905
rect 501933 381871 501967 381905
rect 502001 381871 502035 381905
rect 502069 381871 502103 381905
rect 502137 381871 502153 381905
rect 500863 381859 502153 381871
rect 497103 381557 498393 381569
rect 497103 381523 497119 381557
rect 497153 381523 497187 381557
rect 497221 381523 497255 381557
rect 497289 381523 497323 381557
rect 497357 381523 497391 381557
rect 497425 381523 497459 381557
rect 497493 381523 497527 381557
rect 497561 381523 497595 381557
rect 497629 381523 497663 381557
rect 497697 381523 497731 381557
rect 497765 381523 497799 381557
rect 497833 381523 497867 381557
rect 497901 381523 497935 381557
rect 497969 381523 498003 381557
rect 498037 381523 498071 381557
rect 498105 381523 498139 381557
rect 498173 381523 498207 381557
rect 498241 381523 498275 381557
rect 498309 381523 498343 381557
rect 498377 381523 498393 381557
rect 497103 381511 498393 381523
rect 493343 381375 494633 381387
rect 493343 381341 493359 381375
rect 493393 381341 493427 381375
rect 493461 381341 493495 381375
rect 493529 381341 493563 381375
rect 493597 381341 493631 381375
rect 493665 381341 493699 381375
rect 493733 381341 493767 381375
rect 493801 381341 493835 381375
rect 493869 381341 493903 381375
rect 493937 381341 493971 381375
rect 494005 381341 494039 381375
rect 494073 381341 494107 381375
rect 494141 381341 494175 381375
rect 494209 381341 494243 381375
rect 494277 381341 494311 381375
rect 494345 381341 494379 381375
rect 494413 381341 494447 381375
rect 494481 381341 494515 381375
rect 494549 381341 494583 381375
rect 494617 381341 494633 381375
rect 493343 381329 494633 381341
rect 523423 381833 524713 381845
rect 523423 381799 523439 381833
rect 523473 381799 523507 381833
rect 523541 381799 523575 381833
rect 523609 381799 523643 381833
rect 523677 381799 523711 381833
rect 523745 381799 523779 381833
rect 523813 381799 523847 381833
rect 523881 381799 523915 381833
rect 523949 381799 523983 381833
rect 524017 381799 524051 381833
rect 524085 381799 524119 381833
rect 524153 381799 524187 381833
rect 524221 381799 524255 381833
rect 524289 381799 524323 381833
rect 524357 381799 524391 381833
rect 524425 381799 524459 381833
rect 524493 381799 524527 381833
rect 524561 381799 524595 381833
rect 524629 381799 524663 381833
rect 524697 381799 524713 381833
rect 523423 381787 524713 381799
rect 500863 381447 502153 381459
rect 500863 381413 500879 381447
rect 500913 381413 500947 381447
rect 500981 381413 501015 381447
rect 501049 381413 501083 381447
rect 501117 381413 501151 381447
rect 501185 381413 501219 381447
rect 501253 381413 501287 381447
rect 501321 381413 501355 381447
rect 501389 381413 501423 381447
rect 501457 381413 501491 381447
rect 501525 381413 501559 381447
rect 501593 381413 501627 381447
rect 501661 381413 501695 381447
rect 501729 381413 501763 381447
rect 501797 381413 501831 381447
rect 501865 381413 501899 381447
rect 501933 381413 501967 381447
rect 502001 381413 502035 381447
rect 502069 381413 502103 381447
rect 502137 381413 502153 381447
rect 500863 381401 502153 381413
rect 493343 380917 494633 380929
rect 493343 380883 493359 380917
rect 493393 380883 493427 380917
rect 493461 380883 493495 380917
rect 493529 380883 493563 380917
rect 493597 380883 493631 380917
rect 493665 380883 493699 380917
rect 493733 380883 493767 380917
rect 493801 380883 493835 380917
rect 493869 380883 493903 380917
rect 493937 380883 493971 380917
rect 494005 380883 494039 380917
rect 494073 380883 494107 380917
rect 494141 380883 494175 380917
rect 494209 380883 494243 380917
rect 494277 380883 494311 380917
rect 494345 380883 494379 380917
rect 494413 380883 494447 380917
rect 494481 380883 494515 380917
rect 494549 380883 494583 380917
rect 494617 380883 494633 380917
rect 493343 380871 494633 380883
rect 497103 381099 498393 381111
rect 497103 381065 497119 381099
rect 497153 381065 497187 381099
rect 497221 381065 497255 381099
rect 497289 381065 497323 381099
rect 497357 381065 497391 381099
rect 497425 381065 497459 381099
rect 497493 381065 497527 381099
rect 497561 381065 497595 381099
rect 497629 381065 497663 381099
rect 497697 381065 497731 381099
rect 497765 381065 497799 381099
rect 497833 381065 497867 381099
rect 497901 381065 497935 381099
rect 497969 381065 498003 381099
rect 498037 381065 498071 381099
rect 498105 381065 498139 381099
rect 498173 381065 498207 381099
rect 498241 381065 498275 381099
rect 498309 381065 498343 381099
rect 498377 381065 498393 381099
rect 497103 381053 498393 381065
rect 493343 380459 494633 380471
rect 493343 380425 493359 380459
rect 493393 380425 493427 380459
rect 493461 380425 493495 380459
rect 493529 380425 493563 380459
rect 493597 380425 493631 380459
rect 493665 380425 493699 380459
rect 493733 380425 493767 380459
rect 493801 380425 493835 380459
rect 493869 380425 493903 380459
rect 493937 380425 493971 380459
rect 494005 380425 494039 380459
rect 494073 380425 494107 380459
rect 494141 380425 494175 380459
rect 494209 380425 494243 380459
rect 494277 380425 494311 380459
rect 494345 380425 494379 380459
rect 494413 380425 494447 380459
rect 494481 380425 494515 380459
rect 494549 380425 494583 380459
rect 494617 380425 494633 380459
rect 493343 380413 494633 380425
rect 500863 380989 502153 381001
rect 500863 380955 500879 380989
rect 500913 380955 500947 380989
rect 500981 380955 501015 380989
rect 501049 380955 501083 380989
rect 501117 380955 501151 380989
rect 501185 380955 501219 380989
rect 501253 380955 501287 380989
rect 501321 380955 501355 380989
rect 501389 380955 501423 380989
rect 501457 380955 501491 380989
rect 501525 380955 501559 380989
rect 501593 380955 501627 380989
rect 501661 380955 501695 380989
rect 501729 380955 501763 380989
rect 501797 380955 501831 380989
rect 501865 380955 501899 380989
rect 501933 380955 501967 380989
rect 502001 380955 502035 380989
rect 502069 380955 502103 380989
rect 502137 380955 502153 380989
rect 500863 380943 502153 380955
rect 497103 380641 498393 380653
rect 497103 380607 497119 380641
rect 497153 380607 497187 380641
rect 497221 380607 497255 380641
rect 497289 380607 497323 380641
rect 497357 380607 497391 380641
rect 497425 380607 497459 380641
rect 497493 380607 497527 380641
rect 497561 380607 497595 380641
rect 497629 380607 497663 380641
rect 497697 380607 497731 380641
rect 497765 380607 497799 380641
rect 497833 380607 497867 380641
rect 497901 380607 497935 380641
rect 497969 380607 498003 380641
rect 498037 380607 498071 380641
rect 498105 380607 498139 380641
rect 498173 380607 498207 380641
rect 498241 380607 498275 380641
rect 498309 380607 498343 380641
rect 498377 380607 498393 380641
rect 497103 380595 498393 380607
rect 500863 380531 502153 380543
rect 500863 380497 500879 380531
rect 500913 380497 500947 380531
rect 500981 380497 501015 380531
rect 501049 380497 501083 380531
rect 501117 380497 501151 380531
rect 501185 380497 501219 380531
rect 501253 380497 501287 380531
rect 501321 380497 501355 380531
rect 501389 380497 501423 380531
rect 501457 380497 501491 380531
rect 501525 380497 501559 380531
rect 501593 380497 501627 380531
rect 501661 380497 501695 380531
rect 501729 380497 501763 380531
rect 501797 380497 501831 380531
rect 501865 380497 501899 380531
rect 501933 380497 501967 380531
rect 502001 380497 502035 380531
rect 502069 380497 502103 380531
rect 502137 380497 502153 380531
rect 500863 380485 502153 380497
rect 493343 380001 494633 380013
rect 493343 379967 493359 380001
rect 493393 379967 493427 380001
rect 493461 379967 493495 380001
rect 493529 379967 493563 380001
rect 493597 379967 493631 380001
rect 493665 379967 493699 380001
rect 493733 379967 493767 380001
rect 493801 379967 493835 380001
rect 493869 379967 493903 380001
rect 493937 379967 493971 380001
rect 494005 379967 494039 380001
rect 494073 379967 494107 380001
rect 494141 379967 494175 380001
rect 494209 379967 494243 380001
rect 494277 379967 494311 380001
rect 494345 379967 494379 380001
rect 494413 379967 494447 380001
rect 494481 379967 494515 380001
rect 494549 379967 494583 380001
rect 494617 379967 494633 380001
rect 493343 379955 494633 379967
rect 497103 380183 498393 380195
rect 497103 380149 497119 380183
rect 497153 380149 497187 380183
rect 497221 380149 497255 380183
rect 497289 380149 497323 380183
rect 497357 380149 497391 380183
rect 497425 380149 497459 380183
rect 497493 380149 497527 380183
rect 497561 380149 497595 380183
rect 497629 380149 497663 380183
rect 497697 380149 497731 380183
rect 497765 380149 497799 380183
rect 497833 380149 497867 380183
rect 497901 380149 497935 380183
rect 497969 380149 498003 380183
rect 498037 380149 498071 380183
rect 498105 380149 498139 380183
rect 498173 380149 498207 380183
rect 498241 380149 498275 380183
rect 498309 380149 498343 380183
rect 498377 380149 498393 380183
rect 497103 380137 498393 380149
rect 500863 380073 502153 380085
rect 500863 380039 500879 380073
rect 500913 380039 500947 380073
rect 500981 380039 501015 380073
rect 501049 380039 501083 380073
rect 501117 380039 501151 380073
rect 501185 380039 501219 380073
rect 501253 380039 501287 380073
rect 501321 380039 501355 380073
rect 501389 380039 501423 380073
rect 501457 380039 501491 380073
rect 501525 380039 501559 380073
rect 501593 380039 501627 380073
rect 501661 380039 501695 380073
rect 501729 380039 501763 380073
rect 501797 380039 501831 380073
rect 501865 380039 501899 380073
rect 501933 380039 501967 380073
rect 502001 380039 502035 380073
rect 502069 380039 502103 380073
rect 502137 380039 502153 380073
rect 500863 380027 502153 380039
rect 493343 379543 494633 379555
rect 493343 379509 493359 379543
rect 493393 379509 493427 379543
rect 493461 379509 493495 379543
rect 493529 379509 493563 379543
rect 493597 379509 493631 379543
rect 493665 379509 493699 379543
rect 493733 379509 493767 379543
rect 493801 379509 493835 379543
rect 493869 379509 493903 379543
rect 493937 379509 493971 379543
rect 494005 379509 494039 379543
rect 494073 379509 494107 379543
rect 494141 379509 494175 379543
rect 494209 379509 494243 379543
rect 494277 379509 494311 379543
rect 494345 379509 494379 379543
rect 494413 379509 494447 379543
rect 494481 379509 494515 379543
rect 494549 379509 494583 379543
rect 494617 379509 494633 379543
rect 493343 379497 494633 379509
rect 497103 379725 498393 379737
rect 497103 379691 497119 379725
rect 497153 379691 497187 379725
rect 497221 379691 497255 379725
rect 497289 379691 497323 379725
rect 497357 379691 497391 379725
rect 497425 379691 497459 379725
rect 497493 379691 497527 379725
rect 497561 379691 497595 379725
rect 497629 379691 497663 379725
rect 497697 379691 497731 379725
rect 497765 379691 497799 379725
rect 497833 379691 497867 379725
rect 497901 379691 497935 379725
rect 497969 379691 498003 379725
rect 498037 379691 498071 379725
rect 498105 379691 498139 379725
rect 498173 379691 498207 379725
rect 498241 379691 498275 379725
rect 498309 379691 498343 379725
rect 498377 379691 498393 379725
rect 497103 379679 498393 379691
rect 523423 381375 524713 381387
rect 523423 381341 523439 381375
rect 523473 381341 523507 381375
rect 523541 381341 523575 381375
rect 523609 381341 523643 381375
rect 523677 381341 523711 381375
rect 523745 381341 523779 381375
rect 523813 381341 523847 381375
rect 523881 381341 523915 381375
rect 523949 381341 523983 381375
rect 524017 381341 524051 381375
rect 524085 381341 524119 381375
rect 524153 381341 524187 381375
rect 524221 381341 524255 381375
rect 524289 381341 524323 381375
rect 524357 381341 524391 381375
rect 524425 381341 524459 381375
rect 524493 381341 524527 381375
rect 524561 381341 524595 381375
rect 524629 381341 524663 381375
rect 524697 381341 524713 381375
rect 523423 381329 524713 381341
rect 523423 380917 524713 380929
rect 523423 380883 523439 380917
rect 523473 380883 523507 380917
rect 523541 380883 523575 380917
rect 523609 380883 523643 380917
rect 523677 380883 523711 380917
rect 523745 380883 523779 380917
rect 523813 380883 523847 380917
rect 523881 380883 523915 380917
rect 523949 380883 523983 380917
rect 524017 380883 524051 380917
rect 524085 380883 524119 380917
rect 524153 380883 524187 380917
rect 524221 380883 524255 380917
rect 524289 380883 524323 380917
rect 524357 380883 524391 380917
rect 524425 380883 524459 380917
rect 524493 380883 524527 380917
rect 524561 380883 524595 380917
rect 524629 380883 524663 380917
rect 524697 380883 524713 380917
rect 523423 380871 524713 380883
rect 523423 380459 524713 380471
rect 523423 380425 523439 380459
rect 523473 380425 523507 380459
rect 523541 380425 523575 380459
rect 523609 380425 523643 380459
rect 523677 380425 523711 380459
rect 523745 380425 523779 380459
rect 523813 380425 523847 380459
rect 523881 380425 523915 380459
rect 523949 380425 523983 380459
rect 524017 380425 524051 380459
rect 524085 380425 524119 380459
rect 524153 380425 524187 380459
rect 524221 380425 524255 380459
rect 524289 380425 524323 380459
rect 524357 380425 524391 380459
rect 524425 380425 524459 380459
rect 524493 380425 524527 380459
rect 524561 380425 524595 380459
rect 524629 380425 524663 380459
rect 524697 380425 524713 380459
rect 523423 380413 524713 380425
rect 523423 380001 524713 380013
rect 523423 379967 523439 380001
rect 523473 379967 523507 380001
rect 523541 379967 523575 380001
rect 523609 379967 523643 380001
rect 523677 379967 523711 380001
rect 523745 379967 523779 380001
rect 523813 379967 523847 380001
rect 523881 379967 523915 380001
rect 523949 379967 523983 380001
rect 524017 379967 524051 380001
rect 524085 379967 524119 380001
rect 524153 379967 524187 380001
rect 524221 379967 524255 380001
rect 524289 379967 524323 380001
rect 524357 379967 524391 380001
rect 524425 379967 524459 380001
rect 524493 379967 524527 380001
rect 524561 379967 524595 380001
rect 524629 379967 524663 380001
rect 524697 379967 524713 380001
rect 523423 379955 524713 379967
rect 523423 379543 524713 379555
rect 523423 379509 523439 379543
rect 523473 379509 523507 379543
rect 523541 379509 523575 379543
rect 523609 379509 523643 379543
rect 523677 379509 523711 379543
rect 523745 379509 523779 379543
rect 523813 379509 523847 379543
rect 523881 379509 523915 379543
rect 523949 379509 523983 379543
rect 524017 379509 524051 379543
rect 524085 379509 524119 379543
rect 524153 379509 524187 379543
rect 524221 379509 524255 379543
rect 524289 379509 524323 379543
rect 524357 379509 524391 379543
rect 524425 379509 524459 379543
rect 524493 379509 524527 379543
rect 524561 379509 524595 379543
rect 524629 379509 524663 379543
rect 524697 379509 524713 379543
rect 523423 379497 524713 379509
rect 497103 379267 498393 379279
rect 497103 379233 497119 379267
rect 497153 379233 497187 379267
rect 497221 379233 497255 379267
rect 497289 379233 497323 379267
rect 497357 379233 497391 379267
rect 497425 379233 497459 379267
rect 497493 379233 497527 379267
rect 497561 379233 497595 379267
rect 497629 379233 497663 379267
rect 497697 379233 497731 379267
rect 497765 379233 497799 379267
rect 497833 379233 497867 379267
rect 497901 379233 497935 379267
rect 497969 379233 498003 379267
rect 498037 379233 498071 379267
rect 498105 379233 498139 379267
rect 498173 379233 498207 379267
rect 498241 379233 498275 379267
rect 498309 379233 498343 379267
rect 498377 379233 498393 379267
rect 497103 379221 498393 379233
rect 493343 379085 494633 379097
rect 493343 379051 493359 379085
rect 493393 379051 493427 379085
rect 493461 379051 493495 379085
rect 493529 379051 493563 379085
rect 493597 379051 493631 379085
rect 493665 379051 493699 379085
rect 493733 379051 493767 379085
rect 493801 379051 493835 379085
rect 493869 379051 493903 379085
rect 493937 379051 493971 379085
rect 494005 379051 494039 379085
rect 494073 379051 494107 379085
rect 494141 379051 494175 379085
rect 494209 379051 494243 379085
rect 494277 379051 494311 379085
rect 494345 379051 494379 379085
rect 494413 379051 494447 379085
rect 494481 379051 494515 379085
rect 494549 379051 494583 379085
rect 494617 379051 494633 379085
rect 493343 379039 494633 379051
rect 523423 379085 524713 379097
rect 523423 379051 523439 379085
rect 523473 379051 523507 379085
rect 523541 379051 523575 379085
rect 523609 379051 523643 379085
rect 523677 379051 523711 379085
rect 523745 379051 523779 379085
rect 523813 379051 523847 379085
rect 523881 379051 523915 379085
rect 523949 379051 523983 379085
rect 524017 379051 524051 379085
rect 524085 379051 524119 379085
rect 524153 379051 524187 379085
rect 524221 379051 524255 379085
rect 524289 379051 524323 379085
rect 524357 379051 524391 379085
rect 524425 379051 524459 379085
rect 524493 379051 524527 379085
rect 524561 379051 524595 379085
rect 524629 379051 524663 379085
rect 524697 379051 524713 379085
rect 523423 379039 524713 379051
rect 497103 378809 498393 378821
rect 497103 378775 497119 378809
rect 497153 378775 497187 378809
rect 497221 378775 497255 378809
rect 497289 378775 497323 378809
rect 497357 378775 497391 378809
rect 497425 378775 497459 378809
rect 497493 378775 497527 378809
rect 497561 378775 497595 378809
rect 497629 378775 497663 378809
rect 497697 378775 497731 378809
rect 497765 378775 497799 378809
rect 497833 378775 497867 378809
rect 497901 378775 497935 378809
rect 497969 378775 498003 378809
rect 498037 378775 498071 378809
rect 498105 378775 498139 378809
rect 498173 378775 498207 378809
rect 498241 378775 498275 378809
rect 498309 378775 498343 378809
rect 498377 378775 498393 378809
rect 497103 378763 498393 378775
rect 493343 378627 494633 378639
rect 493343 378593 493359 378627
rect 493393 378593 493427 378627
rect 493461 378593 493495 378627
rect 493529 378593 493563 378627
rect 493597 378593 493631 378627
rect 493665 378593 493699 378627
rect 493733 378593 493767 378627
rect 493801 378593 493835 378627
rect 493869 378593 493903 378627
rect 493937 378593 493971 378627
rect 494005 378593 494039 378627
rect 494073 378593 494107 378627
rect 494141 378593 494175 378627
rect 494209 378593 494243 378627
rect 494277 378593 494311 378627
rect 494345 378593 494379 378627
rect 494413 378593 494447 378627
rect 494481 378593 494515 378627
rect 494549 378593 494583 378627
rect 494617 378593 494633 378627
rect 493343 378581 494633 378593
rect 523423 378627 524713 378639
rect 523423 378593 523439 378627
rect 523473 378593 523507 378627
rect 523541 378593 523575 378627
rect 523609 378593 523643 378627
rect 523677 378593 523711 378627
rect 523745 378593 523779 378627
rect 523813 378593 523847 378627
rect 523881 378593 523915 378627
rect 523949 378593 523983 378627
rect 524017 378593 524051 378627
rect 524085 378593 524119 378627
rect 524153 378593 524187 378627
rect 524221 378593 524255 378627
rect 524289 378593 524323 378627
rect 524357 378593 524391 378627
rect 524425 378593 524459 378627
rect 524493 378593 524527 378627
rect 524561 378593 524595 378627
rect 524629 378593 524663 378627
rect 524697 378593 524713 378627
rect 523423 378581 524713 378593
rect 493343 378169 494633 378181
rect 493343 378135 493359 378169
rect 493393 378135 493427 378169
rect 493461 378135 493495 378169
rect 493529 378135 493563 378169
rect 493597 378135 493631 378169
rect 493665 378135 493699 378169
rect 493733 378135 493767 378169
rect 493801 378135 493835 378169
rect 493869 378135 493903 378169
rect 493937 378135 493971 378169
rect 494005 378135 494039 378169
rect 494073 378135 494107 378169
rect 494141 378135 494175 378169
rect 494209 378135 494243 378169
rect 494277 378135 494311 378169
rect 494345 378135 494379 378169
rect 494413 378135 494447 378169
rect 494481 378135 494515 378169
rect 494549 378135 494583 378169
rect 494617 378135 494633 378169
rect 493343 378123 494633 378135
rect 497103 378351 498393 378363
rect 497103 378317 497119 378351
rect 497153 378317 497187 378351
rect 497221 378317 497255 378351
rect 497289 378317 497323 378351
rect 497357 378317 497391 378351
rect 497425 378317 497459 378351
rect 497493 378317 497527 378351
rect 497561 378317 497595 378351
rect 497629 378317 497663 378351
rect 497697 378317 497731 378351
rect 497765 378317 497799 378351
rect 497833 378317 497867 378351
rect 497901 378317 497935 378351
rect 497969 378317 498003 378351
rect 498037 378317 498071 378351
rect 498105 378317 498139 378351
rect 498173 378317 498207 378351
rect 498241 378317 498275 378351
rect 498309 378317 498343 378351
rect 498377 378317 498393 378351
rect 497103 378305 498393 378317
rect 493343 377711 494633 377723
rect 493343 377677 493359 377711
rect 493393 377677 493427 377711
rect 493461 377677 493495 377711
rect 493529 377677 493563 377711
rect 493597 377677 493631 377711
rect 493665 377677 493699 377711
rect 493733 377677 493767 377711
rect 493801 377677 493835 377711
rect 493869 377677 493903 377711
rect 493937 377677 493971 377711
rect 494005 377677 494039 377711
rect 494073 377677 494107 377711
rect 494141 377677 494175 377711
rect 494209 377677 494243 377711
rect 494277 377677 494311 377711
rect 494345 377677 494379 377711
rect 494413 377677 494447 377711
rect 494481 377677 494515 377711
rect 494549 377677 494583 377711
rect 494617 377677 494633 377711
rect 493343 377665 494633 377677
rect 523423 378169 524713 378181
rect 523423 378135 523439 378169
rect 523473 378135 523507 378169
rect 523541 378135 523575 378169
rect 523609 378135 523643 378169
rect 523677 378135 523711 378169
rect 523745 378135 523779 378169
rect 523813 378135 523847 378169
rect 523881 378135 523915 378169
rect 523949 378135 523983 378169
rect 524017 378135 524051 378169
rect 524085 378135 524119 378169
rect 524153 378135 524187 378169
rect 524221 378135 524255 378169
rect 524289 378135 524323 378169
rect 524357 378135 524391 378169
rect 524425 378135 524459 378169
rect 524493 378135 524527 378169
rect 524561 378135 524595 378169
rect 524629 378135 524663 378169
rect 524697 378135 524713 378169
rect 523423 378123 524713 378135
rect 497103 377893 498393 377905
rect 497103 377859 497119 377893
rect 497153 377859 497187 377893
rect 497221 377859 497255 377893
rect 497289 377859 497323 377893
rect 497357 377859 497391 377893
rect 497425 377859 497459 377893
rect 497493 377859 497527 377893
rect 497561 377859 497595 377893
rect 497629 377859 497663 377893
rect 497697 377859 497731 377893
rect 497765 377859 497799 377893
rect 497833 377859 497867 377893
rect 497901 377859 497935 377893
rect 497969 377859 498003 377893
rect 498037 377859 498071 377893
rect 498105 377859 498139 377893
rect 498173 377859 498207 377893
rect 498241 377859 498275 377893
rect 498309 377859 498343 377893
rect 498377 377859 498393 377893
rect 497103 377847 498393 377859
rect 493343 377253 494633 377265
rect 493343 377219 493359 377253
rect 493393 377219 493427 377253
rect 493461 377219 493495 377253
rect 493529 377219 493563 377253
rect 493597 377219 493631 377253
rect 493665 377219 493699 377253
rect 493733 377219 493767 377253
rect 493801 377219 493835 377253
rect 493869 377219 493903 377253
rect 493937 377219 493971 377253
rect 494005 377219 494039 377253
rect 494073 377219 494107 377253
rect 494141 377219 494175 377253
rect 494209 377219 494243 377253
rect 494277 377219 494311 377253
rect 494345 377219 494379 377253
rect 494413 377219 494447 377253
rect 494481 377219 494515 377253
rect 494549 377219 494583 377253
rect 494617 377219 494633 377253
rect 493343 377207 494633 377219
rect 523423 377711 524713 377723
rect 497103 377435 498393 377447
rect 497103 377401 497119 377435
rect 497153 377401 497187 377435
rect 497221 377401 497255 377435
rect 497289 377401 497323 377435
rect 497357 377401 497391 377435
rect 497425 377401 497459 377435
rect 497493 377401 497527 377435
rect 497561 377401 497595 377435
rect 497629 377401 497663 377435
rect 497697 377401 497731 377435
rect 497765 377401 497799 377435
rect 497833 377401 497867 377435
rect 497901 377401 497935 377435
rect 497969 377401 498003 377435
rect 498037 377401 498071 377435
rect 498105 377401 498139 377435
rect 498173 377401 498207 377435
rect 498241 377401 498275 377435
rect 498309 377401 498343 377435
rect 498377 377401 498393 377435
rect 497103 377389 498393 377401
rect 493343 376795 494633 376807
rect 493343 376761 493359 376795
rect 493393 376761 493427 376795
rect 493461 376761 493495 376795
rect 493529 376761 493563 376795
rect 493597 376761 493631 376795
rect 493665 376761 493699 376795
rect 493733 376761 493767 376795
rect 493801 376761 493835 376795
rect 493869 376761 493903 376795
rect 493937 376761 493971 376795
rect 494005 376761 494039 376795
rect 494073 376761 494107 376795
rect 494141 376761 494175 376795
rect 494209 376761 494243 376795
rect 494277 376761 494311 376795
rect 494345 376761 494379 376795
rect 494413 376761 494447 376795
rect 494481 376761 494515 376795
rect 494549 376761 494583 376795
rect 494617 376761 494633 376795
rect 493343 376749 494633 376761
rect 523423 377677 523439 377711
rect 523473 377677 523507 377711
rect 523541 377677 523575 377711
rect 523609 377677 523643 377711
rect 523677 377677 523711 377711
rect 523745 377677 523779 377711
rect 523813 377677 523847 377711
rect 523881 377677 523915 377711
rect 523949 377677 523983 377711
rect 524017 377677 524051 377711
rect 524085 377677 524119 377711
rect 524153 377677 524187 377711
rect 524221 377677 524255 377711
rect 524289 377677 524323 377711
rect 524357 377677 524391 377711
rect 524425 377677 524459 377711
rect 524493 377677 524527 377711
rect 524561 377677 524595 377711
rect 524629 377677 524663 377711
rect 524697 377677 524713 377711
rect 523423 377665 524713 377677
rect 504623 377435 505913 377447
rect 504623 377401 504639 377435
rect 504673 377401 504707 377435
rect 504741 377401 504775 377435
rect 504809 377401 504843 377435
rect 504877 377401 504911 377435
rect 504945 377401 504979 377435
rect 505013 377401 505047 377435
rect 505081 377401 505115 377435
rect 505149 377401 505183 377435
rect 505217 377401 505251 377435
rect 505285 377401 505319 377435
rect 505353 377401 505387 377435
rect 505421 377401 505455 377435
rect 505489 377401 505523 377435
rect 505557 377401 505591 377435
rect 505625 377401 505659 377435
rect 505693 377401 505727 377435
rect 505761 377401 505795 377435
rect 505829 377401 505863 377435
rect 505897 377401 505913 377435
rect 504623 377389 505913 377401
rect 497103 376977 498393 376989
rect 497103 376943 497119 376977
rect 497153 376943 497187 376977
rect 497221 376943 497255 376977
rect 497289 376943 497323 376977
rect 497357 376943 497391 376977
rect 497425 376943 497459 376977
rect 497493 376943 497527 376977
rect 497561 376943 497595 376977
rect 497629 376943 497663 376977
rect 497697 376943 497731 376977
rect 497765 376943 497799 376977
rect 497833 376943 497867 376977
rect 497901 376943 497935 376977
rect 497969 376943 498003 376977
rect 498037 376943 498071 376977
rect 498105 376943 498139 376977
rect 498173 376943 498207 376977
rect 498241 376943 498275 376977
rect 498309 376943 498343 376977
rect 498377 376943 498393 376977
rect 497103 376931 498393 376943
rect 493343 376337 494633 376349
rect 493343 376303 493359 376337
rect 493393 376303 493427 376337
rect 493461 376303 493495 376337
rect 493529 376303 493563 376337
rect 493597 376303 493631 376337
rect 493665 376303 493699 376337
rect 493733 376303 493767 376337
rect 493801 376303 493835 376337
rect 493869 376303 493903 376337
rect 493937 376303 493971 376337
rect 494005 376303 494039 376337
rect 494073 376303 494107 376337
rect 494141 376303 494175 376337
rect 494209 376303 494243 376337
rect 494277 376303 494311 376337
rect 494345 376303 494379 376337
rect 494413 376303 494447 376337
rect 494481 376303 494515 376337
rect 494549 376303 494583 376337
rect 494617 376303 494633 376337
rect 493343 376291 494633 376303
rect 512143 377435 513433 377447
rect 512143 377401 512159 377435
rect 512193 377401 512227 377435
rect 512261 377401 512295 377435
rect 512329 377401 512363 377435
rect 512397 377401 512431 377435
rect 512465 377401 512499 377435
rect 512533 377401 512567 377435
rect 512601 377401 512635 377435
rect 512669 377401 512703 377435
rect 512737 377401 512771 377435
rect 512805 377401 512839 377435
rect 512873 377401 512907 377435
rect 512941 377401 512975 377435
rect 513009 377401 513043 377435
rect 513077 377401 513111 377435
rect 513145 377401 513179 377435
rect 513213 377401 513247 377435
rect 513281 377401 513315 377435
rect 513349 377401 513383 377435
rect 513417 377401 513433 377435
rect 512143 377389 513433 377401
rect 504623 376977 505913 376989
rect 504623 376943 504639 376977
rect 504673 376943 504707 376977
rect 504741 376943 504775 376977
rect 504809 376943 504843 376977
rect 504877 376943 504911 376977
rect 504945 376943 504979 376977
rect 505013 376943 505047 376977
rect 505081 376943 505115 376977
rect 505149 376943 505183 376977
rect 505217 376943 505251 376977
rect 505285 376943 505319 376977
rect 505353 376943 505387 376977
rect 505421 376943 505455 376977
rect 505489 376943 505523 376977
rect 505557 376943 505591 376977
rect 505625 376943 505659 376977
rect 505693 376943 505727 376977
rect 505761 376943 505795 376977
rect 505829 376943 505863 376977
rect 505897 376943 505913 376977
rect 504623 376931 505913 376943
rect 497103 376519 498393 376531
rect 497103 376485 497119 376519
rect 497153 376485 497187 376519
rect 497221 376485 497255 376519
rect 497289 376485 497323 376519
rect 497357 376485 497391 376519
rect 497425 376485 497459 376519
rect 497493 376485 497527 376519
rect 497561 376485 497595 376519
rect 497629 376485 497663 376519
rect 497697 376485 497731 376519
rect 497765 376485 497799 376519
rect 497833 376485 497867 376519
rect 497901 376485 497935 376519
rect 497969 376485 498003 376519
rect 498037 376485 498071 376519
rect 498105 376485 498139 376519
rect 498173 376485 498207 376519
rect 498241 376485 498275 376519
rect 498309 376485 498343 376519
rect 498377 376485 498393 376519
rect 497103 376473 498393 376485
rect 512143 376977 513433 376989
rect 512143 376943 512159 376977
rect 512193 376943 512227 376977
rect 512261 376943 512295 376977
rect 512329 376943 512363 376977
rect 512397 376943 512431 376977
rect 512465 376943 512499 376977
rect 512533 376943 512567 376977
rect 512601 376943 512635 376977
rect 512669 376943 512703 376977
rect 512737 376943 512771 376977
rect 512805 376943 512839 376977
rect 512873 376943 512907 376977
rect 512941 376943 512975 376977
rect 513009 376943 513043 376977
rect 513077 376943 513111 376977
rect 513145 376943 513179 376977
rect 513213 376943 513247 376977
rect 513281 376943 513315 376977
rect 513349 376943 513383 376977
rect 513417 376943 513433 376977
rect 512143 376931 513433 376943
rect 504623 376519 505913 376531
rect 504623 376485 504639 376519
rect 504673 376485 504707 376519
rect 504741 376485 504775 376519
rect 504809 376485 504843 376519
rect 504877 376485 504911 376519
rect 504945 376485 504979 376519
rect 505013 376485 505047 376519
rect 505081 376485 505115 376519
rect 505149 376485 505183 376519
rect 505217 376485 505251 376519
rect 505285 376485 505319 376519
rect 505353 376485 505387 376519
rect 505421 376485 505455 376519
rect 505489 376485 505523 376519
rect 505557 376485 505591 376519
rect 505625 376485 505659 376519
rect 505693 376485 505727 376519
rect 505761 376485 505795 376519
rect 505829 376485 505863 376519
rect 505897 376485 505913 376519
rect 504623 376473 505913 376485
rect 497103 376061 498393 376073
rect 497103 376027 497119 376061
rect 497153 376027 497187 376061
rect 497221 376027 497255 376061
rect 497289 376027 497323 376061
rect 497357 376027 497391 376061
rect 497425 376027 497459 376061
rect 497493 376027 497527 376061
rect 497561 376027 497595 376061
rect 497629 376027 497663 376061
rect 497697 376027 497731 376061
rect 497765 376027 497799 376061
rect 497833 376027 497867 376061
rect 497901 376027 497935 376061
rect 497969 376027 498003 376061
rect 498037 376027 498071 376061
rect 498105 376027 498139 376061
rect 498173 376027 498207 376061
rect 498241 376027 498275 376061
rect 498309 376027 498343 376061
rect 498377 376027 498393 376061
rect 497103 376015 498393 376027
rect 493343 375879 494633 375891
rect 493343 375845 493359 375879
rect 493393 375845 493427 375879
rect 493461 375845 493495 375879
rect 493529 375845 493563 375879
rect 493597 375845 493631 375879
rect 493665 375845 493699 375879
rect 493733 375845 493767 375879
rect 493801 375845 493835 375879
rect 493869 375845 493903 375879
rect 493937 375845 493971 375879
rect 494005 375845 494039 375879
rect 494073 375845 494107 375879
rect 494141 375845 494175 375879
rect 494209 375845 494243 375879
rect 494277 375845 494311 375879
rect 494345 375845 494379 375879
rect 494413 375845 494447 375879
rect 494481 375845 494515 375879
rect 494549 375845 494583 375879
rect 494617 375845 494633 375879
rect 493343 375833 494633 375845
rect 512143 376519 513433 376531
rect 512143 376485 512159 376519
rect 512193 376485 512227 376519
rect 512261 376485 512295 376519
rect 512329 376485 512363 376519
rect 512397 376485 512431 376519
rect 512465 376485 512499 376519
rect 512533 376485 512567 376519
rect 512601 376485 512635 376519
rect 512669 376485 512703 376519
rect 512737 376485 512771 376519
rect 512805 376485 512839 376519
rect 512873 376485 512907 376519
rect 512941 376485 512975 376519
rect 513009 376485 513043 376519
rect 513077 376485 513111 376519
rect 513145 376485 513179 376519
rect 513213 376485 513247 376519
rect 513281 376485 513315 376519
rect 513349 376485 513383 376519
rect 513417 376485 513433 376519
rect 512143 376473 513433 376485
rect 504623 376061 505913 376073
rect 504623 376027 504639 376061
rect 504673 376027 504707 376061
rect 504741 376027 504775 376061
rect 504809 376027 504843 376061
rect 504877 376027 504911 376061
rect 504945 376027 504979 376061
rect 505013 376027 505047 376061
rect 505081 376027 505115 376061
rect 505149 376027 505183 376061
rect 505217 376027 505251 376061
rect 505285 376027 505319 376061
rect 505353 376027 505387 376061
rect 505421 376027 505455 376061
rect 505489 376027 505523 376061
rect 505557 376027 505591 376061
rect 505625 376027 505659 376061
rect 505693 376027 505727 376061
rect 505761 376027 505795 376061
rect 505829 376027 505863 376061
rect 505897 376027 505913 376061
rect 504623 376015 505913 376027
rect 497103 375603 498393 375615
rect 497103 375569 497119 375603
rect 497153 375569 497187 375603
rect 497221 375569 497255 375603
rect 497289 375569 497323 375603
rect 497357 375569 497391 375603
rect 497425 375569 497459 375603
rect 497493 375569 497527 375603
rect 497561 375569 497595 375603
rect 497629 375569 497663 375603
rect 497697 375569 497731 375603
rect 497765 375569 497799 375603
rect 497833 375569 497867 375603
rect 497901 375569 497935 375603
rect 497969 375569 498003 375603
rect 498037 375569 498071 375603
rect 498105 375569 498139 375603
rect 498173 375569 498207 375603
rect 498241 375569 498275 375603
rect 498309 375569 498343 375603
rect 498377 375569 498393 375603
rect 497103 375557 498393 375569
rect 493343 375421 494633 375433
rect 493343 375387 493359 375421
rect 493393 375387 493427 375421
rect 493461 375387 493495 375421
rect 493529 375387 493563 375421
rect 493597 375387 493631 375421
rect 493665 375387 493699 375421
rect 493733 375387 493767 375421
rect 493801 375387 493835 375421
rect 493869 375387 493903 375421
rect 493937 375387 493971 375421
rect 494005 375387 494039 375421
rect 494073 375387 494107 375421
rect 494141 375387 494175 375421
rect 494209 375387 494243 375421
rect 494277 375387 494311 375421
rect 494345 375387 494379 375421
rect 494413 375387 494447 375421
rect 494481 375387 494515 375421
rect 494549 375387 494583 375421
rect 494617 375387 494633 375421
rect 493343 375375 494633 375387
rect 512143 376061 513433 376073
rect 512143 376027 512159 376061
rect 512193 376027 512227 376061
rect 512261 376027 512295 376061
rect 512329 376027 512363 376061
rect 512397 376027 512431 376061
rect 512465 376027 512499 376061
rect 512533 376027 512567 376061
rect 512601 376027 512635 376061
rect 512669 376027 512703 376061
rect 512737 376027 512771 376061
rect 512805 376027 512839 376061
rect 512873 376027 512907 376061
rect 512941 376027 512975 376061
rect 513009 376027 513043 376061
rect 513077 376027 513111 376061
rect 513145 376027 513179 376061
rect 513213 376027 513247 376061
rect 513281 376027 513315 376061
rect 513349 376027 513383 376061
rect 513417 376027 513433 376061
rect 512143 376015 513433 376027
rect 504623 375603 505913 375615
rect 504623 375569 504639 375603
rect 504673 375569 504707 375603
rect 504741 375569 504775 375603
rect 504809 375569 504843 375603
rect 504877 375569 504911 375603
rect 504945 375569 504979 375603
rect 505013 375569 505047 375603
rect 505081 375569 505115 375603
rect 505149 375569 505183 375603
rect 505217 375569 505251 375603
rect 505285 375569 505319 375603
rect 505353 375569 505387 375603
rect 505421 375569 505455 375603
rect 505489 375569 505523 375603
rect 505557 375569 505591 375603
rect 505625 375569 505659 375603
rect 505693 375569 505727 375603
rect 505761 375569 505795 375603
rect 505829 375569 505863 375603
rect 505897 375569 505913 375603
rect 504623 375557 505913 375569
rect 493343 374963 494633 374975
rect 493343 374929 493359 374963
rect 493393 374929 493427 374963
rect 493461 374929 493495 374963
rect 493529 374929 493563 374963
rect 493597 374929 493631 374963
rect 493665 374929 493699 374963
rect 493733 374929 493767 374963
rect 493801 374929 493835 374963
rect 493869 374929 493903 374963
rect 493937 374929 493971 374963
rect 494005 374929 494039 374963
rect 494073 374929 494107 374963
rect 494141 374929 494175 374963
rect 494209 374929 494243 374963
rect 494277 374929 494311 374963
rect 494345 374929 494379 374963
rect 494413 374929 494447 374963
rect 494481 374929 494515 374963
rect 494549 374929 494583 374963
rect 494617 374929 494633 374963
rect 493343 374917 494633 374929
rect 497103 375145 498393 375157
rect 497103 375111 497119 375145
rect 497153 375111 497187 375145
rect 497221 375111 497255 375145
rect 497289 375111 497323 375145
rect 497357 375111 497391 375145
rect 497425 375111 497459 375145
rect 497493 375111 497527 375145
rect 497561 375111 497595 375145
rect 497629 375111 497663 375145
rect 497697 375111 497731 375145
rect 497765 375111 497799 375145
rect 497833 375111 497867 375145
rect 497901 375111 497935 375145
rect 497969 375111 498003 375145
rect 498037 375111 498071 375145
rect 498105 375111 498139 375145
rect 498173 375111 498207 375145
rect 498241 375111 498275 375145
rect 498309 375111 498343 375145
rect 498377 375111 498393 375145
rect 497103 375099 498393 375111
rect 493343 374505 494633 374517
rect 493343 374471 493359 374505
rect 493393 374471 493427 374505
rect 493461 374471 493495 374505
rect 493529 374471 493563 374505
rect 493597 374471 493631 374505
rect 493665 374471 493699 374505
rect 493733 374471 493767 374505
rect 493801 374471 493835 374505
rect 493869 374471 493903 374505
rect 493937 374471 493971 374505
rect 494005 374471 494039 374505
rect 494073 374471 494107 374505
rect 494141 374471 494175 374505
rect 494209 374471 494243 374505
rect 494277 374471 494311 374505
rect 494345 374471 494379 374505
rect 494413 374471 494447 374505
rect 494481 374471 494515 374505
rect 494549 374471 494583 374505
rect 494617 374471 494633 374505
rect 493343 374459 494633 374471
rect 512143 375603 513433 375615
rect 512143 375569 512159 375603
rect 512193 375569 512227 375603
rect 512261 375569 512295 375603
rect 512329 375569 512363 375603
rect 512397 375569 512431 375603
rect 512465 375569 512499 375603
rect 512533 375569 512567 375603
rect 512601 375569 512635 375603
rect 512669 375569 512703 375603
rect 512737 375569 512771 375603
rect 512805 375569 512839 375603
rect 512873 375569 512907 375603
rect 512941 375569 512975 375603
rect 513009 375569 513043 375603
rect 513077 375569 513111 375603
rect 513145 375569 513179 375603
rect 513213 375569 513247 375603
rect 513281 375569 513315 375603
rect 513349 375569 513383 375603
rect 513417 375569 513433 375603
rect 512143 375557 513433 375569
rect 504623 375145 505913 375157
rect 504623 375111 504639 375145
rect 504673 375111 504707 375145
rect 504741 375111 504775 375145
rect 504809 375111 504843 375145
rect 504877 375111 504911 375145
rect 504945 375111 504979 375145
rect 505013 375111 505047 375145
rect 505081 375111 505115 375145
rect 505149 375111 505183 375145
rect 505217 375111 505251 375145
rect 505285 375111 505319 375145
rect 505353 375111 505387 375145
rect 505421 375111 505455 375145
rect 505489 375111 505523 375145
rect 505557 375111 505591 375145
rect 505625 375111 505659 375145
rect 505693 375111 505727 375145
rect 505761 375111 505795 375145
rect 505829 375111 505863 375145
rect 505897 375111 505913 375145
rect 504623 375099 505913 375111
rect 497103 374687 498393 374699
rect 497103 374653 497119 374687
rect 497153 374653 497187 374687
rect 497221 374653 497255 374687
rect 497289 374653 497323 374687
rect 497357 374653 497391 374687
rect 497425 374653 497459 374687
rect 497493 374653 497527 374687
rect 497561 374653 497595 374687
rect 497629 374653 497663 374687
rect 497697 374653 497731 374687
rect 497765 374653 497799 374687
rect 497833 374653 497867 374687
rect 497901 374653 497935 374687
rect 497969 374653 498003 374687
rect 498037 374653 498071 374687
rect 498105 374653 498139 374687
rect 498173 374653 498207 374687
rect 498241 374653 498275 374687
rect 498309 374653 498343 374687
rect 498377 374653 498393 374687
rect 497103 374641 498393 374653
rect 493343 374047 494633 374059
rect 493343 374013 493359 374047
rect 493393 374013 493427 374047
rect 493461 374013 493495 374047
rect 493529 374013 493563 374047
rect 493597 374013 493631 374047
rect 493665 374013 493699 374047
rect 493733 374013 493767 374047
rect 493801 374013 493835 374047
rect 493869 374013 493903 374047
rect 493937 374013 493971 374047
rect 494005 374013 494039 374047
rect 494073 374013 494107 374047
rect 494141 374013 494175 374047
rect 494209 374013 494243 374047
rect 494277 374013 494311 374047
rect 494345 374013 494379 374047
rect 494413 374013 494447 374047
rect 494481 374013 494515 374047
rect 494549 374013 494583 374047
rect 494617 374013 494633 374047
rect 493343 374001 494633 374013
rect 497103 374229 498393 374241
rect 497103 374195 497119 374229
rect 497153 374195 497187 374229
rect 497221 374195 497255 374229
rect 497289 374195 497323 374229
rect 497357 374195 497391 374229
rect 497425 374195 497459 374229
rect 497493 374195 497527 374229
rect 497561 374195 497595 374229
rect 497629 374195 497663 374229
rect 497697 374195 497731 374229
rect 497765 374195 497799 374229
rect 497833 374195 497867 374229
rect 497901 374195 497935 374229
rect 497969 374195 498003 374229
rect 498037 374195 498071 374229
rect 498105 374195 498139 374229
rect 498173 374195 498207 374229
rect 498241 374195 498275 374229
rect 498309 374195 498343 374229
rect 498377 374195 498393 374229
rect 497103 374183 498393 374195
rect 493343 373589 494633 373601
rect 493343 373555 493359 373589
rect 493393 373555 493427 373589
rect 493461 373555 493495 373589
rect 493529 373555 493563 373589
rect 493597 373555 493631 373589
rect 493665 373555 493699 373589
rect 493733 373555 493767 373589
rect 493801 373555 493835 373589
rect 493869 373555 493903 373589
rect 493937 373555 493971 373589
rect 494005 373555 494039 373589
rect 494073 373555 494107 373589
rect 494141 373555 494175 373589
rect 494209 373555 494243 373589
rect 494277 373555 494311 373589
rect 494345 373555 494379 373589
rect 494413 373555 494447 373589
rect 494481 373555 494515 373589
rect 494549 373555 494583 373589
rect 494617 373555 494633 373589
rect 493343 373543 494633 373555
rect 512143 375145 513433 375157
rect 512143 375111 512159 375145
rect 512193 375111 512227 375145
rect 512261 375111 512295 375145
rect 512329 375111 512363 375145
rect 512397 375111 512431 375145
rect 512465 375111 512499 375145
rect 512533 375111 512567 375145
rect 512601 375111 512635 375145
rect 512669 375111 512703 375145
rect 512737 375111 512771 375145
rect 512805 375111 512839 375145
rect 512873 375111 512907 375145
rect 512941 375111 512975 375145
rect 513009 375111 513043 375145
rect 513077 375111 513111 375145
rect 513145 375111 513179 375145
rect 513213 375111 513247 375145
rect 513281 375111 513315 375145
rect 513349 375111 513383 375145
rect 513417 375111 513433 375145
rect 512143 375099 513433 375111
rect 504623 374687 505913 374699
rect 504623 374653 504639 374687
rect 504673 374653 504707 374687
rect 504741 374653 504775 374687
rect 504809 374653 504843 374687
rect 504877 374653 504911 374687
rect 504945 374653 504979 374687
rect 505013 374653 505047 374687
rect 505081 374653 505115 374687
rect 505149 374653 505183 374687
rect 505217 374653 505251 374687
rect 505285 374653 505319 374687
rect 505353 374653 505387 374687
rect 505421 374653 505455 374687
rect 505489 374653 505523 374687
rect 505557 374653 505591 374687
rect 505625 374653 505659 374687
rect 505693 374653 505727 374687
rect 505761 374653 505795 374687
rect 505829 374653 505863 374687
rect 505897 374653 505913 374687
rect 504623 374641 505913 374653
rect 497103 373771 498393 373783
rect 497103 373737 497119 373771
rect 497153 373737 497187 373771
rect 497221 373737 497255 373771
rect 497289 373737 497323 373771
rect 497357 373737 497391 373771
rect 497425 373737 497459 373771
rect 497493 373737 497527 373771
rect 497561 373737 497595 373771
rect 497629 373737 497663 373771
rect 497697 373737 497731 373771
rect 497765 373737 497799 373771
rect 497833 373737 497867 373771
rect 497901 373737 497935 373771
rect 497969 373737 498003 373771
rect 498037 373737 498071 373771
rect 498105 373737 498139 373771
rect 498173 373737 498207 373771
rect 498241 373737 498275 373771
rect 498309 373737 498343 373771
rect 498377 373737 498393 373771
rect 497103 373725 498393 373737
rect 523423 377253 524713 377265
rect 523423 377219 523439 377253
rect 523473 377219 523507 377253
rect 523541 377219 523575 377253
rect 523609 377219 523643 377253
rect 523677 377219 523711 377253
rect 523745 377219 523779 377253
rect 523813 377219 523847 377253
rect 523881 377219 523915 377253
rect 523949 377219 523983 377253
rect 524017 377219 524051 377253
rect 524085 377219 524119 377253
rect 524153 377219 524187 377253
rect 524221 377219 524255 377253
rect 524289 377219 524323 377253
rect 524357 377219 524391 377253
rect 524425 377219 524459 377253
rect 524493 377219 524527 377253
rect 524561 377219 524595 377253
rect 524629 377219 524663 377253
rect 524697 377219 524713 377253
rect 523423 377207 524713 377219
rect 523423 376795 524713 376807
rect 523423 376761 523439 376795
rect 523473 376761 523507 376795
rect 523541 376761 523575 376795
rect 523609 376761 523643 376795
rect 523677 376761 523711 376795
rect 523745 376761 523779 376795
rect 523813 376761 523847 376795
rect 523881 376761 523915 376795
rect 523949 376761 523983 376795
rect 524017 376761 524051 376795
rect 524085 376761 524119 376795
rect 524153 376761 524187 376795
rect 524221 376761 524255 376795
rect 524289 376761 524323 376795
rect 524357 376761 524391 376795
rect 524425 376761 524459 376795
rect 524493 376761 524527 376795
rect 524561 376761 524595 376795
rect 524629 376761 524663 376795
rect 524697 376761 524713 376795
rect 523423 376749 524713 376761
rect 523423 376337 524713 376349
rect 523423 376303 523439 376337
rect 523473 376303 523507 376337
rect 523541 376303 523575 376337
rect 523609 376303 523643 376337
rect 523677 376303 523711 376337
rect 523745 376303 523779 376337
rect 523813 376303 523847 376337
rect 523881 376303 523915 376337
rect 523949 376303 523983 376337
rect 524017 376303 524051 376337
rect 524085 376303 524119 376337
rect 524153 376303 524187 376337
rect 524221 376303 524255 376337
rect 524289 376303 524323 376337
rect 524357 376303 524391 376337
rect 524425 376303 524459 376337
rect 524493 376303 524527 376337
rect 524561 376303 524595 376337
rect 524629 376303 524663 376337
rect 524697 376303 524713 376337
rect 523423 376291 524713 376303
rect 523423 375879 524713 375891
rect 523423 375845 523439 375879
rect 523473 375845 523507 375879
rect 523541 375845 523575 375879
rect 523609 375845 523643 375879
rect 523677 375845 523711 375879
rect 523745 375845 523779 375879
rect 523813 375845 523847 375879
rect 523881 375845 523915 375879
rect 523949 375845 523983 375879
rect 524017 375845 524051 375879
rect 524085 375845 524119 375879
rect 524153 375845 524187 375879
rect 524221 375845 524255 375879
rect 524289 375845 524323 375879
rect 524357 375845 524391 375879
rect 524425 375845 524459 375879
rect 524493 375845 524527 375879
rect 524561 375845 524595 375879
rect 524629 375845 524663 375879
rect 524697 375845 524713 375879
rect 523423 375833 524713 375845
rect 523423 375421 524713 375433
rect 523423 375387 523439 375421
rect 523473 375387 523507 375421
rect 523541 375387 523575 375421
rect 523609 375387 523643 375421
rect 523677 375387 523711 375421
rect 523745 375387 523779 375421
rect 523813 375387 523847 375421
rect 523881 375387 523915 375421
rect 523949 375387 523983 375421
rect 524017 375387 524051 375421
rect 524085 375387 524119 375421
rect 524153 375387 524187 375421
rect 524221 375387 524255 375421
rect 524289 375387 524323 375421
rect 524357 375387 524391 375421
rect 524425 375387 524459 375421
rect 524493 375387 524527 375421
rect 524561 375387 524595 375421
rect 524629 375387 524663 375421
rect 524697 375387 524713 375421
rect 523423 375375 524713 375387
rect 523423 374963 524713 374975
rect 523423 374929 523439 374963
rect 523473 374929 523507 374963
rect 523541 374929 523575 374963
rect 523609 374929 523643 374963
rect 523677 374929 523711 374963
rect 523745 374929 523779 374963
rect 523813 374929 523847 374963
rect 523881 374929 523915 374963
rect 523949 374929 523983 374963
rect 524017 374929 524051 374963
rect 524085 374929 524119 374963
rect 524153 374929 524187 374963
rect 524221 374929 524255 374963
rect 524289 374929 524323 374963
rect 524357 374929 524391 374963
rect 524425 374929 524459 374963
rect 524493 374929 524527 374963
rect 524561 374929 524595 374963
rect 524629 374929 524663 374963
rect 524697 374929 524713 374963
rect 523423 374917 524713 374929
rect 512143 374687 513433 374699
rect 512143 374653 512159 374687
rect 512193 374653 512227 374687
rect 512261 374653 512295 374687
rect 512329 374653 512363 374687
rect 512397 374653 512431 374687
rect 512465 374653 512499 374687
rect 512533 374653 512567 374687
rect 512601 374653 512635 374687
rect 512669 374653 512703 374687
rect 512737 374653 512771 374687
rect 512805 374653 512839 374687
rect 512873 374653 512907 374687
rect 512941 374653 512975 374687
rect 513009 374653 513043 374687
rect 513077 374653 513111 374687
rect 513145 374653 513179 374687
rect 513213 374653 513247 374687
rect 513281 374653 513315 374687
rect 513349 374653 513383 374687
rect 513417 374653 513433 374687
rect 512143 374641 513433 374653
rect 493343 373131 494633 373143
rect 493343 373097 493359 373131
rect 493393 373097 493427 373131
rect 493461 373097 493495 373131
rect 493529 373097 493563 373131
rect 493597 373097 493631 373131
rect 493665 373097 493699 373131
rect 493733 373097 493767 373131
rect 493801 373097 493835 373131
rect 493869 373097 493903 373131
rect 493937 373097 493971 373131
rect 494005 373097 494039 373131
rect 494073 373097 494107 373131
rect 494141 373097 494175 373131
rect 494209 373097 494243 373131
rect 494277 373097 494311 373131
rect 494345 373097 494379 373131
rect 494413 373097 494447 373131
rect 494481 373097 494515 373131
rect 494549 373097 494583 373131
rect 494617 373097 494633 373131
rect 493343 373085 494633 373097
rect 497103 373313 498393 373325
rect 497103 373279 497119 373313
rect 497153 373279 497187 373313
rect 497221 373279 497255 373313
rect 497289 373279 497323 373313
rect 497357 373279 497391 373313
rect 497425 373279 497459 373313
rect 497493 373279 497527 373313
rect 497561 373279 497595 373313
rect 497629 373279 497663 373313
rect 497697 373279 497731 373313
rect 497765 373279 497799 373313
rect 497833 373279 497867 373313
rect 497901 373279 497935 373313
rect 497969 373279 498003 373313
rect 498037 373279 498071 373313
rect 498105 373279 498139 373313
rect 498173 373279 498207 373313
rect 498241 373279 498275 373313
rect 498309 373279 498343 373313
rect 498377 373279 498393 373313
rect 497103 373267 498393 373279
rect 497103 372855 498393 372867
rect 497103 372821 497119 372855
rect 497153 372821 497187 372855
rect 497221 372821 497255 372855
rect 497289 372821 497323 372855
rect 497357 372821 497391 372855
rect 497425 372821 497459 372855
rect 497493 372821 497527 372855
rect 497561 372821 497595 372855
rect 497629 372821 497663 372855
rect 497697 372821 497731 372855
rect 497765 372821 497799 372855
rect 497833 372821 497867 372855
rect 497901 372821 497935 372855
rect 497969 372821 498003 372855
rect 498037 372821 498071 372855
rect 498105 372821 498139 372855
rect 498173 372821 498207 372855
rect 498241 372821 498275 372855
rect 498309 372821 498343 372855
rect 498377 372821 498393 372855
rect 497103 372809 498393 372821
rect 493343 372673 494633 372685
rect 493343 372639 493359 372673
rect 493393 372639 493427 372673
rect 493461 372639 493495 372673
rect 493529 372639 493563 372673
rect 493597 372639 493631 372673
rect 493665 372639 493699 372673
rect 493733 372639 493767 372673
rect 493801 372639 493835 372673
rect 493869 372639 493903 372673
rect 493937 372639 493971 372673
rect 494005 372639 494039 372673
rect 494073 372639 494107 372673
rect 494141 372639 494175 372673
rect 494209 372639 494243 372673
rect 494277 372639 494311 372673
rect 494345 372639 494379 372673
rect 494413 372639 494447 372673
rect 494481 372639 494515 372673
rect 494549 372639 494583 372673
rect 494617 372639 494633 372673
rect 493343 372627 494633 372639
rect 497103 372397 498393 372409
rect 497103 372363 497119 372397
rect 497153 372363 497187 372397
rect 497221 372363 497255 372397
rect 497289 372363 497323 372397
rect 497357 372363 497391 372397
rect 497425 372363 497459 372397
rect 497493 372363 497527 372397
rect 497561 372363 497595 372397
rect 497629 372363 497663 372397
rect 497697 372363 497731 372397
rect 497765 372363 497799 372397
rect 497833 372363 497867 372397
rect 497901 372363 497935 372397
rect 497969 372363 498003 372397
rect 498037 372363 498071 372397
rect 498105 372363 498139 372397
rect 498173 372363 498207 372397
rect 498241 372363 498275 372397
rect 498309 372363 498343 372397
rect 498377 372363 498393 372397
rect 497103 372351 498393 372363
rect 493343 372215 494633 372227
rect 493343 372181 493359 372215
rect 493393 372181 493427 372215
rect 493461 372181 493495 372215
rect 493529 372181 493563 372215
rect 493597 372181 493631 372215
rect 493665 372181 493699 372215
rect 493733 372181 493767 372215
rect 493801 372181 493835 372215
rect 493869 372181 493903 372215
rect 493937 372181 493971 372215
rect 494005 372181 494039 372215
rect 494073 372181 494107 372215
rect 494141 372181 494175 372215
rect 494209 372181 494243 372215
rect 494277 372181 494311 372215
rect 494345 372181 494379 372215
rect 494413 372181 494447 372215
rect 494481 372181 494515 372215
rect 494549 372181 494583 372215
rect 494617 372181 494633 372215
rect 493343 372169 494633 372181
rect 501228 372786 501908 372840
rect 501228 372752 501280 372786
rect 501314 372752 501370 372786
rect 501404 372752 501460 372786
rect 501494 372752 501550 372786
rect 501584 372752 501640 372786
rect 501674 372752 501730 372786
rect 501764 372752 501820 372786
rect 501854 372752 501908 372786
rect 501228 372696 501908 372752
rect 501228 372662 501280 372696
rect 501314 372662 501370 372696
rect 501404 372662 501460 372696
rect 501494 372662 501550 372696
rect 501584 372662 501640 372696
rect 501674 372662 501730 372696
rect 501764 372662 501820 372696
rect 501854 372662 501908 372696
rect 501228 372606 501908 372662
rect 501228 372572 501280 372606
rect 501314 372572 501370 372606
rect 501404 372572 501460 372606
rect 501494 372572 501550 372606
rect 501584 372572 501640 372606
rect 501674 372572 501730 372606
rect 501764 372572 501820 372606
rect 501854 372572 501908 372606
rect 501228 372516 501908 372572
rect 501228 372482 501280 372516
rect 501314 372482 501370 372516
rect 501404 372482 501460 372516
rect 501494 372482 501550 372516
rect 501584 372482 501640 372516
rect 501674 372482 501730 372516
rect 501764 372482 501820 372516
rect 501854 372482 501908 372516
rect 501228 372426 501908 372482
rect 501228 372392 501280 372426
rect 501314 372392 501370 372426
rect 501404 372392 501460 372426
rect 501494 372392 501550 372426
rect 501584 372392 501640 372426
rect 501674 372392 501730 372426
rect 501764 372392 501820 372426
rect 501854 372392 501908 372426
rect 501228 372336 501908 372392
rect 501228 372302 501280 372336
rect 501314 372302 501370 372336
rect 501404 372302 501460 372336
rect 501494 372302 501550 372336
rect 501584 372302 501640 372336
rect 501674 372302 501730 372336
rect 501764 372302 501820 372336
rect 501854 372302 501908 372336
rect 501228 372246 501908 372302
rect 501228 372212 501280 372246
rect 501314 372212 501370 372246
rect 501404 372212 501460 372246
rect 501494 372212 501550 372246
rect 501584 372212 501640 372246
rect 501674 372212 501730 372246
rect 501764 372212 501820 372246
rect 501854 372212 501908 372246
rect 501228 372160 501908 372212
rect 493343 371757 494633 371769
rect 493343 371723 493359 371757
rect 493393 371723 493427 371757
rect 493461 371723 493495 371757
rect 493529 371723 493563 371757
rect 493597 371723 493631 371757
rect 493665 371723 493699 371757
rect 493733 371723 493767 371757
rect 493801 371723 493835 371757
rect 493869 371723 493903 371757
rect 493937 371723 493971 371757
rect 494005 371723 494039 371757
rect 494073 371723 494107 371757
rect 494141 371723 494175 371757
rect 494209 371723 494243 371757
rect 494277 371723 494311 371757
rect 494345 371723 494379 371757
rect 494413 371723 494447 371757
rect 494481 371723 494515 371757
rect 494549 371723 494583 371757
rect 494617 371723 494633 371757
rect 493343 371711 494633 371723
rect 493343 371299 494633 371311
rect 493343 371265 493359 371299
rect 493393 371265 493427 371299
rect 493461 371265 493495 371299
rect 493529 371265 493563 371299
rect 493597 371265 493631 371299
rect 493665 371265 493699 371299
rect 493733 371265 493767 371299
rect 493801 371265 493835 371299
rect 493869 371265 493903 371299
rect 493937 371265 493971 371299
rect 494005 371265 494039 371299
rect 494073 371265 494107 371299
rect 494141 371265 494175 371299
rect 494209 371265 494243 371299
rect 494277 371265 494311 371299
rect 494345 371265 494379 371299
rect 494413 371265 494447 371299
rect 494481 371265 494515 371299
rect 494549 371265 494583 371299
rect 494617 371265 494633 371299
rect 493343 371253 494633 371265
rect 493343 370841 494633 370853
rect 493343 370807 493359 370841
rect 493393 370807 493427 370841
rect 493461 370807 493495 370841
rect 493529 370807 493563 370841
rect 493597 370807 493631 370841
rect 493665 370807 493699 370841
rect 493733 370807 493767 370841
rect 493801 370807 493835 370841
rect 493869 370807 493903 370841
rect 493937 370807 493971 370841
rect 494005 370807 494039 370841
rect 494073 370807 494107 370841
rect 494141 370807 494175 370841
rect 494209 370807 494243 370841
rect 494277 370807 494311 370841
rect 494345 370807 494379 370841
rect 494413 370807 494447 370841
rect 494481 370807 494515 370841
rect 494549 370807 494583 370841
rect 494617 370807 494633 370841
rect 493343 370795 494633 370807
rect 493343 370383 494633 370395
rect 493343 370349 493359 370383
rect 493393 370349 493427 370383
rect 493461 370349 493495 370383
rect 493529 370349 493563 370383
rect 493597 370349 493631 370383
rect 493665 370349 493699 370383
rect 493733 370349 493767 370383
rect 493801 370349 493835 370383
rect 493869 370349 493903 370383
rect 493937 370349 493971 370383
rect 494005 370349 494039 370383
rect 494073 370349 494107 370383
rect 494141 370349 494175 370383
rect 494209 370349 494243 370383
rect 494277 370349 494311 370383
rect 494345 370349 494379 370383
rect 494413 370349 494447 370383
rect 494481 370349 494515 370383
rect 494549 370349 494583 370383
rect 494617 370349 494633 370383
rect 493343 370337 494633 370349
rect 493343 369925 494633 369937
rect 493343 369891 493359 369925
rect 493393 369891 493427 369925
rect 493461 369891 493495 369925
rect 493529 369891 493563 369925
rect 493597 369891 493631 369925
rect 493665 369891 493699 369925
rect 493733 369891 493767 369925
rect 493801 369891 493835 369925
rect 493869 369891 493903 369925
rect 493937 369891 493971 369925
rect 494005 369891 494039 369925
rect 494073 369891 494107 369925
rect 494141 369891 494175 369925
rect 494209 369891 494243 369925
rect 494277 369891 494311 369925
rect 494345 369891 494379 369925
rect 494413 369891 494447 369925
rect 494481 369891 494515 369925
rect 494549 369891 494583 369925
rect 494617 369891 494633 369925
rect 493343 369879 494633 369891
rect 493343 369467 494633 369479
rect 493343 369433 493359 369467
rect 493393 369433 493427 369467
rect 493461 369433 493495 369467
rect 493529 369433 493563 369467
rect 493597 369433 493631 369467
rect 493665 369433 493699 369467
rect 493733 369433 493767 369467
rect 493801 369433 493835 369467
rect 493869 369433 493903 369467
rect 493937 369433 493971 369467
rect 494005 369433 494039 369467
rect 494073 369433 494107 369467
rect 494141 369433 494175 369467
rect 494209 369433 494243 369467
rect 494277 369433 494311 369467
rect 494345 369433 494379 369467
rect 494413 369433 494447 369467
rect 494481 369433 494515 369467
rect 494549 369433 494583 369467
rect 494617 369433 494633 369467
rect 493343 369421 494633 369433
rect 493343 369009 494633 369021
rect 493343 368975 493359 369009
rect 493393 368975 493427 369009
rect 493461 368975 493495 369009
rect 493529 368975 493563 369009
rect 493597 368975 493631 369009
rect 493665 368975 493699 369009
rect 493733 368975 493767 369009
rect 493801 368975 493835 369009
rect 493869 368975 493903 369009
rect 493937 368975 493971 369009
rect 494005 368975 494039 369009
rect 494073 368975 494107 369009
rect 494141 368975 494175 369009
rect 494209 368975 494243 369009
rect 494277 368975 494311 369009
rect 494345 368975 494379 369009
rect 494413 368975 494447 369009
rect 494481 368975 494515 369009
rect 494549 368975 494583 369009
rect 494617 368975 494633 369009
rect 493343 368963 494633 368975
rect 493343 368551 494633 368563
rect 493343 368517 493359 368551
rect 493393 368517 493427 368551
rect 493461 368517 493495 368551
rect 493529 368517 493563 368551
rect 493597 368517 493631 368551
rect 493665 368517 493699 368551
rect 493733 368517 493767 368551
rect 493801 368517 493835 368551
rect 493869 368517 493903 368551
rect 493937 368517 493971 368551
rect 494005 368517 494039 368551
rect 494073 368517 494107 368551
rect 494141 368517 494175 368551
rect 494209 368517 494243 368551
rect 494277 368517 494311 368551
rect 494345 368517 494379 368551
rect 494413 368517 494447 368551
rect 494481 368517 494515 368551
rect 494549 368517 494583 368551
rect 494617 368517 494633 368551
rect 493343 368505 494633 368517
rect 493343 368093 494633 368105
rect 493343 368059 493359 368093
rect 493393 368059 493427 368093
rect 493461 368059 493495 368093
rect 493529 368059 493563 368093
rect 493597 368059 493631 368093
rect 493665 368059 493699 368093
rect 493733 368059 493767 368093
rect 493801 368059 493835 368093
rect 493869 368059 493903 368093
rect 493937 368059 493971 368093
rect 494005 368059 494039 368093
rect 494073 368059 494107 368093
rect 494141 368059 494175 368093
rect 494209 368059 494243 368093
rect 494277 368059 494311 368093
rect 494345 368059 494379 368093
rect 494413 368059 494447 368093
rect 494481 368059 494515 368093
rect 494549 368059 494583 368093
rect 494617 368059 494633 368093
rect 493343 368047 494633 368059
rect 493343 367635 494633 367647
rect 493343 367601 493359 367635
rect 493393 367601 493427 367635
rect 493461 367601 493495 367635
rect 493529 367601 493563 367635
rect 493597 367601 493631 367635
rect 493665 367601 493699 367635
rect 493733 367601 493767 367635
rect 493801 367601 493835 367635
rect 493869 367601 493903 367635
rect 493937 367601 493971 367635
rect 494005 367601 494039 367635
rect 494073 367601 494107 367635
rect 494141 367601 494175 367635
rect 494209 367601 494243 367635
rect 494277 367601 494311 367635
rect 494345 367601 494379 367635
rect 494413 367601 494447 367635
rect 494481 367601 494515 367635
rect 494549 367601 494583 367635
rect 494617 367601 494633 367635
rect 493343 367589 494633 367601
rect 493343 367177 494633 367189
rect 493343 367143 493359 367177
rect 493393 367143 493427 367177
rect 493461 367143 493495 367177
rect 493529 367143 493563 367177
rect 493597 367143 493631 367177
rect 493665 367143 493699 367177
rect 493733 367143 493767 367177
rect 493801 367143 493835 367177
rect 493869 367143 493903 367177
rect 493937 367143 493971 367177
rect 494005 367143 494039 367177
rect 494073 367143 494107 367177
rect 494141 367143 494175 367177
rect 494209 367143 494243 367177
rect 494277 367143 494311 367177
rect 494345 367143 494379 367177
rect 494413 367143 494447 367177
rect 494481 367143 494515 367177
rect 494549 367143 494583 367177
rect 494617 367143 494633 367177
rect 493343 367131 494633 367143
rect 493343 366719 494633 366731
rect 493343 366685 493359 366719
rect 493393 366685 493427 366719
rect 493461 366685 493495 366719
rect 493529 366685 493563 366719
rect 493597 366685 493631 366719
rect 493665 366685 493699 366719
rect 493733 366685 493767 366719
rect 493801 366685 493835 366719
rect 493869 366685 493903 366719
rect 493937 366685 493971 366719
rect 494005 366685 494039 366719
rect 494073 366685 494107 366719
rect 494141 366685 494175 366719
rect 494209 366685 494243 366719
rect 494277 366685 494311 366719
rect 494345 366685 494379 366719
rect 494413 366685 494447 366719
rect 494481 366685 494515 366719
rect 494549 366685 494583 366719
rect 494617 366685 494633 366719
rect 493343 366673 494633 366685
rect 493343 366261 494633 366273
rect 493343 366227 493359 366261
rect 493393 366227 493427 366261
rect 493461 366227 493495 366261
rect 493529 366227 493563 366261
rect 493597 366227 493631 366261
rect 493665 366227 493699 366261
rect 493733 366227 493767 366261
rect 493801 366227 493835 366261
rect 493869 366227 493903 366261
rect 493937 366227 493971 366261
rect 494005 366227 494039 366261
rect 494073 366227 494107 366261
rect 494141 366227 494175 366261
rect 494209 366227 494243 366261
rect 494277 366227 494311 366261
rect 494345 366227 494379 366261
rect 494413 366227 494447 366261
rect 494481 366227 494515 366261
rect 494549 366227 494583 366261
rect 494617 366227 494633 366261
rect 493343 366215 494633 366227
rect 493343 365803 494633 365815
rect 493343 365769 493359 365803
rect 493393 365769 493427 365803
rect 493461 365769 493495 365803
rect 493529 365769 493563 365803
rect 493597 365769 493631 365803
rect 493665 365769 493699 365803
rect 493733 365769 493767 365803
rect 493801 365769 493835 365803
rect 493869 365769 493903 365803
rect 493937 365769 493971 365803
rect 494005 365769 494039 365803
rect 494073 365769 494107 365803
rect 494141 365769 494175 365803
rect 494209 365769 494243 365803
rect 494277 365769 494311 365803
rect 494345 365769 494379 365803
rect 494413 365769 494447 365803
rect 494481 365769 494515 365803
rect 494549 365769 494583 365803
rect 494617 365769 494633 365803
rect 493343 365757 494633 365769
rect 493343 365345 494633 365357
rect 493343 365311 493359 365345
rect 493393 365311 493427 365345
rect 493461 365311 493495 365345
rect 493529 365311 493563 365345
rect 493597 365311 493631 365345
rect 493665 365311 493699 365345
rect 493733 365311 493767 365345
rect 493801 365311 493835 365345
rect 493869 365311 493903 365345
rect 493937 365311 493971 365345
rect 494005 365311 494039 365345
rect 494073 365311 494107 365345
rect 494141 365311 494175 365345
rect 494209 365311 494243 365345
rect 494277 365311 494311 365345
rect 494345 365311 494379 365345
rect 494413 365311 494447 365345
rect 494481 365311 494515 365345
rect 494549 365311 494583 365345
rect 494617 365311 494633 365345
rect 493343 365299 494633 365311
rect 493343 364887 494633 364899
rect 493343 364853 493359 364887
rect 493393 364853 493427 364887
rect 493461 364853 493495 364887
rect 493529 364853 493563 364887
rect 493597 364853 493631 364887
rect 493665 364853 493699 364887
rect 493733 364853 493767 364887
rect 493801 364853 493835 364887
rect 493869 364853 493903 364887
rect 493937 364853 493971 364887
rect 494005 364853 494039 364887
rect 494073 364853 494107 364887
rect 494141 364853 494175 364887
rect 494209 364853 494243 364887
rect 494277 364853 494311 364887
rect 494345 364853 494379 364887
rect 494413 364853 494447 364887
rect 494481 364853 494515 364887
rect 494549 364853 494583 364887
rect 494617 364853 494633 364887
rect 493343 364841 494633 364853
rect 493343 364429 494633 364441
rect 493343 364395 493359 364429
rect 493393 364395 493427 364429
rect 493461 364395 493495 364429
rect 493529 364395 493563 364429
rect 493597 364395 493631 364429
rect 493665 364395 493699 364429
rect 493733 364395 493767 364429
rect 493801 364395 493835 364429
rect 493869 364395 493903 364429
rect 493937 364395 493971 364429
rect 494005 364395 494039 364429
rect 494073 364395 494107 364429
rect 494141 364395 494175 364429
rect 494209 364395 494243 364429
rect 494277 364395 494311 364429
rect 494345 364395 494379 364429
rect 494413 364395 494447 364429
rect 494481 364395 494515 364429
rect 494549 364395 494583 364429
rect 494617 364395 494633 364429
rect 493343 364383 494633 364395
rect 493343 363971 494633 363983
rect 493343 363937 493359 363971
rect 493393 363937 493427 363971
rect 493461 363937 493495 363971
rect 493529 363937 493563 363971
rect 493597 363937 493631 363971
rect 493665 363937 493699 363971
rect 493733 363937 493767 363971
rect 493801 363937 493835 363971
rect 493869 363937 493903 363971
rect 493937 363937 493971 363971
rect 494005 363937 494039 363971
rect 494073 363937 494107 363971
rect 494141 363937 494175 363971
rect 494209 363937 494243 363971
rect 494277 363937 494311 363971
rect 494345 363937 494379 363971
rect 494413 363937 494447 363971
rect 494481 363937 494515 363971
rect 494549 363937 494583 363971
rect 494617 363937 494633 363971
rect 493343 363925 494633 363937
rect 493343 363513 494633 363525
rect 493343 363479 493359 363513
rect 493393 363479 493427 363513
rect 493461 363479 493495 363513
rect 493529 363479 493563 363513
rect 493597 363479 493631 363513
rect 493665 363479 493699 363513
rect 493733 363479 493767 363513
rect 493801 363479 493835 363513
rect 493869 363479 493903 363513
rect 493937 363479 493971 363513
rect 494005 363479 494039 363513
rect 494073 363479 494107 363513
rect 494141 363479 494175 363513
rect 494209 363479 494243 363513
rect 494277 363479 494311 363513
rect 494345 363479 494379 363513
rect 494413 363479 494447 363513
rect 494481 363479 494515 363513
rect 494549 363479 494583 363513
rect 494617 363479 494633 363513
rect 493343 363467 494633 363479
rect 493343 363055 494633 363067
rect 493343 363021 493359 363055
rect 493393 363021 493427 363055
rect 493461 363021 493495 363055
rect 493529 363021 493563 363055
rect 493597 363021 493631 363055
rect 493665 363021 493699 363055
rect 493733 363021 493767 363055
rect 493801 363021 493835 363055
rect 493869 363021 493903 363055
rect 493937 363021 493971 363055
rect 494005 363021 494039 363055
rect 494073 363021 494107 363055
rect 494141 363021 494175 363055
rect 494209 363021 494243 363055
rect 494277 363021 494311 363055
rect 494345 363021 494379 363055
rect 494413 363021 494447 363055
rect 494481 363021 494515 363055
rect 494549 363021 494583 363055
rect 494617 363021 494633 363055
rect 493343 363009 494633 363021
rect 493343 362597 494633 362609
rect 493343 362563 493359 362597
rect 493393 362563 493427 362597
rect 493461 362563 493495 362597
rect 493529 362563 493563 362597
rect 493597 362563 493631 362597
rect 493665 362563 493699 362597
rect 493733 362563 493767 362597
rect 493801 362563 493835 362597
rect 493869 362563 493903 362597
rect 493937 362563 493971 362597
rect 494005 362563 494039 362597
rect 494073 362563 494107 362597
rect 494141 362563 494175 362597
rect 494209 362563 494243 362597
rect 494277 362563 494311 362597
rect 494345 362563 494379 362597
rect 494413 362563 494447 362597
rect 494481 362563 494515 362597
rect 494549 362563 494583 362597
rect 494617 362563 494633 362597
rect 493343 362551 494633 362563
rect 497468 371610 498148 371664
rect 497468 371576 497520 371610
rect 497554 371576 497610 371610
rect 497644 371576 497700 371610
rect 497734 371576 497790 371610
rect 497824 371576 497880 371610
rect 497914 371576 497970 371610
rect 498004 371576 498060 371610
rect 498094 371576 498148 371610
rect 497468 371520 498148 371576
rect 497468 371486 497520 371520
rect 497554 371486 497610 371520
rect 497644 371486 497700 371520
rect 497734 371486 497790 371520
rect 497824 371486 497880 371520
rect 497914 371486 497970 371520
rect 498004 371486 498060 371520
rect 498094 371486 498148 371520
rect 497468 371430 498148 371486
rect 497468 371396 497520 371430
rect 497554 371396 497610 371430
rect 497644 371396 497700 371430
rect 497734 371396 497790 371430
rect 497824 371396 497880 371430
rect 497914 371396 497970 371430
rect 498004 371396 498060 371430
rect 498094 371396 498148 371430
rect 497468 371340 498148 371396
rect 497468 371306 497520 371340
rect 497554 371306 497610 371340
rect 497644 371306 497700 371340
rect 497734 371306 497790 371340
rect 497824 371306 497880 371340
rect 497914 371306 497970 371340
rect 498004 371306 498060 371340
rect 498094 371306 498148 371340
rect 497468 371250 498148 371306
rect 497468 371216 497520 371250
rect 497554 371216 497610 371250
rect 497644 371216 497700 371250
rect 497734 371216 497790 371250
rect 497824 371216 497880 371250
rect 497914 371216 497970 371250
rect 498004 371216 498060 371250
rect 498094 371216 498148 371250
rect 497468 371160 498148 371216
rect 497468 371126 497520 371160
rect 497554 371126 497610 371160
rect 497644 371126 497700 371160
rect 497734 371126 497790 371160
rect 497824 371126 497880 371160
rect 497914 371126 497970 371160
rect 498004 371126 498060 371160
rect 498094 371126 498148 371160
rect 497468 371070 498148 371126
rect 497468 371036 497520 371070
rect 497554 371036 497610 371070
rect 497644 371036 497700 371070
rect 497734 371036 497790 371070
rect 497824 371036 497880 371070
rect 497914 371036 497970 371070
rect 498004 371036 498060 371070
rect 498094 371036 498148 371070
rect 497468 370984 498148 371036
rect 497468 370270 498148 370324
rect 497468 370236 497520 370270
rect 497554 370236 497610 370270
rect 497644 370236 497700 370270
rect 497734 370236 497790 370270
rect 497824 370236 497880 370270
rect 497914 370236 497970 370270
rect 498004 370236 498060 370270
rect 498094 370236 498148 370270
rect 497468 370180 498148 370236
rect 497468 370146 497520 370180
rect 497554 370146 497610 370180
rect 497644 370146 497700 370180
rect 497734 370146 497790 370180
rect 497824 370146 497880 370180
rect 497914 370146 497970 370180
rect 498004 370146 498060 370180
rect 498094 370146 498148 370180
rect 497468 370090 498148 370146
rect 497468 370056 497520 370090
rect 497554 370056 497610 370090
rect 497644 370056 497700 370090
rect 497734 370056 497790 370090
rect 497824 370056 497880 370090
rect 497914 370056 497970 370090
rect 498004 370056 498060 370090
rect 498094 370056 498148 370090
rect 497468 370000 498148 370056
rect 497468 369966 497520 370000
rect 497554 369966 497610 370000
rect 497644 369966 497700 370000
rect 497734 369966 497790 370000
rect 497824 369966 497880 370000
rect 497914 369966 497970 370000
rect 498004 369966 498060 370000
rect 498094 369966 498148 370000
rect 497468 369910 498148 369966
rect 497468 369876 497520 369910
rect 497554 369876 497610 369910
rect 497644 369876 497700 369910
rect 497734 369876 497790 369910
rect 497824 369876 497880 369910
rect 497914 369876 497970 369910
rect 498004 369876 498060 369910
rect 498094 369876 498148 369910
rect 497468 369820 498148 369876
rect 497468 369786 497520 369820
rect 497554 369786 497610 369820
rect 497644 369786 497700 369820
rect 497734 369786 497790 369820
rect 497824 369786 497880 369820
rect 497914 369786 497970 369820
rect 498004 369786 498060 369820
rect 498094 369786 498148 369820
rect 497468 369730 498148 369786
rect 497468 369696 497520 369730
rect 497554 369696 497610 369730
rect 497644 369696 497700 369730
rect 497734 369696 497790 369730
rect 497824 369696 497880 369730
rect 497914 369696 497970 369730
rect 498004 369696 498060 369730
rect 498094 369696 498148 369730
rect 497468 369644 498148 369696
rect 497468 368930 498148 368984
rect 497468 368896 497520 368930
rect 497554 368896 497610 368930
rect 497644 368896 497700 368930
rect 497734 368896 497790 368930
rect 497824 368896 497880 368930
rect 497914 368896 497970 368930
rect 498004 368896 498060 368930
rect 498094 368896 498148 368930
rect 497468 368840 498148 368896
rect 497468 368806 497520 368840
rect 497554 368806 497610 368840
rect 497644 368806 497700 368840
rect 497734 368806 497790 368840
rect 497824 368806 497880 368840
rect 497914 368806 497970 368840
rect 498004 368806 498060 368840
rect 498094 368806 498148 368840
rect 497468 368750 498148 368806
rect 497468 368716 497520 368750
rect 497554 368716 497610 368750
rect 497644 368716 497700 368750
rect 497734 368716 497790 368750
rect 497824 368716 497880 368750
rect 497914 368716 497970 368750
rect 498004 368716 498060 368750
rect 498094 368716 498148 368750
rect 497468 368660 498148 368716
rect 497468 368626 497520 368660
rect 497554 368626 497610 368660
rect 497644 368626 497700 368660
rect 497734 368626 497790 368660
rect 497824 368626 497880 368660
rect 497914 368626 497970 368660
rect 498004 368626 498060 368660
rect 498094 368626 498148 368660
rect 497468 368570 498148 368626
rect 497468 368536 497520 368570
rect 497554 368536 497610 368570
rect 497644 368536 497700 368570
rect 497734 368536 497790 368570
rect 497824 368536 497880 368570
rect 497914 368536 497970 368570
rect 498004 368536 498060 368570
rect 498094 368536 498148 368570
rect 497468 368480 498148 368536
rect 497468 368446 497520 368480
rect 497554 368446 497610 368480
rect 497644 368446 497700 368480
rect 497734 368446 497790 368480
rect 497824 368446 497880 368480
rect 497914 368446 497970 368480
rect 498004 368446 498060 368480
rect 498094 368446 498148 368480
rect 497468 368390 498148 368446
rect 497468 368356 497520 368390
rect 497554 368356 497610 368390
rect 497644 368356 497700 368390
rect 497734 368356 497790 368390
rect 497824 368356 497880 368390
rect 497914 368356 497970 368390
rect 498004 368356 498060 368390
rect 498094 368356 498148 368390
rect 497468 368304 498148 368356
rect 497468 367590 498148 367644
rect 497468 367556 497520 367590
rect 497554 367556 497610 367590
rect 497644 367556 497700 367590
rect 497734 367556 497790 367590
rect 497824 367556 497880 367590
rect 497914 367556 497970 367590
rect 498004 367556 498060 367590
rect 498094 367556 498148 367590
rect 497468 367500 498148 367556
rect 497468 367466 497520 367500
rect 497554 367466 497610 367500
rect 497644 367466 497700 367500
rect 497734 367466 497790 367500
rect 497824 367466 497880 367500
rect 497914 367466 497970 367500
rect 498004 367466 498060 367500
rect 498094 367466 498148 367500
rect 497468 367410 498148 367466
rect 497468 367376 497520 367410
rect 497554 367376 497610 367410
rect 497644 367376 497700 367410
rect 497734 367376 497790 367410
rect 497824 367376 497880 367410
rect 497914 367376 497970 367410
rect 498004 367376 498060 367410
rect 498094 367376 498148 367410
rect 497468 367320 498148 367376
rect 497468 367286 497520 367320
rect 497554 367286 497610 367320
rect 497644 367286 497700 367320
rect 497734 367286 497790 367320
rect 497824 367286 497880 367320
rect 497914 367286 497970 367320
rect 498004 367286 498060 367320
rect 498094 367286 498148 367320
rect 497468 367230 498148 367286
rect 497468 367196 497520 367230
rect 497554 367196 497610 367230
rect 497644 367196 497700 367230
rect 497734 367196 497790 367230
rect 497824 367196 497880 367230
rect 497914 367196 497970 367230
rect 498004 367196 498060 367230
rect 498094 367196 498148 367230
rect 497468 367140 498148 367196
rect 497468 367106 497520 367140
rect 497554 367106 497610 367140
rect 497644 367106 497700 367140
rect 497734 367106 497790 367140
rect 497824 367106 497880 367140
rect 497914 367106 497970 367140
rect 498004 367106 498060 367140
rect 498094 367106 498148 367140
rect 497468 367050 498148 367106
rect 497468 367016 497520 367050
rect 497554 367016 497610 367050
rect 497644 367016 497700 367050
rect 497734 367016 497790 367050
rect 497824 367016 497880 367050
rect 497914 367016 497970 367050
rect 498004 367016 498060 367050
rect 498094 367016 498148 367050
rect 497468 366964 498148 367016
rect 497468 366250 498148 366304
rect 497468 366216 497520 366250
rect 497554 366216 497610 366250
rect 497644 366216 497700 366250
rect 497734 366216 497790 366250
rect 497824 366216 497880 366250
rect 497914 366216 497970 366250
rect 498004 366216 498060 366250
rect 498094 366216 498148 366250
rect 497468 366160 498148 366216
rect 497468 366126 497520 366160
rect 497554 366126 497610 366160
rect 497644 366126 497700 366160
rect 497734 366126 497790 366160
rect 497824 366126 497880 366160
rect 497914 366126 497970 366160
rect 498004 366126 498060 366160
rect 498094 366126 498148 366160
rect 497468 366070 498148 366126
rect 497468 366036 497520 366070
rect 497554 366036 497610 366070
rect 497644 366036 497700 366070
rect 497734 366036 497790 366070
rect 497824 366036 497880 366070
rect 497914 366036 497970 366070
rect 498004 366036 498060 366070
rect 498094 366036 498148 366070
rect 497468 365980 498148 366036
rect 497468 365946 497520 365980
rect 497554 365946 497610 365980
rect 497644 365946 497700 365980
rect 497734 365946 497790 365980
rect 497824 365946 497880 365980
rect 497914 365946 497970 365980
rect 498004 365946 498060 365980
rect 498094 365946 498148 365980
rect 497468 365890 498148 365946
rect 497468 365856 497520 365890
rect 497554 365856 497610 365890
rect 497644 365856 497700 365890
rect 497734 365856 497790 365890
rect 497824 365856 497880 365890
rect 497914 365856 497970 365890
rect 498004 365856 498060 365890
rect 498094 365856 498148 365890
rect 497468 365800 498148 365856
rect 497468 365766 497520 365800
rect 497554 365766 497610 365800
rect 497644 365766 497700 365800
rect 497734 365766 497790 365800
rect 497824 365766 497880 365800
rect 497914 365766 497970 365800
rect 498004 365766 498060 365800
rect 498094 365766 498148 365800
rect 497468 365710 498148 365766
rect 497468 365676 497520 365710
rect 497554 365676 497610 365710
rect 497644 365676 497700 365710
rect 497734 365676 497790 365710
rect 497824 365676 497880 365710
rect 497914 365676 497970 365710
rect 498004 365676 498060 365710
rect 498094 365676 498148 365710
rect 497468 365624 498148 365676
rect 497468 364910 498148 364964
rect 497468 364876 497520 364910
rect 497554 364876 497610 364910
rect 497644 364876 497700 364910
rect 497734 364876 497790 364910
rect 497824 364876 497880 364910
rect 497914 364876 497970 364910
rect 498004 364876 498060 364910
rect 498094 364876 498148 364910
rect 497468 364820 498148 364876
rect 497468 364786 497520 364820
rect 497554 364786 497610 364820
rect 497644 364786 497700 364820
rect 497734 364786 497790 364820
rect 497824 364786 497880 364820
rect 497914 364786 497970 364820
rect 498004 364786 498060 364820
rect 498094 364786 498148 364820
rect 497468 364730 498148 364786
rect 497468 364696 497520 364730
rect 497554 364696 497610 364730
rect 497644 364696 497700 364730
rect 497734 364696 497790 364730
rect 497824 364696 497880 364730
rect 497914 364696 497970 364730
rect 498004 364696 498060 364730
rect 498094 364696 498148 364730
rect 497468 364640 498148 364696
rect 497468 364606 497520 364640
rect 497554 364606 497610 364640
rect 497644 364606 497700 364640
rect 497734 364606 497790 364640
rect 497824 364606 497880 364640
rect 497914 364606 497970 364640
rect 498004 364606 498060 364640
rect 498094 364606 498148 364640
rect 497468 364550 498148 364606
rect 497468 364516 497520 364550
rect 497554 364516 497610 364550
rect 497644 364516 497700 364550
rect 497734 364516 497790 364550
rect 497824 364516 497880 364550
rect 497914 364516 497970 364550
rect 498004 364516 498060 364550
rect 498094 364516 498148 364550
rect 497468 364460 498148 364516
rect 497468 364426 497520 364460
rect 497554 364426 497610 364460
rect 497644 364426 497700 364460
rect 497734 364426 497790 364460
rect 497824 364426 497880 364460
rect 497914 364426 497970 364460
rect 498004 364426 498060 364460
rect 498094 364426 498148 364460
rect 497468 364370 498148 364426
rect 497468 364336 497520 364370
rect 497554 364336 497610 364370
rect 497644 364336 497700 364370
rect 497734 364336 497790 364370
rect 497824 364336 497880 364370
rect 497914 364336 497970 364370
rect 498004 364336 498060 364370
rect 498094 364336 498148 364370
rect 497468 364284 498148 364336
rect 497468 363570 498148 363624
rect 497468 363536 497520 363570
rect 497554 363536 497610 363570
rect 497644 363536 497700 363570
rect 497734 363536 497790 363570
rect 497824 363536 497880 363570
rect 497914 363536 497970 363570
rect 498004 363536 498060 363570
rect 498094 363536 498148 363570
rect 497468 363480 498148 363536
rect 497468 363446 497520 363480
rect 497554 363446 497610 363480
rect 497644 363446 497700 363480
rect 497734 363446 497790 363480
rect 497824 363446 497880 363480
rect 497914 363446 497970 363480
rect 498004 363446 498060 363480
rect 498094 363446 498148 363480
rect 497468 363390 498148 363446
rect 497468 363356 497520 363390
rect 497554 363356 497610 363390
rect 497644 363356 497700 363390
rect 497734 363356 497790 363390
rect 497824 363356 497880 363390
rect 497914 363356 497970 363390
rect 498004 363356 498060 363390
rect 498094 363356 498148 363390
rect 497468 363300 498148 363356
rect 497468 363266 497520 363300
rect 497554 363266 497610 363300
rect 497644 363266 497700 363300
rect 497734 363266 497790 363300
rect 497824 363266 497880 363300
rect 497914 363266 497970 363300
rect 498004 363266 498060 363300
rect 498094 363266 498148 363300
rect 497468 363210 498148 363266
rect 497468 363176 497520 363210
rect 497554 363176 497610 363210
rect 497644 363176 497700 363210
rect 497734 363176 497790 363210
rect 497824 363176 497880 363210
rect 497914 363176 497970 363210
rect 498004 363176 498060 363210
rect 498094 363176 498148 363210
rect 497468 363120 498148 363176
rect 497468 363086 497520 363120
rect 497554 363086 497610 363120
rect 497644 363086 497700 363120
rect 497734 363086 497790 363120
rect 497824 363086 497880 363120
rect 497914 363086 497970 363120
rect 498004 363086 498060 363120
rect 498094 363086 498148 363120
rect 497468 363030 498148 363086
rect 497468 362996 497520 363030
rect 497554 362996 497610 363030
rect 497644 362996 497700 363030
rect 497734 362996 497790 363030
rect 497824 362996 497880 363030
rect 497914 362996 497970 363030
rect 498004 362996 498060 363030
rect 498094 362996 498148 363030
rect 497468 362944 498148 362996
rect 501228 371446 501908 371500
rect 501228 371412 501280 371446
rect 501314 371412 501370 371446
rect 501404 371412 501460 371446
rect 501494 371412 501550 371446
rect 501584 371412 501640 371446
rect 501674 371412 501730 371446
rect 501764 371412 501820 371446
rect 501854 371412 501908 371446
rect 501228 371356 501908 371412
rect 501228 371322 501280 371356
rect 501314 371322 501370 371356
rect 501404 371322 501460 371356
rect 501494 371322 501550 371356
rect 501584 371322 501640 371356
rect 501674 371322 501730 371356
rect 501764 371322 501820 371356
rect 501854 371322 501908 371356
rect 501228 371266 501908 371322
rect 501228 371232 501280 371266
rect 501314 371232 501370 371266
rect 501404 371232 501460 371266
rect 501494 371232 501550 371266
rect 501584 371232 501640 371266
rect 501674 371232 501730 371266
rect 501764 371232 501820 371266
rect 501854 371232 501908 371266
rect 501228 371176 501908 371232
rect 501228 371142 501280 371176
rect 501314 371142 501370 371176
rect 501404 371142 501460 371176
rect 501494 371142 501550 371176
rect 501584 371142 501640 371176
rect 501674 371142 501730 371176
rect 501764 371142 501820 371176
rect 501854 371142 501908 371176
rect 501228 371086 501908 371142
rect 501228 371052 501280 371086
rect 501314 371052 501370 371086
rect 501404 371052 501460 371086
rect 501494 371052 501550 371086
rect 501584 371052 501640 371086
rect 501674 371052 501730 371086
rect 501764 371052 501820 371086
rect 501854 371052 501908 371086
rect 501228 370996 501908 371052
rect 501228 370962 501280 370996
rect 501314 370962 501370 370996
rect 501404 370962 501460 370996
rect 501494 370962 501550 370996
rect 501584 370962 501640 370996
rect 501674 370962 501730 370996
rect 501764 370962 501820 370996
rect 501854 370962 501908 370996
rect 501228 370906 501908 370962
rect 501228 370872 501280 370906
rect 501314 370872 501370 370906
rect 501404 370872 501460 370906
rect 501494 370872 501550 370906
rect 501584 370872 501640 370906
rect 501674 370872 501730 370906
rect 501764 370872 501820 370906
rect 501854 370872 501908 370906
rect 501228 370820 501908 370872
rect 501228 370106 501908 370160
rect 501228 370072 501280 370106
rect 501314 370072 501370 370106
rect 501404 370072 501460 370106
rect 501494 370072 501550 370106
rect 501584 370072 501640 370106
rect 501674 370072 501730 370106
rect 501764 370072 501820 370106
rect 501854 370072 501908 370106
rect 501228 370016 501908 370072
rect 501228 369982 501280 370016
rect 501314 369982 501370 370016
rect 501404 369982 501460 370016
rect 501494 369982 501550 370016
rect 501584 369982 501640 370016
rect 501674 369982 501730 370016
rect 501764 369982 501820 370016
rect 501854 369982 501908 370016
rect 501228 369926 501908 369982
rect 501228 369892 501280 369926
rect 501314 369892 501370 369926
rect 501404 369892 501460 369926
rect 501494 369892 501550 369926
rect 501584 369892 501640 369926
rect 501674 369892 501730 369926
rect 501764 369892 501820 369926
rect 501854 369892 501908 369926
rect 501228 369836 501908 369892
rect 501228 369802 501280 369836
rect 501314 369802 501370 369836
rect 501404 369802 501460 369836
rect 501494 369802 501550 369836
rect 501584 369802 501640 369836
rect 501674 369802 501730 369836
rect 501764 369802 501820 369836
rect 501854 369802 501908 369836
rect 501228 369746 501908 369802
rect 501228 369712 501280 369746
rect 501314 369712 501370 369746
rect 501404 369712 501460 369746
rect 501494 369712 501550 369746
rect 501584 369712 501640 369746
rect 501674 369712 501730 369746
rect 501764 369712 501820 369746
rect 501854 369712 501908 369746
rect 501228 369656 501908 369712
rect 501228 369622 501280 369656
rect 501314 369622 501370 369656
rect 501404 369622 501460 369656
rect 501494 369622 501550 369656
rect 501584 369622 501640 369656
rect 501674 369622 501730 369656
rect 501764 369622 501820 369656
rect 501854 369622 501908 369656
rect 501228 369566 501908 369622
rect 501228 369532 501280 369566
rect 501314 369532 501370 369566
rect 501404 369532 501460 369566
rect 501494 369532 501550 369566
rect 501584 369532 501640 369566
rect 501674 369532 501730 369566
rect 501764 369532 501820 369566
rect 501854 369532 501908 369566
rect 501228 369480 501908 369532
rect 501228 368766 501908 368820
rect 501228 368732 501280 368766
rect 501314 368732 501370 368766
rect 501404 368732 501460 368766
rect 501494 368732 501550 368766
rect 501584 368732 501640 368766
rect 501674 368732 501730 368766
rect 501764 368732 501820 368766
rect 501854 368732 501908 368766
rect 501228 368676 501908 368732
rect 501228 368642 501280 368676
rect 501314 368642 501370 368676
rect 501404 368642 501460 368676
rect 501494 368642 501550 368676
rect 501584 368642 501640 368676
rect 501674 368642 501730 368676
rect 501764 368642 501820 368676
rect 501854 368642 501908 368676
rect 501228 368586 501908 368642
rect 501228 368552 501280 368586
rect 501314 368552 501370 368586
rect 501404 368552 501460 368586
rect 501494 368552 501550 368586
rect 501584 368552 501640 368586
rect 501674 368552 501730 368586
rect 501764 368552 501820 368586
rect 501854 368552 501908 368586
rect 501228 368496 501908 368552
rect 501228 368462 501280 368496
rect 501314 368462 501370 368496
rect 501404 368462 501460 368496
rect 501494 368462 501550 368496
rect 501584 368462 501640 368496
rect 501674 368462 501730 368496
rect 501764 368462 501820 368496
rect 501854 368462 501908 368496
rect 501228 368406 501908 368462
rect 501228 368372 501280 368406
rect 501314 368372 501370 368406
rect 501404 368372 501460 368406
rect 501494 368372 501550 368406
rect 501584 368372 501640 368406
rect 501674 368372 501730 368406
rect 501764 368372 501820 368406
rect 501854 368372 501908 368406
rect 501228 368316 501908 368372
rect 501228 368282 501280 368316
rect 501314 368282 501370 368316
rect 501404 368282 501460 368316
rect 501494 368282 501550 368316
rect 501584 368282 501640 368316
rect 501674 368282 501730 368316
rect 501764 368282 501820 368316
rect 501854 368282 501908 368316
rect 501228 368226 501908 368282
rect 501228 368192 501280 368226
rect 501314 368192 501370 368226
rect 501404 368192 501460 368226
rect 501494 368192 501550 368226
rect 501584 368192 501640 368226
rect 501674 368192 501730 368226
rect 501764 368192 501820 368226
rect 501854 368192 501908 368226
rect 501228 368140 501908 368192
rect 501228 367426 501908 367480
rect 501228 367392 501280 367426
rect 501314 367392 501370 367426
rect 501404 367392 501460 367426
rect 501494 367392 501550 367426
rect 501584 367392 501640 367426
rect 501674 367392 501730 367426
rect 501764 367392 501820 367426
rect 501854 367392 501908 367426
rect 501228 367336 501908 367392
rect 501228 367302 501280 367336
rect 501314 367302 501370 367336
rect 501404 367302 501460 367336
rect 501494 367302 501550 367336
rect 501584 367302 501640 367336
rect 501674 367302 501730 367336
rect 501764 367302 501820 367336
rect 501854 367302 501908 367336
rect 501228 367246 501908 367302
rect 501228 367212 501280 367246
rect 501314 367212 501370 367246
rect 501404 367212 501460 367246
rect 501494 367212 501550 367246
rect 501584 367212 501640 367246
rect 501674 367212 501730 367246
rect 501764 367212 501820 367246
rect 501854 367212 501908 367246
rect 501228 367156 501908 367212
rect 501228 367122 501280 367156
rect 501314 367122 501370 367156
rect 501404 367122 501460 367156
rect 501494 367122 501550 367156
rect 501584 367122 501640 367156
rect 501674 367122 501730 367156
rect 501764 367122 501820 367156
rect 501854 367122 501908 367156
rect 501228 367066 501908 367122
rect 501228 367032 501280 367066
rect 501314 367032 501370 367066
rect 501404 367032 501460 367066
rect 501494 367032 501550 367066
rect 501584 367032 501640 367066
rect 501674 367032 501730 367066
rect 501764 367032 501820 367066
rect 501854 367032 501908 367066
rect 501228 366976 501908 367032
rect 501228 366942 501280 366976
rect 501314 366942 501370 366976
rect 501404 366942 501460 366976
rect 501494 366942 501550 366976
rect 501584 366942 501640 366976
rect 501674 366942 501730 366976
rect 501764 366942 501820 366976
rect 501854 366942 501908 366976
rect 501228 366886 501908 366942
rect 501228 366852 501280 366886
rect 501314 366852 501370 366886
rect 501404 366852 501460 366886
rect 501494 366852 501550 366886
rect 501584 366852 501640 366886
rect 501674 366852 501730 366886
rect 501764 366852 501820 366886
rect 501854 366852 501908 366886
rect 501228 366800 501908 366852
rect 501228 366086 501908 366140
rect 501228 366052 501280 366086
rect 501314 366052 501370 366086
rect 501404 366052 501460 366086
rect 501494 366052 501550 366086
rect 501584 366052 501640 366086
rect 501674 366052 501730 366086
rect 501764 366052 501820 366086
rect 501854 366052 501908 366086
rect 501228 365996 501908 366052
rect 501228 365962 501280 365996
rect 501314 365962 501370 365996
rect 501404 365962 501460 365996
rect 501494 365962 501550 365996
rect 501584 365962 501640 365996
rect 501674 365962 501730 365996
rect 501764 365962 501820 365996
rect 501854 365962 501908 365996
rect 501228 365906 501908 365962
rect 501228 365872 501280 365906
rect 501314 365872 501370 365906
rect 501404 365872 501460 365906
rect 501494 365872 501550 365906
rect 501584 365872 501640 365906
rect 501674 365872 501730 365906
rect 501764 365872 501820 365906
rect 501854 365872 501908 365906
rect 501228 365816 501908 365872
rect 501228 365782 501280 365816
rect 501314 365782 501370 365816
rect 501404 365782 501460 365816
rect 501494 365782 501550 365816
rect 501584 365782 501640 365816
rect 501674 365782 501730 365816
rect 501764 365782 501820 365816
rect 501854 365782 501908 365816
rect 501228 365726 501908 365782
rect 501228 365692 501280 365726
rect 501314 365692 501370 365726
rect 501404 365692 501460 365726
rect 501494 365692 501550 365726
rect 501584 365692 501640 365726
rect 501674 365692 501730 365726
rect 501764 365692 501820 365726
rect 501854 365692 501908 365726
rect 501228 365636 501908 365692
rect 501228 365602 501280 365636
rect 501314 365602 501370 365636
rect 501404 365602 501460 365636
rect 501494 365602 501550 365636
rect 501584 365602 501640 365636
rect 501674 365602 501730 365636
rect 501764 365602 501820 365636
rect 501854 365602 501908 365636
rect 501228 365546 501908 365602
rect 501228 365512 501280 365546
rect 501314 365512 501370 365546
rect 501404 365512 501460 365546
rect 501494 365512 501550 365546
rect 501584 365512 501640 365546
rect 501674 365512 501730 365546
rect 501764 365512 501820 365546
rect 501854 365512 501908 365546
rect 501228 365460 501908 365512
rect 501228 364746 501908 364800
rect 501228 364712 501280 364746
rect 501314 364712 501370 364746
rect 501404 364712 501460 364746
rect 501494 364712 501550 364746
rect 501584 364712 501640 364746
rect 501674 364712 501730 364746
rect 501764 364712 501820 364746
rect 501854 364712 501908 364746
rect 501228 364656 501908 364712
rect 501228 364622 501280 364656
rect 501314 364622 501370 364656
rect 501404 364622 501460 364656
rect 501494 364622 501550 364656
rect 501584 364622 501640 364656
rect 501674 364622 501730 364656
rect 501764 364622 501820 364656
rect 501854 364622 501908 364656
rect 501228 364566 501908 364622
rect 501228 364532 501280 364566
rect 501314 364532 501370 364566
rect 501404 364532 501460 364566
rect 501494 364532 501550 364566
rect 501584 364532 501640 364566
rect 501674 364532 501730 364566
rect 501764 364532 501820 364566
rect 501854 364532 501908 364566
rect 501228 364476 501908 364532
rect 501228 364442 501280 364476
rect 501314 364442 501370 364476
rect 501404 364442 501460 364476
rect 501494 364442 501550 364476
rect 501584 364442 501640 364476
rect 501674 364442 501730 364476
rect 501764 364442 501820 364476
rect 501854 364442 501908 364476
rect 501228 364386 501908 364442
rect 501228 364352 501280 364386
rect 501314 364352 501370 364386
rect 501404 364352 501460 364386
rect 501494 364352 501550 364386
rect 501584 364352 501640 364386
rect 501674 364352 501730 364386
rect 501764 364352 501820 364386
rect 501854 364352 501908 364386
rect 501228 364296 501908 364352
rect 501228 364262 501280 364296
rect 501314 364262 501370 364296
rect 501404 364262 501460 364296
rect 501494 364262 501550 364296
rect 501584 364262 501640 364296
rect 501674 364262 501730 364296
rect 501764 364262 501820 364296
rect 501854 364262 501908 364296
rect 501228 364206 501908 364262
rect 501228 364172 501280 364206
rect 501314 364172 501370 364206
rect 501404 364172 501460 364206
rect 501494 364172 501550 364206
rect 501584 364172 501640 364206
rect 501674 364172 501730 364206
rect 501764 364172 501820 364206
rect 501854 364172 501908 364206
rect 501228 364120 501908 364172
rect 501228 363406 501908 363460
rect 501228 363372 501280 363406
rect 501314 363372 501370 363406
rect 501404 363372 501460 363406
rect 501494 363372 501550 363406
rect 501584 363372 501640 363406
rect 501674 363372 501730 363406
rect 501764 363372 501820 363406
rect 501854 363372 501908 363406
rect 501228 363316 501908 363372
rect 501228 363282 501280 363316
rect 501314 363282 501370 363316
rect 501404 363282 501460 363316
rect 501494 363282 501550 363316
rect 501584 363282 501640 363316
rect 501674 363282 501730 363316
rect 501764 363282 501820 363316
rect 501854 363282 501908 363316
rect 501228 363226 501908 363282
rect 501228 363192 501280 363226
rect 501314 363192 501370 363226
rect 501404 363192 501460 363226
rect 501494 363192 501550 363226
rect 501584 363192 501640 363226
rect 501674 363192 501730 363226
rect 501764 363192 501820 363226
rect 501854 363192 501908 363226
rect 501228 363136 501908 363192
rect 501228 363102 501280 363136
rect 501314 363102 501370 363136
rect 501404 363102 501460 363136
rect 501494 363102 501550 363136
rect 501584 363102 501640 363136
rect 501674 363102 501730 363136
rect 501764 363102 501820 363136
rect 501854 363102 501908 363136
rect 501228 363046 501908 363102
rect 501228 363012 501280 363046
rect 501314 363012 501370 363046
rect 501404 363012 501460 363046
rect 501494 363012 501550 363046
rect 501584 363012 501640 363046
rect 501674 363012 501730 363046
rect 501764 363012 501820 363046
rect 501854 363012 501908 363046
rect 501228 362956 501908 363012
rect 501228 362922 501280 362956
rect 501314 362922 501370 362956
rect 501404 362922 501460 362956
rect 501494 362922 501550 362956
rect 501584 362922 501640 362956
rect 501674 362922 501730 362956
rect 501764 362922 501820 362956
rect 501854 362922 501908 362956
rect 501228 362866 501908 362922
rect 501228 362832 501280 362866
rect 501314 362832 501370 362866
rect 501404 362832 501460 362866
rect 501494 362832 501550 362866
rect 501584 362832 501640 362866
rect 501674 362832 501730 362866
rect 501764 362832 501820 362866
rect 501854 362832 501908 362866
rect 501228 362780 501908 362832
rect 504988 372786 505668 372840
rect 504988 372752 505040 372786
rect 505074 372752 505130 372786
rect 505164 372752 505220 372786
rect 505254 372752 505310 372786
rect 505344 372752 505400 372786
rect 505434 372752 505490 372786
rect 505524 372752 505580 372786
rect 505614 372752 505668 372786
rect 504988 372696 505668 372752
rect 504988 372662 505040 372696
rect 505074 372662 505130 372696
rect 505164 372662 505220 372696
rect 505254 372662 505310 372696
rect 505344 372662 505400 372696
rect 505434 372662 505490 372696
rect 505524 372662 505580 372696
rect 505614 372662 505668 372696
rect 504988 372606 505668 372662
rect 504988 372572 505040 372606
rect 505074 372572 505130 372606
rect 505164 372572 505220 372606
rect 505254 372572 505310 372606
rect 505344 372572 505400 372606
rect 505434 372572 505490 372606
rect 505524 372572 505580 372606
rect 505614 372572 505668 372606
rect 504988 372516 505668 372572
rect 504988 372482 505040 372516
rect 505074 372482 505130 372516
rect 505164 372482 505220 372516
rect 505254 372482 505310 372516
rect 505344 372482 505400 372516
rect 505434 372482 505490 372516
rect 505524 372482 505580 372516
rect 505614 372482 505668 372516
rect 504988 372426 505668 372482
rect 504988 372392 505040 372426
rect 505074 372392 505130 372426
rect 505164 372392 505220 372426
rect 505254 372392 505310 372426
rect 505344 372392 505400 372426
rect 505434 372392 505490 372426
rect 505524 372392 505580 372426
rect 505614 372392 505668 372426
rect 504988 372336 505668 372392
rect 504988 372302 505040 372336
rect 505074 372302 505130 372336
rect 505164 372302 505220 372336
rect 505254 372302 505310 372336
rect 505344 372302 505400 372336
rect 505434 372302 505490 372336
rect 505524 372302 505580 372336
rect 505614 372302 505668 372336
rect 504988 372246 505668 372302
rect 504988 372212 505040 372246
rect 505074 372212 505130 372246
rect 505164 372212 505220 372246
rect 505254 372212 505310 372246
rect 505344 372212 505400 372246
rect 505434 372212 505490 372246
rect 505524 372212 505580 372246
rect 505614 372212 505668 372246
rect 504988 372160 505668 372212
rect 504988 371446 505668 371500
rect 504988 371412 505040 371446
rect 505074 371412 505130 371446
rect 505164 371412 505220 371446
rect 505254 371412 505310 371446
rect 505344 371412 505400 371446
rect 505434 371412 505490 371446
rect 505524 371412 505580 371446
rect 505614 371412 505668 371446
rect 504988 371356 505668 371412
rect 504988 371322 505040 371356
rect 505074 371322 505130 371356
rect 505164 371322 505220 371356
rect 505254 371322 505310 371356
rect 505344 371322 505400 371356
rect 505434 371322 505490 371356
rect 505524 371322 505580 371356
rect 505614 371322 505668 371356
rect 504988 371266 505668 371322
rect 504988 371232 505040 371266
rect 505074 371232 505130 371266
rect 505164 371232 505220 371266
rect 505254 371232 505310 371266
rect 505344 371232 505400 371266
rect 505434 371232 505490 371266
rect 505524 371232 505580 371266
rect 505614 371232 505668 371266
rect 504988 371176 505668 371232
rect 504988 371142 505040 371176
rect 505074 371142 505130 371176
rect 505164 371142 505220 371176
rect 505254 371142 505310 371176
rect 505344 371142 505400 371176
rect 505434 371142 505490 371176
rect 505524 371142 505580 371176
rect 505614 371142 505668 371176
rect 504988 371086 505668 371142
rect 504988 371052 505040 371086
rect 505074 371052 505130 371086
rect 505164 371052 505220 371086
rect 505254 371052 505310 371086
rect 505344 371052 505400 371086
rect 505434 371052 505490 371086
rect 505524 371052 505580 371086
rect 505614 371052 505668 371086
rect 504988 370996 505668 371052
rect 504988 370962 505040 370996
rect 505074 370962 505130 370996
rect 505164 370962 505220 370996
rect 505254 370962 505310 370996
rect 505344 370962 505400 370996
rect 505434 370962 505490 370996
rect 505524 370962 505580 370996
rect 505614 370962 505668 370996
rect 504988 370906 505668 370962
rect 504988 370872 505040 370906
rect 505074 370872 505130 370906
rect 505164 370872 505220 370906
rect 505254 370872 505310 370906
rect 505344 370872 505400 370906
rect 505434 370872 505490 370906
rect 505524 370872 505580 370906
rect 505614 370872 505668 370906
rect 504988 370820 505668 370872
rect 504988 370106 505668 370160
rect 504988 370072 505040 370106
rect 505074 370072 505130 370106
rect 505164 370072 505220 370106
rect 505254 370072 505310 370106
rect 505344 370072 505400 370106
rect 505434 370072 505490 370106
rect 505524 370072 505580 370106
rect 505614 370072 505668 370106
rect 504988 370016 505668 370072
rect 504988 369982 505040 370016
rect 505074 369982 505130 370016
rect 505164 369982 505220 370016
rect 505254 369982 505310 370016
rect 505344 369982 505400 370016
rect 505434 369982 505490 370016
rect 505524 369982 505580 370016
rect 505614 369982 505668 370016
rect 504988 369926 505668 369982
rect 504988 369892 505040 369926
rect 505074 369892 505130 369926
rect 505164 369892 505220 369926
rect 505254 369892 505310 369926
rect 505344 369892 505400 369926
rect 505434 369892 505490 369926
rect 505524 369892 505580 369926
rect 505614 369892 505668 369926
rect 504988 369836 505668 369892
rect 504988 369802 505040 369836
rect 505074 369802 505130 369836
rect 505164 369802 505220 369836
rect 505254 369802 505310 369836
rect 505344 369802 505400 369836
rect 505434 369802 505490 369836
rect 505524 369802 505580 369836
rect 505614 369802 505668 369836
rect 504988 369746 505668 369802
rect 504988 369712 505040 369746
rect 505074 369712 505130 369746
rect 505164 369712 505220 369746
rect 505254 369712 505310 369746
rect 505344 369712 505400 369746
rect 505434 369712 505490 369746
rect 505524 369712 505580 369746
rect 505614 369712 505668 369746
rect 504988 369656 505668 369712
rect 504988 369622 505040 369656
rect 505074 369622 505130 369656
rect 505164 369622 505220 369656
rect 505254 369622 505310 369656
rect 505344 369622 505400 369656
rect 505434 369622 505490 369656
rect 505524 369622 505580 369656
rect 505614 369622 505668 369656
rect 504988 369566 505668 369622
rect 504988 369532 505040 369566
rect 505074 369532 505130 369566
rect 505164 369532 505220 369566
rect 505254 369532 505310 369566
rect 505344 369532 505400 369566
rect 505434 369532 505490 369566
rect 505524 369532 505580 369566
rect 505614 369532 505668 369566
rect 504988 369480 505668 369532
rect 504988 368766 505668 368820
rect 504988 368732 505040 368766
rect 505074 368732 505130 368766
rect 505164 368732 505220 368766
rect 505254 368732 505310 368766
rect 505344 368732 505400 368766
rect 505434 368732 505490 368766
rect 505524 368732 505580 368766
rect 505614 368732 505668 368766
rect 504988 368676 505668 368732
rect 504988 368642 505040 368676
rect 505074 368642 505130 368676
rect 505164 368642 505220 368676
rect 505254 368642 505310 368676
rect 505344 368642 505400 368676
rect 505434 368642 505490 368676
rect 505524 368642 505580 368676
rect 505614 368642 505668 368676
rect 504988 368586 505668 368642
rect 504988 368552 505040 368586
rect 505074 368552 505130 368586
rect 505164 368552 505220 368586
rect 505254 368552 505310 368586
rect 505344 368552 505400 368586
rect 505434 368552 505490 368586
rect 505524 368552 505580 368586
rect 505614 368552 505668 368586
rect 504988 368496 505668 368552
rect 504988 368462 505040 368496
rect 505074 368462 505130 368496
rect 505164 368462 505220 368496
rect 505254 368462 505310 368496
rect 505344 368462 505400 368496
rect 505434 368462 505490 368496
rect 505524 368462 505580 368496
rect 505614 368462 505668 368496
rect 504988 368406 505668 368462
rect 504988 368372 505040 368406
rect 505074 368372 505130 368406
rect 505164 368372 505220 368406
rect 505254 368372 505310 368406
rect 505344 368372 505400 368406
rect 505434 368372 505490 368406
rect 505524 368372 505580 368406
rect 505614 368372 505668 368406
rect 504988 368316 505668 368372
rect 504988 368282 505040 368316
rect 505074 368282 505130 368316
rect 505164 368282 505220 368316
rect 505254 368282 505310 368316
rect 505344 368282 505400 368316
rect 505434 368282 505490 368316
rect 505524 368282 505580 368316
rect 505614 368282 505668 368316
rect 504988 368226 505668 368282
rect 504988 368192 505040 368226
rect 505074 368192 505130 368226
rect 505164 368192 505220 368226
rect 505254 368192 505310 368226
rect 505344 368192 505400 368226
rect 505434 368192 505490 368226
rect 505524 368192 505580 368226
rect 505614 368192 505668 368226
rect 504988 368140 505668 368192
rect 504988 367426 505668 367480
rect 504988 367392 505040 367426
rect 505074 367392 505130 367426
rect 505164 367392 505220 367426
rect 505254 367392 505310 367426
rect 505344 367392 505400 367426
rect 505434 367392 505490 367426
rect 505524 367392 505580 367426
rect 505614 367392 505668 367426
rect 504988 367336 505668 367392
rect 504988 367302 505040 367336
rect 505074 367302 505130 367336
rect 505164 367302 505220 367336
rect 505254 367302 505310 367336
rect 505344 367302 505400 367336
rect 505434 367302 505490 367336
rect 505524 367302 505580 367336
rect 505614 367302 505668 367336
rect 504988 367246 505668 367302
rect 504988 367212 505040 367246
rect 505074 367212 505130 367246
rect 505164 367212 505220 367246
rect 505254 367212 505310 367246
rect 505344 367212 505400 367246
rect 505434 367212 505490 367246
rect 505524 367212 505580 367246
rect 505614 367212 505668 367246
rect 504988 367156 505668 367212
rect 504988 367122 505040 367156
rect 505074 367122 505130 367156
rect 505164 367122 505220 367156
rect 505254 367122 505310 367156
rect 505344 367122 505400 367156
rect 505434 367122 505490 367156
rect 505524 367122 505580 367156
rect 505614 367122 505668 367156
rect 504988 367066 505668 367122
rect 504988 367032 505040 367066
rect 505074 367032 505130 367066
rect 505164 367032 505220 367066
rect 505254 367032 505310 367066
rect 505344 367032 505400 367066
rect 505434 367032 505490 367066
rect 505524 367032 505580 367066
rect 505614 367032 505668 367066
rect 504988 366976 505668 367032
rect 504988 366942 505040 366976
rect 505074 366942 505130 366976
rect 505164 366942 505220 366976
rect 505254 366942 505310 366976
rect 505344 366942 505400 366976
rect 505434 366942 505490 366976
rect 505524 366942 505580 366976
rect 505614 366942 505668 366976
rect 504988 366886 505668 366942
rect 504988 366852 505040 366886
rect 505074 366852 505130 366886
rect 505164 366852 505220 366886
rect 505254 366852 505310 366886
rect 505344 366852 505400 366886
rect 505434 366852 505490 366886
rect 505524 366852 505580 366886
rect 505614 366852 505668 366886
rect 504988 366800 505668 366852
rect 504988 366086 505668 366140
rect 504988 366052 505040 366086
rect 505074 366052 505130 366086
rect 505164 366052 505220 366086
rect 505254 366052 505310 366086
rect 505344 366052 505400 366086
rect 505434 366052 505490 366086
rect 505524 366052 505580 366086
rect 505614 366052 505668 366086
rect 504988 365996 505668 366052
rect 504988 365962 505040 365996
rect 505074 365962 505130 365996
rect 505164 365962 505220 365996
rect 505254 365962 505310 365996
rect 505344 365962 505400 365996
rect 505434 365962 505490 365996
rect 505524 365962 505580 365996
rect 505614 365962 505668 365996
rect 504988 365906 505668 365962
rect 504988 365872 505040 365906
rect 505074 365872 505130 365906
rect 505164 365872 505220 365906
rect 505254 365872 505310 365906
rect 505344 365872 505400 365906
rect 505434 365872 505490 365906
rect 505524 365872 505580 365906
rect 505614 365872 505668 365906
rect 504988 365816 505668 365872
rect 504988 365782 505040 365816
rect 505074 365782 505130 365816
rect 505164 365782 505220 365816
rect 505254 365782 505310 365816
rect 505344 365782 505400 365816
rect 505434 365782 505490 365816
rect 505524 365782 505580 365816
rect 505614 365782 505668 365816
rect 504988 365726 505668 365782
rect 504988 365692 505040 365726
rect 505074 365692 505130 365726
rect 505164 365692 505220 365726
rect 505254 365692 505310 365726
rect 505344 365692 505400 365726
rect 505434 365692 505490 365726
rect 505524 365692 505580 365726
rect 505614 365692 505668 365726
rect 504988 365636 505668 365692
rect 504988 365602 505040 365636
rect 505074 365602 505130 365636
rect 505164 365602 505220 365636
rect 505254 365602 505310 365636
rect 505344 365602 505400 365636
rect 505434 365602 505490 365636
rect 505524 365602 505580 365636
rect 505614 365602 505668 365636
rect 504988 365546 505668 365602
rect 504988 365512 505040 365546
rect 505074 365512 505130 365546
rect 505164 365512 505220 365546
rect 505254 365512 505310 365546
rect 505344 365512 505400 365546
rect 505434 365512 505490 365546
rect 505524 365512 505580 365546
rect 505614 365512 505668 365546
rect 504988 365460 505668 365512
rect 504988 364746 505668 364800
rect 504988 364712 505040 364746
rect 505074 364712 505130 364746
rect 505164 364712 505220 364746
rect 505254 364712 505310 364746
rect 505344 364712 505400 364746
rect 505434 364712 505490 364746
rect 505524 364712 505580 364746
rect 505614 364712 505668 364746
rect 504988 364656 505668 364712
rect 504988 364622 505040 364656
rect 505074 364622 505130 364656
rect 505164 364622 505220 364656
rect 505254 364622 505310 364656
rect 505344 364622 505400 364656
rect 505434 364622 505490 364656
rect 505524 364622 505580 364656
rect 505614 364622 505668 364656
rect 504988 364566 505668 364622
rect 504988 364532 505040 364566
rect 505074 364532 505130 364566
rect 505164 364532 505220 364566
rect 505254 364532 505310 364566
rect 505344 364532 505400 364566
rect 505434 364532 505490 364566
rect 505524 364532 505580 364566
rect 505614 364532 505668 364566
rect 504988 364476 505668 364532
rect 504988 364442 505040 364476
rect 505074 364442 505130 364476
rect 505164 364442 505220 364476
rect 505254 364442 505310 364476
rect 505344 364442 505400 364476
rect 505434 364442 505490 364476
rect 505524 364442 505580 364476
rect 505614 364442 505668 364476
rect 504988 364386 505668 364442
rect 504988 364352 505040 364386
rect 505074 364352 505130 364386
rect 505164 364352 505220 364386
rect 505254 364352 505310 364386
rect 505344 364352 505400 364386
rect 505434 364352 505490 364386
rect 505524 364352 505580 364386
rect 505614 364352 505668 364386
rect 504988 364296 505668 364352
rect 504988 364262 505040 364296
rect 505074 364262 505130 364296
rect 505164 364262 505220 364296
rect 505254 364262 505310 364296
rect 505344 364262 505400 364296
rect 505434 364262 505490 364296
rect 505524 364262 505580 364296
rect 505614 364262 505668 364296
rect 504988 364206 505668 364262
rect 504988 364172 505040 364206
rect 505074 364172 505130 364206
rect 505164 364172 505220 364206
rect 505254 364172 505310 364206
rect 505344 364172 505400 364206
rect 505434 364172 505490 364206
rect 505524 364172 505580 364206
rect 505614 364172 505668 364206
rect 504988 364120 505668 364172
rect 504988 363406 505668 363460
rect 504988 363372 505040 363406
rect 505074 363372 505130 363406
rect 505164 363372 505220 363406
rect 505254 363372 505310 363406
rect 505344 363372 505400 363406
rect 505434 363372 505490 363406
rect 505524 363372 505580 363406
rect 505614 363372 505668 363406
rect 504988 363316 505668 363372
rect 504988 363282 505040 363316
rect 505074 363282 505130 363316
rect 505164 363282 505220 363316
rect 505254 363282 505310 363316
rect 505344 363282 505400 363316
rect 505434 363282 505490 363316
rect 505524 363282 505580 363316
rect 505614 363282 505668 363316
rect 504988 363226 505668 363282
rect 504988 363192 505040 363226
rect 505074 363192 505130 363226
rect 505164 363192 505220 363226
rect 505254 363192 505310 363226
rect 505344 363192 505400 363226
rect 505434 363192 505490 363226
rect 505524 363192 505580 363226
rect 505614 363192 505668 363226
rect 504988 363136 505668 363192
rect 504988 363102 505040 363136
rect 505074 363102 505130 363136
rect 505164 363102 505220 363136
rect 505254 363102 505310 363136
rect 505344 363102 505400 363136
rect 505434 363102 505490 363136
rect 505524 363102 505580 363136
rect 505614 363102 505668 363136
rect 504988 363046 505668 363102
rect 504988 363012 505040 363046
rect 505074 363012 505130 363046
rect 505164 363012 505220 363046
rect 505254 363012 505310 363046
rect 505344 363012 505400 363046
rect 505434 363012 505490 363046
rect 505524 363012 505580 363046
rect 505614 363012 505668 363046
rect 504988 362956 505668 363012
rect 504988 362922 505040 362956
rect 505074 362922 505130 362956
rect 505164 362922 505220 362956
rect 505254 362922 505310 362956
rect 505344 362922 505400 362956
rect 505434 362922 505490 362956
rect 505524 362922 505580 362956
rect 505614 362922 505668 362956
rect 504988 362866 505668 362922
rect 504988 362832 505040 362866
rect 505074 362832 505130 362866
rect 505164 362832 505220 362866
rect 505254 362832 505310 362866
rect 505344 362832 505400 362866
rect 505434 362832 505490 362866
rect 505524 362832 505580 362866
rect 505614 362832 505668 362866
rect 504988 362780 505668 362832
rect 508748 372786 509428 372840
rect 508748 372752 508800 372786
rect 508834 372752 508890 372786
rect 508924 372752 508980 372786
rect 509014 372752 509070 372786
rect 509104 372752 509160 372786
rect 509194 372752 509250 372786
rect 509284 372752 509340 372786
rect 509374 372752 509428 372786
rect 508748 372696 509428 372752
rect 508748 372662 508800 372696
rect 508834 372662 508890 372696
rect 508924 372662 508980 372696
rect 509014 372662 509070 372696
rect 509104 372662 509160 372696
rect 509194 372662 509250 372696
rect 509284 372662 509340 372696
rect 509374 372662 509428 372696
rect 508748 372606 509428 372662
rect 508748 372572 508800 372606
rect 508834 372572 508890 372606
rect 508924 372572 508980 372606
rect 509014 372572 509070 372606
rect 509104 372572 509160 372606
rect 509194 372572 509250 372606
rect 509284 372572 509340 372606
rect 509374 372572 509428 372606
rect 508748 372516 509428 372572
rect 508748 372482 508800 372516
rect 508834 372482 508890 372516
rect 508924 372482 508980 372516
rect 509014 372482 509070 372516
rect 509104 372482 509160 372516
rect 509194 372482 509250 372516
rect 509284 372482 509340 372516
rect 509374 372482 509428 372516
rect 508748 372426 509428 372482
rect 508748 372392 508800 372426
rect 508834 372392 508890 372426
rect 508924 372392 508980 372426
rect 509014 372392 509070 372426
rect 509104 372392 509160 372426
rect 509194 372392 509250 372426
rect 509284 372392 509340 372426
rect 509374 372392 509428 372426
rect 508748 372336 509428 372392
rect 508748 372302 508800 372336
rect 508834 372302 508890 372336
rect 508924 372302 508980 372336
rect 509014 372302 509070 372336
rect 509104 372302 509160 372336
rect 509194 372302 509250 372336
rect 509284 372302 509340 372336
rect 509374 372302 509428 372336
rect 508748 372246 509428 372302
rect 508748 372212 508800 372246
rect 508834 372212 508890 372246
rect 508924 372212 508980 372246
rect 509014 372212 509070 372246
rect 509104 372212 509160 372246
rect 509194 372212 509250 372246
rect 509284 372212 509340 372246
rect 509374 372212 509428 372246
rect 508748 372160 509428 372212
rect 508748 371446 509428 371500
rect 508748 371412 508800 371446
rect 508834 371412 508890 371446
rect 508924 371412 508980 371446
rect 509014 371412 509070 371446
rect 509104 371412 509160 371446
rect 509194 371412 509250 371446
rect 509284 371412 509340 371446
rect 509374 371412 509428 371446
rect 508748 371356 509428 371412
rect 508748 371322 508800 371356
rect 508834 371322 508890 371356
rect 508924 371322 508980 371356
rect 509014 371322 509070 371356
rect 509104 371322 509160 371356
rect 509194 371322 509250 371356
rect 509284 371322 509340 371356
rect 509374 371322 509428 371356
rect 508748 371266 509428 371322
rect 508748 371232 508800 371266
rect 508834 371232 508890 371266
rect 508924 371232 508980 371266
rect 509014 371232 509070 371266
rect 509104 371232 509160 371266
rect 509194 371232 509250 371266
rect 509284 371232 509340 371266
rect 509374 371232 509428 371266
rect 508748 371176 509428 371232
rect 508748 371142 508800 371176
rect 508834 371142 508890 371176
rect 508924 371142 508980 371176
rect 509014 371142 509070 371176
rect 509104 371142 509160 371176
rect 509194 371142 509250 371176
rect 509284 371142 509340 371176
rect 509374 371142 509428 371176
rect 508748 371086 509428 371142
rect 508748 371052 508800 371086
rect 508834 371052 508890 371086
rect 508924 371052 508980 371086
rect 509014 371052 509070 371086
rect 509104 371052 509160 371086
rect 509194 371052 509250 371086
rect 509284 371052 509340 371086
rect 509374 371052 509428 371086
rect 508748 370996 509428 371052
rect 508748 370962 508800 370996
rect 508834 370962 508890 370996
rect 508924 370962 508980 370996
rect 509014 370962 509070 370996
rect 509104 370962 509160 370996
rect 509194 370962 509250 370996
rect 509284 370962 509340 370996
rect 509374 370962 509428 370996
rect 508748 370906 509428 370962
rect 508748 370872 508800 370906
rect 508834 370872 508890 370906
rect 508924 370872 508980 370906
rect 509014 370872 509070 370906
rect 509104 370872 509160 370906
rect 509194 370872 509250 370906
rect 509284 370872 509340 370906
rect 509374 370872 509428 370906
rect 508748 370820 509428 370872
rect 508748 370106 509428 370160
rect 508748 370072 508800 370106
rect 508834 370072 508890 370106
rect 508924 370072 508980 370106
rect 509014 370072 509070 370106
rect 509104 370072 509160 370106
rect 509194 370072 509250 370106
rect 509284 370072 509340 370106
rect 509374 370072 509428 370106
rect 508748 370016 509428 370072
rect 508748 369982 508800 370016
rect 508834 369982 508890 370016
rect 508924 369982 508980 370016
rect 509014 369982 509070 370016
rect 509104 369982 509160 370016
rect 509194 369982 509250 370016
rect 509284 369982 509340 370016
rect 509374 369982 509428 370016
rect 508748 369926 509428 369982
rect 508748 369892 508800 369926
rect 508834 369892 508890 369926
rect 508924 369892 508980 369926
rect 509014 369892 509070 369926
rect 509104 369892 509160 369926
rect 509194 369892 509250 369926
rect 509284 369892 509340 369926
rect 509374 369892 509428 369926
rect 508748 369836 509428 369892
rect 508748 369802 508800 369836
rect 508834 369802 508890 369836
rect 508924 369802 508980 369836
rect 509014 369802 509070 369836
rect 509104 369802 509160 369836
rect 509194 369802 509250 369836
rect 509284 369802 509340 369836
rect 509374 369802 509428 369836
rect 508748 369746 509428 369802
rect 508748 369712 508800 369746
rect 508834 369712 508890 369746
rect 508924 369712 508980 369746
rect 509014 369712 509070 369746
rect 509104 369712 509160 369746
rect 509194 369712 509250 369746
rect 509284 369712 509340 369746
rect 509374 369712 509428 369746
rect 508748 369656 509428 369712
rect 508748 369622 508800 369656
rect 508834 369622 508890 369656
rect 508924 369622 508980 369656
rect 509014 369622 509070 369656
rect 509104 369622 509160 369656
rect 509194 369622 509250 369656
rect 509284 369622 509340 369656
rect 509374 369622 509428 369656
rect 508748 369566 509428 369622
rect 508748 369532 508800 369566
rect 508834 369532 508890 369566
rect 508924 369532 508980 369566
rect 509014 369532 509070 369566
rect 509104 369532 509160 369566
rect 509194 369532 509250 369566
rect 509284 369532 509340 369566
rect 509374 369532 509428 369566
rect 508748 369480 509428 369532
rect 508748 368766 509428 368820
rect 508748 368732 508800 368766
rect 508834 368732 508890 368766
rect 508924 368732 508980 368766
rect 509014 368732 509070 368766
rect 509104 368732 509160 368766
rect 509194 368732 509250 368766
rect 509284 368732 509340 368766
rect 509374 368732 509428 368766
rect 508748 368676 509428 368732
rect 508748 368642 508800 368676
rect 508834 368642 508890 368676
rect 508924 368642 508980 368676
rect 509014 368642 509070 368676
rect 509104 368642 509160 368676
rect 509194 368642 509250 368676
rect 509284 368642 509340 368676
rect 509374 368642 509428 368676
rect 508748 368586 509428 368642
rect 508748 368552 508800 368586
rect 508834 368552 508890 368586
rect 508924 368552 508980 368586
rect 509014 368552 509070 368586
rect 509104 368552 509160 368586
rect 509194 368552 509250 368586
rect 509284 368552 509340 368586
rect 509374 368552 509428 368586
rect 508748 368496 509428 368552
rect 508748 368462 508800 368496
rect 508834 368462 508890 368496
rect 508924 368462 508980 368496
rect 509014 368462 509070 368496
rect 509104 368462 509160 368496
rect 509194 368462 509250 368496
rect 509284 368462 509340 368496
rect 509374 368462 509428 368496
rect 508748 368406 509428 368462
rect 508748 368372 508800 368406
rect 508834 368372 508890 368406
rect 508924 368372 508980 368406
rect 509014 368372 509070 368406
rect 509104 368372 509160 368406
rect 509194 368372 509250 368406
rect 509284 368372 509340 368406
rect 509374 368372 509428 368406
rect 508748 368316 509428 368372
rect 508748 368282 508800 368316
rect 508834 368282 508890 368316
rect 508924 368282 508980 368316
rect 509014 368282 509070 368316
rect 509104 368282 509160 368316
rect 509194 368282 509250 368316
rect 509284 368282 509340 368316
rect 509374 368282 509428 368316
rect 508748 368226 509428 368282
rect 508748 368192 508800 368226
rect 508834 368192 508890 368226
rect 508924 368192 508980 368226
rect 509014 368192 509070 368226
rect 509104 368192 509160 368226
rect 509194 368192 509250 368226
rect 509284 368192 509340 368226
rect 509374 368192 509428 368226
rect 508748 368140 509428 368192
rect 508748 367426 509428 367480
rect 508748 367392 508800 367426
rect 508834 367392 508890 367426
rect 508924 367392 508980 367426
rect 509014 367392 509070 367426
rect 509104 367392 509160 367426
rect 509194 367392 509250 367426
rect 509284 367392 509340 367426
rect 509374 367392 509428 367426
rect 508748 367336 509428 367392
rect 508748 367302 508800 367336
rect 508834 367302 508890 367336
rect 508924 367302 508980 367336
rect 509014 367302 509070 367336
rect 509104 367302 509160 367336
rect 509194 367302 509250 367336
rect 509284 367302 509340 367336
rect 509374 367302 509428 367336
rect 508748 367246 509428 367302
rect 508748 367212 508800 367246
rect 508834 367212 508890 367246
rect 508924 367212 508980 367246
rect 509014 367212 509070 367246
rect 509104 367212 509160 367246
rect 509194 367212 509250 367246
rect 509284 367212 509340 367246
rect 509374 367212 509428 367246
rect 508748 367156 509428 367212
rect 508748 367122 508800 367156
rect 508834 367122 508890 367156
rect 508924 367122 508980 367156
rect 509014 367122 509070 367156
rect 509104 367122 509160 367156
rect 509194 367122 509250 367156
rect 509284 367122 509340 367156
rect 509374 367122 509428 367156
rect 508748 367066 509428 367122
rect 508748 367032 508800 367066
rect 508834 367032 508890 367066
rect 508924 367032 508980 367066
rect 509014 367032 509070 367066
rect 509104 367032 509160 367066
rect 509194 367032 509250 367066
rect 509284 367032 509340 367066
rect 509374 367032 509428 367066
rect 508748 366976 509428 367032
rect 508748 366942 508800 366976
rect 508834 366942 508890 366976
rect 508924 366942 508980 366976
rect 509014 366942 509070 366976
rect 509104 366942 509160 366976
rect 509194 366942 509250 366976
rect 509284 366942 509340 366976
rect 509374 366942 509428 366976
rect 508748 366886 509428 366942
rect 508748 366852 508800 366886
rect 508834 366852 508890 366886
rect 508924 366852 508980 366886
rect 509014 366852 509070 366886
rect 509104 366852 509160 366886
rect 509194 366852 509250 366886
rect 509284 366852 509340 366886
rect 509374 366852 509428 366886
rect 508748 366800 509428 366852
rect 508748 366086 509428 366140
rect 508748 366052 508800 366086
rect 508834 366052 508890 366086
rect 508924 366052 508980 366086
rect 509014 366052 509070 366086
rect 509104 366052 509160 366086
rect 509194 366052 509250 366086
rect 509284 366052 509340 366086
rect 509374 366052 509428 366086
rect 508748 365996 509428 366052
rect 508748 365962 508800 365996
rect 508834 365962 508890 365996
rect 508924 365962 508980 365996
rect 509014 365962 509070 365996
rect 509104 365962 509160 365996
rect 509194 365962 509250 365996
rect 509284 365962 509340 365996
rect 509374 365962 509428 365996
rect 508748 365906 509428 365962
rect 508748 365872 508800 365906
rect 508834 365872 508890 365906
rect 508924 365872 508980 365906
rect 509014 365872 509070 365906
rect 509104 365872 509160 365906
rect 509194 365872 509250 365906
rect 509284 365872 509340 365906
rect 509374 365872 509428 365906
rect 508748 365816 509428 365872
rect 508748 365782 508800 365816
rect 508834 365782 508890 365816
rect 508924 365782 508980 365816
rect 509014 365782 509070 365816
rect 509104 365782 509160 365816
rect 509194 365782 509250 365816
rect 509284 365782 509340 365816
rect 509374 365782 509428 365816
rect 508748 365726 509428 365782
rect 508748 365692 508800 365726
rect 508834 365692 508890 365726
rect 508924 365692 508980 365726
rect 509014 365692 509070 365726
rect 509104 365692 509160 365726
rect 509194 365692 509250 365726
rect 509284 365692 509340 365726
rect 509374 365692 509428 365726
rect 508748 365636 509428 365692
rect 508748 365602 508800 365636
rect 508834 365602 508890 365636
rect 508924 365602 508980 365636
rect 509014 365602 509070 365636
rect 509104 365602 509160 365636
rect 509194 365602 509250 365636
rect 509284 365602 509340 365636
rect 509374 365602 509428 365636
rect 508748 365546 509428 365602
rect 508748 365512 508800 365546
rect 508834 365512 508890 365546
rect 508924 365512 508980 365546
rect 509014 365512 509070 365546
rect 509104 365512 509160 365546
rect 509194 365512 509250 365546
rect 509284 365512 509340 365546
rect 509374 365512 509428 365546
rect 508748 365460 509428 365512
rect 508748 364746 509428 364800
rect 508748 364712 508800 364746
rect 508834 364712 508890 364746
rect 508924 364712 508980 364746
rect 509014 364712 509070 364746
rect 509104 364712 509160 364746
rect 509194 364712 509250 364746
rect 509284 364712 509340 364746
rect 509374 364712 509428 364746
rect 508748 364656 509428 364712
rect 508748 364622 508800 364656
rect 508834 364622 508890 364656
rect 508924 364622 508980 364656
rect 509014 364622 509070 364656
rect 509104 364622 509160 364656
rect 509194 364622 509250 364656
rect 509284 364622 509340 364656
rect 509374 364622 509428 364656
rect 508748 364566 509428 364622
rect 508748 364532 508800 364566
rect 508834 364532 508890 364566
rect 508924 364532 508980 364566
rect 509014 364532 509070 364566
rect 509104 364532 509160 364566
rect 509194 364532 509250 364566
rect 509284 364532 509340 364566
rect 509374 364532 509428 364566
rect 508748 364476 509428 364532
rect 508748 364442 508800 364476
rect 508834 364442 508890 364476
rect 508924 364442 508980 364476
rect 509014 364442 509070 364476
rect 509104 364442 509160 364476
rect 509194 364442 509250 364476
rect 509284 364442 509340 364476
rect 509374 364442 509428 364476
rect 508748 364386 509428 364442
rect 508748 364352 508800 364386
rect 508834 364352 508890 364386
rect 508924 364352 508980 364386
rect 509014 364352 509070 364386
rect 509104 364352 509160 364386
rect 509194 364352 509250 364386
rect 509284 364352 509340 364386
rect 509374 364352 509428 364386
rect 508748 364296 509428 364352
rect 508748 364262 508800 364296
rect 508834 364262 508890 364296
rect 508924 364262 508980 364296
rect 509014 364262 509070 364296
rect 509104 364262 509160 364296
rect 509194 364262 509250 364296
rect 509284 364262 509340 364296
rect 509374 364262 509428 364296
rect 508748 364206 509428 364262
rect 508748 364172 508800 364206
rect 508834 364172 508890 364206
rect 508924 364172 508980 364206
rect 509014 364172 509070 364206
rect 509104 364172 509160 364206
rect 509194 364172 509250 364206
rect 509284 364172 509340 364206
rect 509374 364172 509428 364206
rect 508748 364120 509428 364172
rect 508748 363406 509428 363460
rect 508748 363372 508800 363406
rect 508834 363372 508890 363406
rect 508924 363372 508980 363406
rect 509014 363372 509070 363406
rect 509104 363372 509160 363406
rect 509194 363372 509250 363406
rect 509284 363372 509340 363406
rect 509374 363372 509428 363406
rect 508748 363316 509428 363372
rect 508748 363282 508800 363316
rect 508834 363282 508890 363316
rect 508924 363282 508980 363316
rect 509014 363282 509070 363316
rect 509104 363282 509160 363316
rect 509194 363282 509250 363316
rect 509284 363282 509340 363316
rect 509374 363282 509428 363316
rect 508748 363226 509428 363282
rect 508748 363192 508800 363226
rect 508834 363192 508890 363226
rect 508924 363192 508980 363226
rect 509014 363192 509070 363226
rect 509104 363192 509160 363226
rect 509194 363192 509250 363226
rect 509284 363192 509340 363226
rect 509374 363192 509428 363226
rect 508748 363136 509428 363192
rect 508748 363102 508800 363136
rect 508834 363102 508890 363136
rect 508924 363102 508980 363136
rect 509014 363102 509070 363136
rect 509104 363102 509160 363136
rect 509194 363102 509250 363136
rect 509284 363102 509340 363136
rect 509374 363102 509428 363136
rect 508748 363046 509428 363102
rect 508748 363012 508800 363046
rect 508834 363012 508890 363046
rect 508924 363012 508980 363046
rect 509014 363012 509070 363046
rect 509104 363012 509160 363046
rect 509194 363012 509250 363046
rect 509284 363012 509340 363046
rect 509374 363012 509428 363046
rect 508748 362956 509428 363012
rect 508748 362922 508800 362956
rect 508834 362922 508890 362956
rect 508924 362922 508980 362956
rect 509014 362922 509070 362956
rect 509104 362922 509160 362956
rect 509194 362922 509250 362956
rect 509284 362922 509340 362956
rect 509374 362922 509428 362956
rect 508748 362866 509428 362922
rect 508748 362832 508800 362866
rect 508834 362832 508890 362866
rect 508924 362832 508980 362866
rect 509014 362832 509070 362866
rect 509104 362832 509160 362866
rect 509194 362832 509250 362866
rect 509284 362832 509340 362866
rect 509374 362832 509428 362866
rect 508748 362780 509428 362832
rect 512508 372786 513188 372840
rect 512508 372752 512560 372786
rect 512594 372752 512650 372786
rect 512684 372752 512740 372786
rect 512774 372752 512830 372786
rect 512864 372752 512920 372786
rect 512954 372752 513010 372786
rect 513044 372752 513100 372786
rect 513134 372752 513188 372786
rect 512508 372696 513188 372752
rect 512508 372662 512560 372696
rect 512594 372662 512650 372696
rect 512684 372662 512740 372696
rect 512774 372662 512830 372696
rect 512864 372662 512920 372696
rect 512954 372662 513010 372696
rect 513044 372662 513100 372696
rect 513134 372662 513188 372696
rect 512508 372606 513188 372662
rect 512508 372572 512560 372606
rect 512594 372572 512650 372606
rect 512684 372572 512740 372606
rect 512774 372572 512830 372606
rect 512864 372572 512920 372606
rect 512954 372572 513010 372606
rect 513044 372572 513100 372606
rect 513134 372572 513188 372606
rect 512508 372516 513188 372572
rect 512508 372482 512560 372516
rect 512594 372482 512650 372516
rect 512684 372482 512740 372516
rect 512774 372482 512830 372516
rect 512864 372482 512920 372516
rect 512954 372482 513010 372516
rect 513044 372482 513100 372516
rect 513134 372482 513188 372516
rect 512508 372426 513188 372482
rect 512508 372392 512560 372426
rect 512594 372392 512650 372426
rect 512684 372392 512740 372426
rect 512774 372392 512830 372426
rect 512864 372392 512920 372426
rect 512954 372392 513010 372426
rect 513044 372392 513100 372426
rect 513134 372392 513188 372426
rect 512508 372336 513188 372392
rect 512508 372302 512560 372336
rect 512594 372302 512650 372336
rect 512684 372302 512740 372336
rect 512774 372302 512830 372336
rect 512864 372302 512920 372336
rect 512954 372302 513010 372336
rect 513044 372302 513100 372336
rect 513134 372302 513188 372336
rect 512508 372246 513188 372302
rect 512508 372212 512560 372246
rect 512594 372212 512650 372246
rect 512684 372212 512740 372246
rect 512774 372212 512830 372246
rect 512864 372212 512920 372246
rect 512954 372212 513010 372246
rect 513044 372212 513100 372246
rect 513134 372212 513188 372246
rect 512508 372160 513188 372212
rect 523423 374505 524713 374517
rect 523423 374471 523439 374505
rect 523473 374471 523507 374505
rect 523541 374471 523575 374505
rect 523609 374471 523643 374505
rect 523677 374471 523711 374505
rect 523745 374471 523779 374505
rect 523813 374471 523847 374505
rect 523881 374471 523915 374505
rect 523949 374471 523983 374505
rect 524017 374471 524051 374505
rect 524085 374471 524119 374505
rect 524153 374471 524187 374505
rect 524221 374471 524255 374505
rect 524289 374471 524323 374505
rect 524357 374471 524391 374505
rect 524425 374471 524459 374505
rect 524493 374471 524527 374505
rect 524561 374471 524595 374505
rect 524629 374471 524663 374505
rect 524697 374471 524713 374505
rect 523423 374459 524713 374471
rect 523423 374047 524713 374059
rect 523423 374013 523439 374047
rect 523473 374013 523507 374047
rect 523541 374013 523575 374047
rect 523609 374013 523643 374047
rect 523677 374013 523711 374047
rect 523745 374013 523779 374047
rect 523813 374013 523847 374047
rect 523881 374013 523915 374047
rect 523949 374013 523983 374047
rect 524017 374013 524051 374047
rect 524085 374013 524119 374047
rect 524153 374013 524187 374047
rect 524221 374013 524255 374047
rect 524289 374013 524323 374047
rect 524357 374013 524391 374047
rect 524425 374013 524459 374047
rect 524493 374013 524527 374047
rect 524561 374013 524595 374047
rect 524629 374013 524663 374047
rect 524697 374013 524713 374047
rect 523423 374001 524713 374013
rect 523423 373589 524713 373601
rect 523423 373555 523439 373589
rect 523473 373555 523507 373589
rect 523541 373555 523575 373589
rect 523609 373555 523643 373589
rect 523677 373555 523711 373589
rect 523745 373555 523779 373589
rect 523813 373555 523847 373589
rect 523881 373555 523915 373589
rect 523949 373555 523983 373589
rect 524017 373555 524051 373589
rect 524085 373555 524119 373589
rect 524153 373555 524187 373589
rect 524221 373555 524255 373589
rect 524289 373555 524323 373589
rect 524357 373555 524391 373589
rect 524425 373555 524459 373589
rect 524493 373555 524527 373589
rect 524561 373555 524595 373589
rect 524629 373555 524663 373589
rect 524697 373555 524713 373589
rect 523423 373543 524713 373555
rect 523423 373131 524713 373143
rect 523423 373097 523439 373131
rect 523473 373097 523507 373131
rect 523541 373097 523575 373131
rect 523609 373097 523643 373131
rect 523677 373097 523711 373131
rect 523745 373097 523779 373131
rect 523813 373097 523847 373131
rect 523881 373097 523915 373131
rect 523949 373097 523983 373131
rect 524017 373097 524051 373131
rect 524085 373097 524119 373131
rect 524153 373097 524187 373131
rect 524221 373097 524255 373131
rect 524289 373097 524323 373131
rect 524357 373097 524391 373131
rect 524425 373097 524459 373131
rect 524493 373097 524527 373131
rect 524561 373097 524595 373131
rect 524629 373097 524663 373131
rect 524697 373097 524713 373131
rect 523423 373085 524713 373097
rect 523423 372673 524713 372685
rect 523423 372639 523439 372673
rect 523473 372639 523507 372673
rect 523541 372639 523575 372673
rect 523609 372639 523643 372673
rect 523677 372639 523711 372673
rect 523745 372639 523779 372673
rect 523813 372639 523847 372673
rect 523881 372639 523915 372673
rect 523949 372639 523983 372673
rect 524017 372639 524051 372673
rect 524085 372639 524119 372673
rect 524153 372639 524187 372673
rect 524221 372639 524255 372673
rect 524289 372639 524323 372673
rect 524357 372639 524391 372673
rect 524425 372639 524459 372673
rect 524493 372639 524527 372673
rect 524561 372639 524595 372673
rect 524629 372639 524663 372673
rect 524697 372639 524713 372673
rect 523423 372627 524713 372639
rect 523423 372215 524713 372227
rect 523423 372181 523439 372215
rect 523473 372181 523507 372215
rect 523541 372181 523575 372215
rect 523609 372181 523643 372215
rect 523677 372181 523711 372215
rect 523745 372181 523779 372215
rect 523813 372181 523847 372215
rect 523881 372181 523915 372215
rect 523949 372181 523983 372215
rect 524017 372181 524051 372215
rect 524085 372181 524119 372215
rect 524153 372181 524187 372215
rect 524221 372181 524255 372215
rect 524289 372181 524323 372215
rect 524357 372181 524391 372215
rect 524425 372181 524459 372215
rect 524493 372181 524527 372215
rect 524561 372181 524595 372215
rect 524629 372181 524663 372215
rect 524697 372181 524713 372215
rect 523423 372169 524713 372181
rect 512508 371446 513188 371500
rect 512508 371412 512560 371446
rect 512594 371412 512650 371446
rect 512684 371412 512740 371446
rect 512774 371412 512830 371446
rect 512864 371412 512920 371446
rect 512954 371412 513010 371446
rect 513044 371412 513100 371446
rect 513134 371412 513188 371446
rect 512508 371356 513188 371412
rect 512508 371322 512560 371356
rect 512594 371322 512650 371356
rect 512684 371322 512740 371356
rect 512774 371322 512830 371356
rect 512864 371322 512920 371356
rect 512954 371322 513010 371356
rect 513044 371322 513100 371356
rect 513134 371322 513188 371356
rect 512508 371266 513188 371322
rect 512508 371232 512560 371266
rect 512594 371232 512650 371266
rect 512684 371232 512740 371266
rect 512774 371232 512830 371266
rect 512864 371232 512920 371266
rect 512954 371232 513010 371266
rect 513044 371232 513100 371266
rect 513134 371232 513188 371266
rect 512508 371176 513188 371232
rect 512508 371142 512560 371176
rect 512594 371142 512650 371176
rect 512684 371142 512740 371176
rect 512774 371142 512830 371176
rect 512864 371142 512920 371176
rect 512954 371142 513010 371176
rect 513044 371142 513100 371176
rect 513134 371142 513188 371176
rect 512508 371086 513188 371142
rect 512508 371052 512560 371086
rect 512594 371052 512650 371086
rect 512684 371052 512740 371086
rect 512774 371052 512830 371086
rect 512864 371052 512920 371086
rect 512954 371052 513010 371086
rect 513044 371052 513100 371086
rect 513134 371052 513188 371086
rect 512508 370996 513188 371052
rect 512508 370962 512560 370996
rect 512594 370962 512650 370996
rect 512684 370962 512740 370996
rect 512774 370962 512830 370996
rect 512864 370962 512920 370996
rect 512954 370962 513010 370996
rect 513044 370962 513100 370996
rect 513134 370962 513188 370996
rect 512508 370906 513188 370962
rect 512508 370872 512560 370906
rect 512594 370872 512650 370906
rect 512684 370872 512740 370906
rect 512774 370872 512830 370906
rect 512864 370872 512920 370906
rect 512954 370872 513010 370906
rect 513044 370872 513100 370906
rect 513134 370872 513188 370906
rect 512508 370820 513188 370872
rect 512508 370106 513188 370160
rect 512508 370072 512560 370106
rect 512594 370072 512650 370106
rect 512684 370072 512740 370106
rect 512774 370072 512830 370106
rect 512864 370072 512920 370106
rect 512954 370072 513010 370106
rect 513044 370072 513100 370106
rect 513134 370072 513188 370106
rect 512508 370016 513188 370072
rect 512508 369982 512560 370016
rect 512594 369982 512650 370016
rect 512684 369982 512740 370016
rect 512774 369982 512830 370016
rect 512864 369982 512920 370016
rect 512954 369982 513010 370016
rect 513044 369982 513100 370016
rect 513134 369982 513188 370016
rect 512508 369926 513188 369982
rect 512508 369892 512560 369926
rect 512594 369892 512650 369926
rect 512684 369892 512740 369926
rect 512774 369892 512830 369926
rect 512864 369892 512920 369926
rect 512954 369892 513010 369926
rect 513044 369892 513100 369926
rect 513134 369892 513188 369926
rect 512508 369836 513188 369892
rect 512508 369802 512560 369836
rect 512594 369802 512650 369836
rect 512684 369802 512740 369836
rect 512774 369802 512830 369836
rect 512864 369802 512920 369836
rect 512954 369802 513010 369836
rect 513044 369802 513100 369836
rect 513134 369802 513188 369836
rect 512508 369746 513188 369802
rect 512508 369712 512560 369746
rect 512594 369712 512650 369746
rect 512684 369712 512740 369746
rect 512774 369712 512830 369746
rect 512864 369712 512920 369746
rect 512954 369712 513010 369746
rect 513044 369712 513100 369746
rect 513134 369712 513188 369746
rect 512508 369656 513188 369712
rect 512508 369622 512560 369656
rect 512594 369622 512650 369656
rect 512684 369622 512740 369656
rect 512774 369622 512830 369656
rect 512864 369622 512920 369656
rect 512954 369622 513010 369656
rect 513044 369622 513100 369656
rect 513134 369622 513188 369656
rect 512508 369566 513188 369622
rect 512508 369532 512560 369566
rect 512594 369532 512650 369566
rect 512684 369532 512740 369566
rect 512774 369532 512830 369566
rect 512864 369532 512920 369566
rect 512954 369532 513010 369566
rect 513044 369532 513100 369566
rect 513134 369532 513188 369566
rect 512508 369480 513188 369532
rect 523423 371757 524713 371769
rect 523423 371723 523439 371757
rect 523473 371723 523507 371757
rect 523541 371723 523575 371757
rect 523609 371723 523643 371757
rect 523677 371723 523711 371757
rect 523745 371723 523779 371757
rect 523813 371723 523847 371757
rect 523881 371723 523915 371757
rect 523949 371723 523983 371757
rect 524017 371723 524051 371757
rect 524085 371723 524119 371757
rect 524153 371723 524187 371757
rect 524221 371723 524255 371757
rect 524289 371723 524323 371757
rect 524357 371723 524391 371757
rect 524425 371723 524459 371757
rect 524493 371723 524527 371757
rect 524561 371723 524595 371757
rect 524629 371723 524663 371757
rect 524697 371723 524713 371757
rect 523423 371711 524713 371723
rect 523423 371299 524713 371311
rect 523423 371265 523439 371299
rect 523473 371265 523507 371299
rect 523541 371265 523575 371299
rect 523609 371265 523643 371299
rect 523677 371265 523711 371299
rect 523745 371265 523779 371299
rect 523813 371265 523847 371299
rect 523881 371265 523915 371299
rect 523949 371265 523983 371299
rect 524017 371265 524051 371299
rect 524085 371265 524119 371299
rect 524153 371265 524187 371299
rect 524221 371265 524255 371299
rect 524289 371265 524323 371299
rect 524357 371265 524391 371299
rect 524425 371265 524459 371299
rect 524493 371265 524527 371299
rect 524561 371265 524595 371299
rect 524629 371265 524663 371299
rect 524697 371265 524713 371299
rect 523423 371253 524713 371265
rect 523423 370841 524713 370853
rect 523423 370807 523439 370841
rect 523473 370807 523507 370841
rect 523541 370807 523575 370841
rect 523609 370807 523643 370841
rect 523677 370807 523711 370841
rect 523745 370807 523779 370841
rect 523813 370807 523847 370841
rect 523881 370807 523915 370841
rect 523949 370807 523983 370841
rect 524017 370807 524051 370841
rect 524085 370807 524119 370841
rect 524153 370807 524187 370841
rect 524221 370807 524255 370841
rect 524289 370807 524323 370841
rect 524357 370807 524391 370841
rect 524425 370807 524459 370841
rect 524493 370807 524527 370841
rect 524561 370807 524595 370841
rect 524629 370807 524663 370841
rect 524697 370807 524713 370841
rect 523423 370795 524713 370807
rect 523423 370383 524713 370395
rect 523423 370349 523439 370383
rect 523473 370349 523507 370383
rect 523541 370349 523575 370383
rect 523609 370349 523643 370383
rect 523677 370349 523711 370383
rect 523745 370349 523779 370383
rect 523813 370349 523847 370383
rect 523881 370349 523915 370383
rect 523949 370349 523983 370383
rect 524017 370349 524051 370383
rect 524085 370349 524119 370383
rect 524153 370349 524187 370383
rect 524221 370349 524255 370383
rect 524289 370349 524323 370383
rect 524357 370349 524391 370383
rect 524425 370349 524459 370383
rect 524493 370349 524527 370383
rect 524561 370349 524595 370383
rect 524629 370349 524663 370383
rect 524697 370349 524713 370383
rect 523423 370337 524713 370349
rect 523423 369925 524713 369937
rect 523423 369891 523439 369925
rect 523473 369891 523507 369925
rect 523541 369891 523575 369925
rect 523609 369891 523643 369925
rect 523677 369891 523711 369925
rect 523745 369891 523779 369925
rect 523813 369891 523847 369925
rect 523881 369891 523915 369925
rect 523949 369891 523983 369925
rect 524017 369891 524051 369925
rect 524085 369891 524119 369925
rect 524153 369891 524187 369925
rect 524221 369891 524255 369925
rect 524289 369891 524323 369925
rect 524357 369891 524391 369925
rect 524425 369891 524459 369925
rect 524493 369891 524527 369925
rect 524561 369891 524595 369925
rect 524629 369891 524663 369925
rect 524697 369891 524713 369925
rect 523423 369879 524713 369891
rect 523423 369467 524713 369479
rect 523423 369433 523439 369467
rect 523473 369433 523507 369467
rect 523541 369433 523575 369467
rect 523609 369433 523643 369467
rect 523677 369433 523711 369467
rect 523745 369433 523779 369467
rect 523813 369433 523847 369467
rect 523881 369433 523915 369467
rect 523949 369433 523983 369467
rect 524017 369433 524051 369467
rect 524085 369433 524119 369467
rect 524153 369433 524187 369467
rect 524221 369433 524255 369467
rect 524289 369433 524323 369467
rect 524357 369433 524391 369467
rect 524425 369433 524459 369467
rect 524493 369433 524527 369467
rect 524561 369433 524595 369467
rect 524629 369433 524663 369467
rect 524697 369433 524713 369467
rect 523423 369421 524713 369433
rect 512508 368766 513188 368820
rect 512508 368732 512560 368766
rect 512594 368732 512650 368766
rect 512684 368732 512740 368766
rect 512774 368732 512830 368766
rect 512864 368732 512920 368766
rect 512954 368732 513010 368766
rect 513044 368732 513100 368766
rect 513134 368732 513188 368766
rect 512508 368676 513188 368732
rect 512508 368642 512560 368676
rect 512594 368642 512650 368676
rect 512684 368642 512740 368676
rect 512774 368642 512830 368676
rect 512864 368642 512920 368676
rect 512954 368642 513010 368676
rect 513044 368642 513100 368676
rect 513134 368642 513188 368676
rect 512508 368586 513188 368642
rect 512508 368552 512560 368586
rect 512594 368552 512650 368586
rect 512684 368552 512740 368586
rect 512774 368552 512830 368586
rect 512864 368552 512920 368586
rect 512954 368552 513010 368586
rect 513044 368552 513100 368586
rect 513134 368552 513188 368586
rect 512508 368496 513188 368552
rect 512508 368462 512560 368496
rect 512594 368462 512650 368496
rect 512684 368462 512740 368496
rect 512774 368462 512830 368496
rect 512864 368462 512920 368496
rect 512954 368462 513010 368496
rect 513044 368462 513100 368496
rect 513134 368462 513188 368496
rect 512508 368406 513188 368462
rect 512508 368372 512560 368406
rect 512594 368372 512650 368406
rect 512684 368372 512740 368406
rect 512774 368372 512830 368406
rect 512864 368372 512920 368406
rect 512954 368372 513010 368406
rect 513044 368372 513100 368406
rect 513134 368372 513188 368406
rect 512508 368316 513188 368372
rect 512508 368282 512560 368316
rect 512594 368282 512650 368316
rect 512684 368282 512740 368316
rect 512774 368282 512830 368316
rect 512864 368282 512920 368316
rect 512954 368282 513010 368316
rect 513044 368282 513100 368316
rect 513134 368282 513188 368316
rect 512508 368226 513188 368282
rect 512508 368192 512560 368226
rect 512594 368192 512650 368226
rect 512684 368192 512740 368226
rect 512774 368192 512830 368226
rect 512864 368192 512920 368226
rect 512954 368192 513010 368226
rect 513044 368192 513100 368226
rect 513134 368192 513188 368226
rect 512508 368140 513188 368192
rect 512508 367426 513188 367480
rect 512508 367392 512560 367426
rect 512594 367392 512650 367426
rect 512684 367392 512740 367426
rect 512774 367392 512830 367426
rect 512864 367392 512920 367426
rect 512954 367392 513010 367426
rect 513044 367392 513100 367426
rect 513134 367392 513188 367426
rect 512508 367336 513188 367392
rect 512508 367302 512560 367336
rect 512594 367302 512650 367336
rect 512684 367302 512740 367336
rect 512774 367302 512830 367336
rect 512864 367302 512920 367336
rect 512954 367302 513010 367336
rect 513044 367302 513100 367336
rect 513134 367302 513188 367336
rect 512508 367246 513188 367302
rect 512508 367212 512560 367246
rect 512594 367212 512650 367246
rect 512684 367212 512740 367246
rect 512774 367212 512830 367246
rect 512864 367212 512920 367246
rect 512954 367212 513010 367246
rect 513044 367212 513100 367246
rect 513134 367212 513188 367246
rect 512508 367156 513188 367212
rect 512508 367122 512560 367156
rect 512594 367122 512650 367156
rect 512684 367122 512740 367156
rect 512774 367122 512830 367156
rect 512864 367122 512920 367156
rect 512954 367122 513010 367156
rect 513044 367122 513100 367156
rect 513134 367122 513188 367156
rect 512508 367066 513188 367122
rect 512508 367032 512560 367066
rect 512594 367032 512650 367066
rect 512684 367032 512740 367066
rect 512774 367032 512830 367066
rect 512864 367032 512920 367066
rect 512954 367032 513010 367066
rect 513044 367032 513100 367066
rect 513134 367032 513188 367066
rect 512508 366976 513188 367032
rect 512508 366942 512560 366976
rect 512594 366942 512650 366976
rect 512684 366942 512740 366976
rect 512774 366942 512830 366976
rect 512864 366942 512920 366976
rect 512954 366942 513010 366976
rect 513044 366942 513100 366976
rect 513134 366942 513188 366976
rect 512508 366886 513188 366942
rect 512508 366852 512560 366886
rect 512594 366852 512650 366886
rect 512684 366852 512740 366886
rect 512774 366852 512830 366886
rect 512864 366852 512920 366886
rect 512954 366852 513010 366886
rect 513044 366852 513100 366886
rect 513134 366852 513188 366886
rect 512508 366800 513188 366852
rect 523423 369009 524713 369021
rect 523423 368975 523439 369009
rect 523473 368975 523507 369009
rect 523541 368975 523575 369009
rect 523609 368975 523643 369009
rect 523677 368975 523711 369009
rect 523745 368975 523779 369009
rect 523813 368975 523847 369009
rect 523881 368975 523915 369009
rect 523949 368975 523983 369009
rect 524017 368975 524051 369009
rect 524085 368975 524119 369009
rect 524153 368975 524187 369009
rect 524221 368975 524255 369009
rect 524289 368975 524323 369009
rect 524357 368975 524391 369009
rect 524425 368975 524459 369009
rect 524493 368975 524527 369009
rect 524561 368975 524595 369009
rect 524629 368975 524663 369009
rect 524697 368975 524713 369009
rect 523423 368963 524713 368975
rect 523423 368551 524713 368563
rect 523423 368517 523439 368551
rect 523473 368517 523507 368551
rect 523541 368517 523575 368551
rect 523609 368517 523643 368551
rect 523677 368517 523711 368551
rect 523745 368517 523779 368551
rect 523813 368517 523847 368551
rect 523881 368517 523915 368551
rect 523949 368517 523983 368551
rect 524017 368517 524051 368551
rect 524085 368517 524119 368551
rect 524153 368517 524187 368551
rect 524221 368517 524255 368551
rect 524289 368517 524323 368551
rect 524357 368517 524391 368551
rect 524425 368517 524459 368551
rect 524493 368517 524527 368551
rect 524561 368517 524595 368551
rect 524629 368517 524663 368551
rect 524697 368517 524713 368551
rect 523423 368505 524713 368517
rect 523423 368093 524713 368105
rect 523423 368059 523439 368093
rect 523473 368059 523507 368093
rect 523541 368059 523575 368093
rect 523609 368059 523643 368093
rect 523677 368059 523711 368093
rect 523745 368059 523779 368093
rect 523813 368059 523847 368093
rect 523881 368059 523915 368093
rect 523949 368059 523983 368093
rect 524017 368059 524051 368093
rect 524085 368059 524119 368093
rect 524153 368059 524187 368093
rect 524221 368059 524255 368093
rect 524289 368059 524323 368093
rect 524357 368059 524391 368093
rect 524425 368059 524459 368093
rect 524493 368059 524527 368093
rect 524561 368059 524595 368093
rect 524629 368059 524663 368093
rect 524697 368059 524713 368093
rect 523423 368047 524713 368059
rect 523423 367635 524713 367647
rect 523423 367601 523439 367635
rect 523473 367601 523507 367635
rect 523541 367601 523575 367635
rect 523609 367601 523643 367635
rect 523677 367601 523711 367635
rect 523745 367601 523779 367635
rect 523813 367601 523847 367635
rect 523881 367601 523915 367635
rect 523949 367601 523983 367635
rect 524017 367601 524051 367635
rect 524085 367601 524119 367635
rect 524153 367601 524187 367635
rect 524221 367601 524255 367635
rect 524289 367601 524323 367635
rect 524357 367601 524391 367635
rect 524425 367601 524459 367635
rect 524493 367601 524527 367635
rect 524561 367601 524595 367635
rect 524629 367601 524663 367635
rect 524697 367601 524713 367635
rect 523423 367589 524713 367601
rect 523423 367177 524713 367189
rect 523423 367143 523439 367177
rect 523473 367143 523507 367177
rect 523541 367143 523575 367177
rect 523609 367143 523643 367177
rect 523677 367143 523711 367177
rect 523745 367143 523779 367177
rect 523813 367143 523847 367177
rect 523881 367143 523915 367177
rect 523949 367143 523983 367177
rect 524017 367143 524051 367177
rect 524085 367143 524119 367177
rect 524153 367143 524187 367177
rect 524221 367143 524255 367177
rect 524289 367143 524323 367177
rect 524357 367143 524391 367177
rect 524425 367143 524459 367177
rect 524493 367143 524527 367177
rect 524561 367143 524595 367177
rect 524629 367143 524663 367177
rect 524697 367143 524713 367177
rect 523423 367131 524713 367143
rect 523423 366719 524713 366731
rect 523423 366685 523439 366719
rect 523473 366685 523507 366719
rect 523541 366685 523575 366719
rect 523609 366685 523643 366719
rect 523677 366685 523711 366719
rect 523745 366685 523779 366719
rect 523813 366685 523847 366719
rect 523881 366685 523915 366719
rect 523949 366685 523983 366719
rect 524017 366685 524051 366719
rect 524085 366685 524119 366719
rect 524153 366685 524187 366719
rect 524221 366685 524255 366719
rect 524289 366685 524323 366719
rect 524357 366685 524391 366719
rect 524425 366685 524459 366719
rect 524493 366685 524527 366719
rect 524561 366685 524595 366719
rect 524629 366685 524663 366719
rect 524697 366685 524713 366719
rect 523423 366673 524713 366685
rect 512508 366086 513188 366140
rect 512508 366052 512560 366086
rect 512594 366052 512650 366086
rect 512684 366052 512740 366086
rect 512774 366052 512830 366086
rect 512864 366052 512920 366086
rect 512954 366052 513010 366086
rect 513044 366052 513100 366086
rect 513134 366052 513188 366086
rect 512508 365996 513188 366052
rect 512508 365962 512560 365996
rect 512594 365962 512650 365996
rect 512684 365962 512740 365996
rect 512774 365962 512830 365996
rect 512864 365962 512920 365996
rect 512954 365962 513010 365996
rect 513044 365962 513100 365996
rect 513134 365962 513188 365996
rect 512508 365906 513188 365962
rect 512508 365872 512560 365906
rect 512594 365872 512650 365906
rect 512684 365872 512740 365906
rect 512774 365872 512830 365906
rect 512864 365872 512920 365906
rect 512954 365872 513010 365906
rect 513044 365872 513100 365906
rect 513134 365872 513188 365906
rect 512508 365816 513188 365872
rect 512508 365782 512560 365816
rect 512594 365782 512650 365816
rect 512684 365782 512740 365816
rect 512774 365782 512830 365816
rect 512864 365782 512920 365816
rect 512954 365782 513010 365816
rect 513044 365782 513100 365816
rect 513134 365782 513188 365816
rect 512508 365726 513188 365782
rect 512508 365692 512560 365726
rect 512594 365692 512650 365726
rect 512684 365692 512740 365726
rect 512774 365692 512830 365726
rect 512864 365692 512920 365726
rect 512954 365692 513010 365726
rect 513044 365692 513100 365726
rect 513134 365692 513188 365726
rect 512508 365636 513188 365692
rect 512508 365602 512560 365636
rect 512594 365602 512650 365636
rect 512684 365602 512740 365636
rect 512774 365602 512830 365636
rect 512864 365602 512920 365636
rect 512954 365602 513010 365636
rect 513044 365602 513100 365636
rect 513134 365602 513188 365636
rect 512508 365546 513188 365602
rect 512508 365512 512560 365546
rect 512594 365512 512650 365546
rect 512684 365512 512740 365546
rect 512774 365512 512830 365546
rect 512864 365512 512920 365546
rect 512954 365512 513010 365546
rect 513044 365512 513100 365546
rect 513134 365512 513188 365546
rect 512508 365460 513188 365512
rect 512508 364746 513188 364800
rect 512508 364712 512560 364746
rect 512594 364712 512650 364746
rect 512684 364712 512740 364746
rect 512774 364712 512830 364746
rect 512864 364712 512920 364746
rect 512954 364712 513010 364746
rect 513044 364712 513100 364746
rect 513134 364712 513188 364746
rect 512508 364656 513188 364712
rect 512508 364622 512560 364656
rect 512594 364622 512650 364656
rect 512684 364622 512740 364656
rect 512774 364622 512830 364656
rect 512864 364622 512920 364656
rect 512954 364622 513010 364656
rect 513044 364622 513100 364656
rect 513134 364622 513188 364656
rect 512508 364566 513188 364622
rect 512508 364532 512560 364566
rect 512594 364532 512650 364566
rect 512684 364532 512740 364566
rect 512774 364532 512830 364566
rect 512864 364532 512920 364566
rect 512954 364532 513010 364566
rect 513044 364532 513100 364566
rect 513134 364532 513188 364566
rect 512508 364476 513188 364532
rect 512508 364442 512560 364476
rect 512594 364442 512650 364476
rect 512684 364442 512740 364476
rect 512774 364442 512830 364476
rect 512864 364442 512920 364476
rect 512954 364442 513010 364476
rect 513044 364442 513100 364476
rect 513134 364442 513188 364476
rect 512508 364386 513188 364442
rect 512508 364352 512560 364386
rect 512594 364352 512650 364386
rect 512684 364352 512740 364386
rect 512774 364352 512830 364386
rect 512864 364352 512920 364386
rect 512954 364352 513010 364386
rect 513044 364352 513100 364386
rect 513134 364352 513188 364386
rect 512508 364296 513188 364352
rect 512508 364262 512560 364296
rect 512594 364262 512650 364296
rect 512684 364262 512740 364296
rect 512774 364262 512830 364296
rect 512864 364262 512920 364296
rect 512954 364262 513010 364296
rect 513044 364262 513100 364296
rect 513134 364262 513188 364296
rect 512508 364206 513188 364262
rect 512508 364172 512560 364206
rect 512594 364172 512650 364206
rect 512684 364172 512740 364206
rect 512774 364172 512830 364206
rect 512864 364172 512920 364206
rect 512954 364172 513010 364206
rect 513044 364172 513100 364206
rect 513134 364172 513188 364206
rect 512508 364120 513188 364172
rect 523423 366261 524713 366273
rect 523423 366227 523439 366261
rect 523473 366227 523507 366261
rect 523541 366227 523575 366261
rect 523609 366227 523643 366261
rect 523677 366227 523711 366261
rect 523745 366227 523779 366261
rect 523813 366227 523847 366261
rect 523881 366227 523915 366261
rect 523949 366227 523983 366261
rect 524017 366227 524051 366261
rect 524085 366227 524119 366261
rect 524153 366227 524187 366261
rect 524221 366227 524255 366261
rect 524289 366227 524323 366261
rect 524357 366227 524391 366261
rect 524425 366227 524459 366261
rect 524493 366227 524527 366261
rect 524561 366227 524595 366261
rect 524629 366227 524663 366261
rect 524697 366227 524713 366261
rect 523423 366215 524713 366227
rect 523423 365803 524713 365815
rect 523423 365769 523439 365803
rect 523473 365769 523507 365803
rect 523541 365769 523575 365803
rect 523609 365769 523643 365803
rect 523677 365769 523711 365803
rect 523745 365769 523779 365803
rect 523813 365769 523847 365803
rect 523881 365769 523915 365803
rect 523949 365769 523983 365803
rect 524017 365769 524051 365803
rect 524085 365769 524119 365803
rect 524153 365769 524187 365803
rect 524221 365769 524255 365803
rect 524289 365769 524323 365803
rect 524357 365769 524391 365803
rect 524425 365769 524459 365803
rect 524493 365769 524527 365803
rect 524561 365769 524595 365803
rect 524629 365769 524663 365803
rect 524697 365769 524713 365803
rect 523423 365757 524713 365769
rect 523423 365345 524713 365357
rect 523423 365311 523439 365345
rect 523473 365311 523507 365345
rect 523541 365311 523575 365345
rect 523609 365311 523643 365345
rect 523677 365311 523711 365345
rect 523745 365311 523779 365345
rect 523813 365311 523847 365345
rect 523881 365311 523915 365345
rect 523949 365311 523983 365345
rect 524017 365311 524051 365345
rect 524085 365311 524119 365345
rect 524153 365311 524187 365345
rect 524221 365311 524255 365345
rect 524289 365311 524323 365345
rect 524357 365311 524391 365345
rect 524425 365311 524459 365345
rect 524493 365311 524527 365345
rect 524561 365311 524595 365345
rect 524629 365311 524663 365345
rect 524697 365311 524713 365345
rect 523423 365299 524713 365311
rect 523423 364887 524713 364899
rect 523423 364853 523439 364887
rect 523473 364853 523507 364887
rect 523541 364853 523575 364887
rect 523609 364853 523643 364887
rect 523677 364853 523711 364887
rect 523745 364853 523779 364887
rect 523813 364853 523847 364887
rect 523881 364853 523915 364887
rect 523949 364853 523983 364887
rect 524017 364853 524051 364887
rect 524085 364853 524119 364887
rect 524153 364853 524187 364887
rect 524221 364853 524255 364887
rect 524289 364853 524323 364887
rect 524357 364853 524391 364887
rect 524425 364853 524459 364887
rect 524493 364853 524527 364887
rect 524561 364853 524595 364887
rect 524629 364853 524663 364887
rect 524697 364853 524713 364887
rect 523423 364841 524713 364853
rect 523423 364429 524713 364441
rect 523423 364395 523439 364429
rect 523473 364395 523507 364429
rect 523541 364395 523575 364429
rect 523609 364395 523643 364429
rect 523677 364395 523711 364429
rect 523745 364395 523779 364429
rect 523813 364395 523847 364429
rect 523881 364395 523915 364429
rect 523949 364395 523983 364429
rect 524017 364395 524051 364429
rect 524085 364395 524119 364429
rect 524153 364395 524187 364429
rect 524221 364395 524255 364429
rect 524289 364395 524323 364429
rect 524357 364395 524391 364429
rect 524425 364395 524459 364429
rect 524493 364395 524527 364429
rect 524561 364395 524595 364429
rect 524629 364395 524663 364429
rect 524697 364395 524713 364429
rect 523423 364383 524713 364395
rect 523423 363971 524713 363983
rect 523423 363937 523439 363971
rect 523473 363937 523507 363971
rect 523541 363937 523575 363971
rect 523609 363937 523643 363971
rect 523677 363937 523711 363971
rect 523745 363937 523779 363971
rect 523813 363937 523847 363971
rect 523881 363937 523915 363971
rect 523949 363937 523983 363971
rect 524017 363937 524051 363971
rect 524085 363937 524119 363971
rect 524153 363937 524187 363971
rect 524221 363937 524255 363971
rect 524289 363937 524323 363971
rect 524357 363937 524391 363971
rect 524425 363937 524459 363971
rect 524493 363937 524527 363971
rect 524561 363937 524595 363971
rect 524629 363937 524663 363971
rect 524697 363937 524713 363971
rect 523423 363925 524713 363937
rect 512508 363406 513188 363460
rect 512508 363372 512560 363406
rect 512594 363372 512650 363406
rect 512684 363372 512740 363406
rect 512774 363372 512830 363406
rect 512864 363372 512920 363406
rect 512954 363372 513010 363406
rect 513044 363372 513100 363406
rect 513134 363372 513188 363406
rect 512508 363316 513188 363372
rect 512508 363282 512560 363316
rect 512594 363282 512650 363316
rect 512684 363282 512740 363316
rect 512774 363282 512830 363316
rect 512864 363282 512920 363316
rect 512954 363282 513010 363316
rect 513044 363282 513100 363316
rect 513134 363282 513188 363316
rect 512508 363226 513188 363282
rect 512508 363192 512560 363226
rect 512594 363192 512650 363226
rect 512684 363192 512740 363226
rect 512774 363192 512830 363226
rect 512864 363192 512920 363226
rect 512954 363192 513010 363226
rect 513044 363192 513100 363226
rect 513134 363192 513188 363226
rect 512508 363136 513188 363192
rect 512508 363102 512560 363136
rect 512594 363102 512650 363136
rect 512684 363102 512740 363136
rect 512774 363102 512830 363136
rect 512864 363102 512920 363136
rect 512954 363102 513010 363136
rect 513044 363102 513100 363136
rect 513134 363102 513188 363136
rect 512508 363046 513188 363102
rect 512508 363012 512560 363046
rect 512594 363012 512650 363046
rect 512684 363012 512740 363046
rect 512774 363012 512830 363046
rect 512864 363012 512920 363046
rect 512954 363012 513010 363046
rect 513044 363012 513100 363046
rect 513134 363012 513188 363046
rect 512508 362956 513188 363012
rect 512508 362922 512560 362956
rect 512594 362922 512650 362956
rect 512684 362922 512740 362956
rect 512774 362922 512830 362956
rect 512864 362922 512920 362956
rect 512954 362922 513010 362956
rect 513044 362922 513100 362956
rect 513134 362922 513188 362956
rect 512508 362866 513188 362922
rect 512508 362832 512560 362866
rect 512594 362832 512650 362866
rect 512684 362832 512740 362866
rect 512774 362832 512830 362866
rect 512864 362832 512920 362866
rect 512954 362832 513010 362866
rect 513044 362832 513100 362866
rect 513134 362832 513188 362866
rect 512508 362780 513188 362832
rect 523423 363513 524713 363525
rect 523423 363479 523439 363513
rect 523473 363479 523507 363513
rect 523541 363479 523575 363513
rect 523609 363479 523643 363513
rect 523677 363479 523711 363513
rect 523745 363479 523779 363513
rect 523813 363479 523847 363513
rect 523881 363479 523915 363513
rect 523949 363479 523983 363513
rect 524017 363479 524051 363513
rect 524085 363479 524119 363513
rect 524153 363479 524187 363513
rect 524221 363479 524255 363513
rect 524289 363479 524323 363513
rect 524357 363479 524391 363513
rect 524425 363479 524459 363513
rect 524493 363479 524527 363513
rect 524561 363479 524595 363513
rect 524629 363479 524663 363513
rect 524697 363479 524713 363513
rect 523423 363467 524713 363479
rect 523423 363055 524713 363067
rect 523423 363021 523439 363055
rect 523473 363021 523507 363055
rect 523541 363021 523575 363055
rect 523609 363021 523643 363055
rect 523677 363021 523711 363055
rect 523745 363021 523779 363055
rect 523813 363021 523847 363055
rect 523881 363021 523915 363055
rect 523949 363021 523983 363055
rect 524017 363021 524051 363055
rect 524085 363021 524119 363055
rect 524153 363021 524187 363055
rect 524221 363021 524255 363055
rect 524289 363021 524323 363055
rect 524357 363021 524391 363055
rect 524425 363021 524459 363055
rect 524493 363021 524527 363055
rect 524561 363021 524595 363055
rect 524629 363021 524663 363055
rect 524697 363021 524713 363055
rect 523423 363009 524713 363021
rect 523423 362597 524713 362609
rect 523423 362563 523439 362597
rect 523473 362563 523507 362597
rect 523541 362563 523575 362597
rect 523609 362563 523643 362597
rect 523677 362563 523711 362597
rect 523745 362563 523779 362597
rect 523813 362563 523847 362597
rect 523881 362563 523915 362597
rect 523949 362563 523983 362597
rect 524017 362563 524051 362597
rect 524085 362563 524119 362597
rect 524153 362563 524187 362597
rect 524221 362563 524255 362597
rect 524289 362563 524323 362597
rect 524357 362563 524391 362597
rect 524425 362563 524459 362597
rect 524493 362563 524527 362597
rect 524561 362563 524595 362597
rect 524629 362563 524663 362597
rect 524697 362563 524713 362597
rect 523423 362551 524713 362563
rect 574679 358898 574737 358910
rect 574679 357922 574691 358898
rect 574725 357922 574737 358898
rect 574679 357910 574737 357922
rect 574937 358898 574995 358910
rect 574937 357922 574949 358898
rect 574983 357922 574995 358898
rect 574937 357910 574995 357922
rect 575195 358898 575253 358910
rect 575195 357922 575207 358898
rect 575241 357922 575253 358898
rect 575195 357910 575253 357922
rect 575453 358898 575511 358910
rect 575453 357922 575465 358898
rect 575499 357922 575511 358898
rect 575453 357910 575511 357922
rect 575711 358898 575769 358910
rect 575711 357922 575723 358898
rect 575757 357922 575769 358898
rect 575711 357910 575769 357922
rect 575969 358898 576027 358910
rect 575969 357922 575981 358898
rect 576015 357922 576027 358898
rect 575969 357910 576027 357922
rect 576227 358898 576285 358910
rect 576227 357922 576239 358898
rect 576273 357922 576285 358898
rect 576227 357910 576285 357922
rect 576485 358898 576543 358910
rect 576485 357922 576497 358898
rect 576531 357922 576543 358898
rect 576485 357910 576543 357922
rect 576743 358898 576801 358910
rect 576743 357922 576755 358898
rect 576789 357922 576801 358898
rect 576743 357910 576801 357922
rect 577001 358898 577059 358910
rect 577001 357922 577013 358898
rect 577047 357922 577059 358898
rect 577001 357910 577059 357922
rect 577259 358898 577317 358910
rect 577259 357922 577271 358898
rect 577305 357922 577317 358898
rect 577259 357910 577317 357922
rect 577517 358898 577575 358910
rect 577517 357922 577529 358898
rect 577563 357922 577575 358898
rect 577517 357910 577575 357922
rect 577775 358898 577833 358910
rect 577775 357922 577787 358898
rect 577821 357922 577833 358898
rect 577775 357910 577833 357922
rect 578033 358898 578091 358910
rect 578033 357922 578045 358898
rect 578079 357922 578091 358898
rect 578033 357910 578091 357922
rect 578291 358898 578349 358910
rect 578291 357922 578303 358898
rect 578337 357922 578349 358898
rect 578291 357910 578349 357922
rect 578549 358898 578607 358910
rect 578549 357922 578561 358898
rect 578595 357922 578607 358898
rect 578549 357910 578607 357922
rect 578807 358898 578865 358910
rect 578807 357922 578819 358898
rect 578853 357922 578865 358898
rect 578807 357910 578865 357922
rect 579065 358898 579123 358910
rect 579065 357922 579077 358898
rect 579111 357922 579123 358898
rect 579065 357910 579123 357922
rect 579323 358898 579381 358910
rect 579323 357922 579335 358898
rect 579369 357922 579381 358898
rect 579323 357910 579381 357922
rect 579581 358898 579639 358910
rect 579581 357922 579593 358898
rect 579627 357922 579639 358898
rect 579581 357910 579639 357922
rect 579839 358898 579897 358910
rect 579839 357922 579851 358898
rect 579885 357922 579897 358898
rect 579839 357910 579897 357922
rect 575127 312730 575185 312742
rect 575127 311754 575139 312730
rect 575173 311754 575185 312730
rect 575127 311742 575185 311754
rect 575385 312730 575443 312742
rect 575385 311754 575397 312730
rect 575431 311754 575443 312730
rect 575385 311742 575443 311754
rect 575643 312730 575701 312742
rect 575643 311754 575655 312730
rect 575689 311754 575701 312730
rect 575643 311742 575701 311754
rect 575901 312730 575959 312742
rect 575901 311754 575913 312730
rect 575947 311754 575959 312730
rect 575901 311742 575959 311754
rect 576159 312730 576217 312742
rect 576159 311754 576171 312730
rect 576205 311754 576217 312730
rect 576159 311742 576217 311754
rect 576417 312730 576475 312742
rect 576417 311754 576429 312730
rect 576463 311754 576475 312730
rect 576417 311742 576475 311754
rect 576675 312730 576733 312742
rect 576675 311754 576687 312730
rect 576721 311754 576733 312730
rect 576675 311742 576733 311754
rect 576933 312730 576991 312742
rect 576933 311754 576945 312730
rect 576979 311754 576991 312730
rect 576933 311742 576991 311754
rect 577191 312730 577249 312742
rect 577191 311754 577203 312730
rect 577237 311754 577249 312730
rect 577191 311742 577249 311754
rect 577449 312730 577507 312742
rect 577449 311754 577461 312730
rect 577495 311754 577507 312730
rect 577449 311742 577507 311754
rect 577707 312730 577765 312742
rect 577707 311754 577719 312730
rect 577753 311754 577765 312730
rect 577707 311742 577765 311754
rect 577965 312730 578023 312742
rect 577965 311754 577977 312730
rect 578011 311754 578023 312730
rect 577965 311742 578023 311754
rect 578223 312730 578281 312742
rect 578223 311754 578235 312730
rect 578269 311754 578281 312730
rect 578223 311742 578281 311754
rect 578481 312730 578539 312742
rect 578481 311754 578493 312730
rect 578527 311754 578539 312730
rect 578481 311742 578539 311754
rect 578739 312730 578797 312742
rect 578739 311754 578751 312730
rect 578785 311754 578797 312730
rect 578739 311742 578797 311754
rect 578997 312730 579055 312742
rect 578997 311754 579009 312730
rect 579043 311754 579055 312730
rect 578997 311742 579055 311754
rect 579255 312730 579313 312742
rect 579255 311754 579267 312730
rect 579301 311754 579313 312730
rect 579255 311742 579313 311754
rect 579513 312730 579571 312742
rect 579513 311754 579525 312730
rect 579559 311754 579571 312730
rect 579513 311742 579571 311754
rect 579771 312730 579829 312742
rect 579771 311754 579783 312730
rect 579817 311754 579829 312730
rect 579771 311742 579829 311754
rect 580029 312730 580087 312742
rect 580029 311754 580041 312730
rect 580075 311754 580087 312730
rect 580029 311742 580087 311754
rect 580287 312730 580345 312742
rect 580287 311754 580299 312730
rect 580333 311754 580345 312730
rect 580287 311742 580345 311754
<< ndiffc >>
rect 560661 492452 560695 493428
rect 560919 492452 560953 493428
rect 561177 492452 561211 493428
rect 561435 492452 561469 493428
rect 561693 492452 561727 493428
rect 561951 492452 561985 493428
rect 562209 492452 562243 493428
rect 562467 492452 562501 493428
rect 562725 492452 562759 493428
rect 562983 492452 563017 493428
rect 563241 492452 563275 493428
rect 563499 492452 563533 493428
rect 563757 492452 563791 493428
rect 564015 492452 564049 493428
rect 564273 492452 564307 493428
rect 564531 492452 564565 493428
rect 564789 492452 564823 493428
rect 565047 492452 565081 493428
rect 565305 492452 565339 493428
rect 565563 492452 565597 493428
rect 565821 492452 565855 493428
rect 560701 403310 560735 404286
rect 560959 403310 560993 404286
rect 561217 403310 561251 404286
rect 561475 403310 561509 404286
rect 561733 403310 561767 404286
rect 561991 403310 562025 404286
rect 562249 403310 562283 404286
rect 562507 403310 562541 404286
rect 562765 403310 562799 404286
rect 563023 403310 563057 404286
rect 563281 403310 563315 404286
rect 563539 403310 563573 404286
rect 563797 403310 563831 404286
rect 564055 403310 564089 404286
rect 564313 403310 564347 404286
rect 564571 403310 564605 404286
rect 564829 403310 564863 404286
rect 565087 403310 565121 404286
rect 565345 403310 565379 404286
rect 565603 403310 565637 404286
rect 565861 403310 565895 404286
rect 497391 400790 497425 400824
rect 497459 400790 497493 400824
rect 497527 400790 497561 400824
rect 497595 400790 497629 400824
rect 497663 400790 497697 400824
rect 497731 400790 497765 400824
rect 497799 400790 497833 400824
rect 497867 400790 497901 400824
rect 497935 400790 497969 400824
rect 498003 400790 498037 400824
rect 498071 400790 498105 400824
rect 497391 400332 497425 400366
rect 497459 400332 497493 400366
rect 497527 400332 497561 400366
rect 497595 400332 497629 400366
rect 497663 400332 497697 400366
rect 497731 400332 497765 400366
rect 497799 400332 497833 400366
rect 497867 400332 497901 400366
rect 497935 400332 497969 400366
rect 498003 400332 498037 400366
rect 498071 400332 498105 400366
rect 493631 390990 493665 391024
rect 493699 390990 493733 391024
rect 493767 390990 493801 391024
rect 493835 390990 493869 391024
rect 493903 390990 493937 391024
rect 493971 390990 494005 391024
rect 494039 390990 494073 391024
rect 494107 390990 494141 391024
rect 494175 390990 494209 391024
rect 494243 390990 494277 391024
rect 494311 390990 494345 391024
rect 493631 390532 493665 390566
rect 493699 390532 493733 390566
rect 493767 390532 493801 390566
rect 493835 390532 493869 390566
rect 493903 390532 493937 390566
rect 493971 390532 494005 390566
rect 494039 390532 494073 390566
rect 494107 390532 494141 390566
rect 494175 390532 494209 390566
rect 494243 390532 494277 390566
rect 494311 390532 494345 390566
rect 504911 389490 504945 389524
rect 504979 389490 505013 389524
rect 505047 389490 505081 389524
rect 505115 389490 505149 389524
rect 505183 389490 505217 389524
rect 505251 389490 505285 389524
rect 505319 389490 505353 389524
rect 505387 389490 505421 389524
rect 505455 389490 505489 389524
rect 505523 389490 505557 389524
rect 505591 389490 505625 389524
rect 516191 389490 516225 389524
rect 516259 389490 516293 389524
rect 516327 389490 516361 389524
rect 516395 389490 516429 389524
rect 516463 389490 516497 389524
rect 516531 389490 516565 389524
rect 516599 389490 516633 389524
rect 516667 389490 516701 389524
rect 516735 389490 516769 389524
rect 516803 389490 516837 389524
rect 516871 389490 516905 389524
rect 504911 389032 504945 389066
rect 504979 389032 505013 389066
rect 505047 389032 505081 389066
rect 505115 389032 505149 389066
rect 505183 389032 505217 389066
rect 505251 389032 505285 389066
rect 505319 389032 505353 389066
rect 505387 389032 505421 389066
rect 505455 389032 505489 389066
rect 505523 389032 505557 389066
rect 505591 389032 505625 389066
rect 516191 389032 516225 389066
rect 516259 389032 516293 389066
rect 516327 389032 516361 389066
rect 516395 389032 516429 389066
rect 516463 389032 516497 389066
rect 516531 389032 516565 389066
rect 516599 389032 516633 389066
rect 516667 389032 516701 389066
rect 516735 389032 516769 389066
rect 516803 389032 516837 389066
rect 516871 389032 516905 389066
rect 504911 388574 504945 388608
rect 504979 388574 505013 388608
rect 505047 388574 505081 388608
rect 505115 388574 505149 388608
rect 505183 388574 505217 388608
rect 505251 388574 505285 388608
rect 505319 388574 505353 388608
rect 505387 388574 505421 388608
rect 505455 388574 505489 388608
rect 505523 388574 505557 388608
rect 505591 388574 505625 388608
rect 516191 388574 516225 388608
rect 516259 388574 516293 388608
rect 516327 388574 516361 388608
rect 516395 388574 516429 388608
rect 516463 388574 516497 388608
rect 516531 388574 516565 388608
rect 516599 388574 516633 388608
rect 516667 388574 516701 388608
rect 516735 388574 516769 388608
rect 516803 388574 516837 388608
rect 516871 388574 516905 388608
rect 504911 388116 504945 388150
rect 504979 388116 505013 388150
rect 505047 388116 505081 388150
rect 505115 388116 505149 388150
rect 505183 388116 505217 388150
rect 505251 388116 505285 388150
rect 505319 388116 505353 388150
rect 505387 388116 505421 388150
rect 505455 388116 505489 388150
rect 505523 388116 505557 388150
rect 505591 388116 505625 388150
rect 516191 388116 516225 388150
rect 516259 388116 516293 388150
rect 516327 388116 516361 388150
rect 516395 388116 516429 388150
rect 516463 388116 516497 388150
rect 516531 388116 516565 388150
rect 516599 388116 516633 388150
rect 516667 388116 516701 388150
rect 516735 388116 516769 388150
rect 516803 388116 516837 388150
rect 516871 388116 516905 388150
rect 504911 387658 504945 387692
rect 504979 387658 505013 387692
rect 505047 387658 505081 387692
rect 505115 387658 505149 387692
rect 505183 387658 505217 387692
rect 505251 387658 505285 387692
rect 505319 387658 505353 387692
rect 505387 387658 505421 387692
rect 505455 387658 505489 387692
rect 505523 387658 505557 387692
rect 505591 387658 505625 387692
rect 504911 387200 504945 387234
rect 504979 387200 505013 387234
rect 505047 387200 505081 387234
rect 505115 387200 505149 387234
rect 505183 387200 505217 387234
rect 505251 387200 505285 387234
rect 505319 387200 505353 387234
rect 505387 387200 505421 387234
rect 505455 387200 505489 387234
rect 505523 387200 505557 387234
rect 505591 387200 505625 387234
rect 504911 386742 504945 386776
rect 504979 386742 505013 386776
rect 505047 386742 505081 386776
rect 505115 386742 505149 386776
rect 505183 386742 505217 386776
rect 505251 386742 505285 386776
rect 505319 386742 505353 386776
rect 505387 386742 505421 386776
rect 505455 386742 505489 386776
rect 505523 386742 505557 386776
rect 505591 386742 505625 386776
rect 504911 386284 504945 386318
rect 504979 386284 505013 386318
rect 505047 386284 505081 386318
rect 505115 386284 505149 386318
rect 505183 386284 505217 386318
rect 505251 386284 505285 386318
rect 505319 386284 505353 386318
rect 505387 386284 505421 386318
rect 505455 386284 505489 386318
rect 505523 386284 505557 386318
rect 505591 386284 505625 386318
rect 504911 385826 504945 385860
rect 504979 385826 505013 385860
rect 505047 385826 505081 385860
rect 505115 385826 505149 385860
rect 505183 385826 505217 385860
rect 505251 385826 505285 385860
rect 505319 385826 505353 385860
rect 505387 385826 505421 385860
rect 505455 385826 505489 385860
rect 505523 385826 505557 385860
rect 505591 385826 505625 385860
rect 504911 385368 504945 385402
rect 504979 385368 505013 385402
rect 505047 385368 505081 385402
rect 505115 385368 505149 385402
rect 505183 385368 505217 385402
rect 505251 385368 505285 385402
rect 505319 385368 505353 385402
rect 505387 385368 505421 385402
rect 505455 385368 505489 385402
rect 505523 385368 505557 385402
rect 505591 385368 505625 385402
rect 516191 387658 516225 387692
rect 516259 387658 516293 387692
rect 516327 387658 516361 387692
rect 516395 387658 516429 387692
rect 516463 387658 516497 387692
rect 516531 387658 516565 387692
rect 516599 387658 516633 387692
rect 516667 387658 516701 387692
rect 516735 387658 516769 387692
rect 516803 387658 516837 387692
rect 516871 387658 516905 387692
rect 516191 387200 516225 387234
rect 516259 387200 516293 387234
rect 516327 387200 516361 387234
rect 516395 387200 516429 387234
rect 516463 387200 516497 387234
rect 516531 387200 516565 387234
rect 516599 387200 516633 387234
rect 516667 387200 516701 387234
rect 516735 387200 516769 387234
rect 516803 387200 516837 387234
rect 516871 387200 516905 387234
rect 516191 386742 516225 386776
rect 516259 386742 516293 386776
rect 516327 386742 516361 386776
rect 516395 386742 516429 386776
rect 516463 386742 516497 386776
rect 516531 386742 516565 386776
rect 516599 386742 516633 386776
rect 516667 386742 516701 386776
rect 516735 386742 516769 386776
rect 516803 386742 516837 386776
rect 516871 386742 516905 386776
rect 516191 386284 516225 386318
rect 516259 386284 516293 386318
rect 516327 386284 516361 386318
rect 516395 386284 516429 386318
rect 516463 386284 516497 386318
rect 516531 386284 516565 386318
rect 516599 386284 516633 386318
rect 516667 386284 516701 386318
rect 516735 386284 516769 386318
rect 516803 386284 516837 386318
rect 516871 386284 516905 386318
rect 516191 385826 516225 385860
rect 516259 385826 516293 385860
rect 516327 385826 516361 385860
rect 516395 385826 516429 385860
rect 516463 385826 516497 385860
rect 516531 385826 516565 385860
rect 516599 385826 516633 385860
rect 516667 385826 516701 385860
rect 516735 385826 516769 385860
rect 516803 385826 516837 385860
rect 516871 385826 516905 385860
rect 516191 385368 516225 385402
rect 516259 385368 516293 385402
rect 516327 385368 516361 385402
rect 516395 385368 516429 385402
rect 516463 385368 516497 385402
rect 516531 385368 516565 385402
rect 516599 385368 516633 385402
rect 516667 385368 516701 385402
rect 516735 385368 516769 385402
rect 516803 385368 516837 385402
rect 516871 385368 516905 385402
rect 501151 377632 501185 377666
rect 501219 377632 501253 377666
rect 501287 377632 501321 377666
rect 501355 377632 501389 377666
rect 501423 377632 501457 377666
rect 501491 377632 501525 377666
rect 501559 377632 501593 377666
rect 501627 377632 501661 377666
rect 501695 377632 501729 377666
rect 501763 377632 501797 377666
rect 501831 377632 501865 377666
rect 501151 377174 501185 377208
rect 501219 377174 501253 377208
rect 501287 377174 501321 377208
rect 501355 377174 501389 377208
rect 501423 377174 501457 377208
rect 501491 377174 501525 377208
rect 501559 377174 501593 377208
rect 501627 377174 501661 377208
rect 501695 377174 501729 377208
rect 501763 377174 501797 377208
rect 501831 377174 501865 377208
rect 501151 376716 501185 376750
rect 501219 376716 501253 376750
rect 501287 376716 501321 376750
rect 501355 376716 501389 376750
rect 501423 376716 501457 376750
rect 501491 376716 501525 376750
rect 501559 376716 501593 376750
rect 501627 376716 501661 376750
rect 501695 376716 501729 376750
rect 501763 376716 501797 376750
rect 501831 376716 501865 376750
rect 501151 376258 501185 376292
rect 501219 376258 501253 376292
rect 501287 376258 501321 376292
rect 501355 376258 501389 376292
rect 501423 376258 501457 376292
rect 501491 376258 501525 376292
rect 501559 376258 501593 376292
rect 501627 376258 501661 376292
rect 501695 376258 501729 376292
rect 501763 376258 501797 376292
rect 501831 376258 501865 376292
rect 501151 375800 501185 375834
rect 501219 375800 501253 375834
rect 501287 375800 501321 375834
rect 501355 375800 501389 375834
rect 501423 375800 501457 375834
rect 501491 375800 501525 375834
rect 501559 375800 501593 375834
rect 501627 375800 501661 375834
rect 501695 375800 501729 375834
rect 501763 375800 501797 375834
rect 501831 375800 501865 375834
rect 501151 375342 501185 375376
rect 501219 375342 501253 375376
rect 501287 375342 501321 375376
rect 501355 375342 501389 375376
rect 501423 375342 501457 375376
rect 501491 375342 501525 375376
rect 501559 375342 501593 375376
rect 501627 375342 501661 375376
rect 501695 375342 501729 375376
rect 501763 375342 501797 375376
rect 501831 375342 501865 375376
rect 501151 374884 501185 374918
rect 501219 374884 501253 374918
rect 501287 374884 501321 374918
rect 501355 374884 501389 374918
rect 501423 374884 501457 374918
rect 501491 374884 501525 374918
rect 501559 374884 501593 374918
rect 501627 374884 501661 374918
rect 501695 374884 501729 374918
rect 501763 374884 501797 374918
rect 501831 374884 501865 374918
rect 501151 374426 501185 374460
rect 501219 374426 501253 374460
rect 501287 374426 501321 374460
rect 501355 374426 501389 374460
rect 501423 374426 501457 374460
rect 501491 374426 501525 374460
rect 501559 374426 501593 374460
rect 501627 374426 501661 374460
rect 501695 374426 501729 374460
rect 501763 374426 501797 374460
rect 501831 374426 501865 374460
rect 501151 373968 501185 374002
rect 501219 373968 501253 374002
rect 501287 373968 501321 374002
rect 501355 373968 501389 374002
rect 501423 373968 501457 374002
rect 501491 373968 501525 374002
rect 501559 373968 501593 374002
rect 501627 373968 501661 374002
rect 501695 373968 501729 374002
rect 501763 373968 501797 374002
rect 501831 373968 501865 374002
rect 501151 373510 501185 373544
rect 501219 373510 501253 373544
rect 501287 373510 501321 373544
rect 501355 373510 501389 373544
rect 501423 373510 501457 373544
rect 501491 373510 501525 373544
rect 501559 373510 501593 373544
rect 501627 373510 501661 373544
rect 501695 373510 501729 373544
rect 501763 373510 501797 373544
rect 501831 373510 501865 373544
rect 560553 357992 560587 358968
rect 560811 357992 560845 358968
rect 561069 357992 561103 358968
rect 561327 357992 561361 358968
rect 561585 357992 561619 358968
rect 561843 357992 561877 358968
rect 562101 357992 562135 358968
rect 562359 357992 562393 358968
rect 562617 357992 562651 358968
rect 562875 357992 562909 358968
rect 563133 357992 563167 358968
rect 563391 357992 563425 358968
rect 563649 357992 563683 358968
rect 563907 357992 563941 358968
rect 564165 357992 564199 358968
rect 564423 357992 564457 358968
rect 564681 357992 564715 358968
rect 564939 357992 564973 358968
rect 565197 357992 565231 358968
rect 565455 357992 565489 358968
rect 565713 357992 565747 358968
rect 560415 311684 560449 312660
rect 560673 311684 560707 312660
rect 560931 311684 560965 312660
rect 561189 311684 561223 312660
rect 561447 311684 561481 312660
rect 561705 311684 561739 312660
rect 561963 311684 561997 312660
rect 562221 311684 562255 312660
rect 562479 311684 562513 312660
rect 562737 311684 562771 312660
rect 562995 311684 563029 312660
rect 563253 311684 563287 312660
rect 563511 311684 563545 312660
rect 563769 311684 563803 312660
rect 564027 311684 564061 312660
rect 564285 311684 564319 312660
rect 564543 311684 564577 312660
rect 564801 311684 564835 312660
rect 565059 311684 565093 312660
rect 565317 311684 565351 312660
rect 565575 311684 565609 312660
<< pdiffc >>
rect 575217 492226 575251 493202
rect 575475 492226 575509 493202
rect 575733 492226 575767 493202
rect 575991 492226 576025 493202
rect 576249 492226 576283 493202
rect 576507 492226 576541 493202
rect 576765 492226 576799 493202
rect 577023 492226 577057 493202
rect 577281 492226 577315 493202
rect 577539 492226 577573 493202
rect 577797 492226 577831 493202
rect 578055 492226 578089 493202
rect 578313 492226 578347 493202
rect 578571 492226 578605 493202
rect 578829 492226 578863 493202
rect 579087 492226 579121 493202
rect 579345 492226 579379 493202
rect 579603 492226 579637 493202
rect 579861 492226 579895 493202
rect 580119 492226 580153 493202
rect 580377 492226 580411 493202
rect 574495 403350 574529 404326
rect 574753 403350 574787 404326
rect 575011 403350 575045 404326
rect 575269 403350 575303 404326
rect 575527 403350 575561 404326
rect 575785 403350 575819 404326
rect 576043 403350 576077 404326
rect 576301 403350 576335 404326
rect 576559 403350 576593 404326
rect 576817 403350 576851 404326
rect 577075 403350 577109 404326
rect 577333 403350 577367 404326
rect 577591 403350 577625 404326
rect 577849 403350 577883 404326
rect 578107 403350 578141 404326
rect 578365 403350 578399 404326
rect 578623 403350 578657 404326
rect 578881 403350 578915 404326
rect 579139 403350 579173 404326
rect 579397 403350 579431 404326
rect 579655 403350 579689 404326
rect 505040 402544 505074 402578
rect 505130 402544 505164 402578
rect 505220 402544 505254 402578
rect 505310 402544 505344 402578
rect 505400 402544 505434 402578
rect 505490 402544 505524 402578
rect 505580 402544 505614 402578
rect 505040 402454 505074 402488
rect 505130 402454 505164 402488
rect 505220 402454 505254 402488
rect 505310 402454 505344 402488
rect 505400 402454 505434 402488
rect 505490 402454 505524 402488
rect 505580 402454 505614 402488
rect 505040 402364 505074 402398
rect 505130 402364 505164 402398
rect 505220 402364 505254 402398
rect 505310 402364 505344 402398
rect 505400 402364 505434 402398
rect 505490 402364 505524 402398
rect 505580 402364 505614 402398
rect 505040 402274 505074 402308
rect 505130 402274 505164 402308
rect 505220 402274 505254 402308
rect 505310 402274 505344 402308
rect 505400 402274 505434 402308
rect 505490 402274 505524 402308
rect 505580 402274 505614 402308
rect 505040 402184 505074 402218
rect 505130 402184 505164 402218
rect 505220 402184 505254 402218
rect 505310 402184 505344 402218
rect 505400 402184 505434 402218
rect 505490 402184 505524 402218
rect 505580 402184 505614 402218
rect 505040 402094 505074 402128
rect 505130 402094 505164 402128
rect 505220 402094 505254 402128
rect 505310 402094 505344 402128
rect 505400 402094 505434 402128
rect 505490 402094 505524 402128
rect 505580 402094 505614 402128
rect 505040 402004 505074 402038
rect 505130 402004 505164 402038
rect 505220 402004 505254 402038
rect 505310 402004 505344 402038
rect 505400 402004 505434 402038
rect 505490 402004 505524 402038
rect 505580 402004 505614 402038
rect 497119 399843 497153 399877
rect 497187 399843 497221 399877
rect 497255 399843 497289 399877
rect 497323 399843 497357 399877
rect 497391 399843 497425 399877
rect 497459 399843 497493 399877
rect 497527 399843 497561 399877
rect 497595 399843 497629 399877
rect 497663 399843 497697 399877
rect 497731 399843 497765 399877
rect 497799 399843 497833 399877
rect 497867 399843 497901 399877
rect 497935 399843 497969 399877
rect 498003 399843 498037 399877
rect 498071 399843 498105 399877
rect 498139 399843 498173 399877
rect 498207 399843 498241 399877
rect 498275 399843 498309 399877
rect 498343 399843 498377 399877
rect 497119 399385 497153 399419
rect 497187 399385 497221 399419
rect 497255 399385 497289 399419
rect 497323 399385 497357 399419
rect 497391 399385 497425 399419
rect 497459 399385 497493 399419
rect 497527 399385 497561 399419
rect 497595 399385 497629 399419
rect 497663 399385 497697 399419
rect 497731 399385 497765 399419
rect 497799 399385 497833 399419
rect 497867 399385 497901 399419
rect 497935 399385 497969 399419
rect 498003 399385 498037 399419
rect 498071 399385 498105 399419
rect 498139 399385 498173 399419
rect 498207 399385 498241 399419
rect 498275 399385 498309 399419
rect 498343 399385 498377 399419
rect 497119 398927 497153 398961
rect 497187 398927 497221 398961
rect 497255 398927 497289 398961
rect 497323 398927 497357 398961
rect 497391 398927 497425 398961
rect 497459 398927 497493 398961
rect 497527 398927 497561 398961
rect 497595 398927 497629 398961
rect 497663 398927 497697 398961
rect 497731 398927 497765 398961
rect 497799 398927 497833 398961
rect 497867 398927 497901 398961
rect 497935 398927 497969 398961
rect 498003 398927 498037 398961
rect 498071 398927 498105 398961
rect 498139 398927 498173 398961
rect 498207 398927 498241 398961
rect 498275 398927 498309 398961
rect 498343 398927 498377 398961
rect 497119 398469 497153 398503
rect 497187 398469 497221 398503
rect 497255 398469 497289 398503
rect 497323 398469 497357 398503
rect 497391 398469 497425 398503
rect 497459 398469 497493 398503
rect 497527 398469 497561 398503
rect 497595 398469 497629 398503
rect 497663 398469 497697 398503
rect 497731 398469 497765 398503
rect 497799 398469 497833 398503
rect 497867 398469 497901 398503
rect 497935 398469 497969 398503
rect 498003 398469 498037 398503
rect 498071 398469 498105 398503
rect 498139 398469 498173 398503
rect 498207 398469 498241 398503
rect 498275 398469 498309 398503
rect 498343 398469 498377 398503
rect 497119 398011 497153 398045
rect 497187 398011 497221 398045
rect 497255 398011 497289 398045
rect 497323 398011 497357 398045
rect 497391 398011 497425 398045
rect 497459 398011 497493 398045
rect 497527 398011 497561 398045
rect 497595 398011 497629 398045
rect 497663 398011 497697 398045
rect 497731 398011 497765 398045
rect 497799 398011 497833 398045
rect 497867 398011 497901 398045
rect 497935 398011 497969 398045
rect 498003 398011 498037 398045
rect 498071 398011 498105 398045
rect 498139 398011 498173 398045
rect 498207 398011 498241 398045
rect 498275 398011 498309 398045
rect 498343 398011 498377 398045
rect 497119 397553 497153 397587
rect 497187 397553 497221 397587
rect 497255 397553 497289 397587
rect 497323 397553 497357 397587
rect 497391 397553 497425 397587
rect 497459 397553 497493 397587
rect 497527 397553 497561 397587
rect 497595 397553 497629 397587
rect 497663 397553 497697 397587
rect 497731 397553 497765 397587
rect 497799 397553 497833 397587
rect 497867 397553 497901 397587
rect 497935 397553 497969 397587
rect 498003 397553 498037 397587
rect 498071 397553 498105 397587
rect 498139 397553 498173 397587
rect 498207 397553 498241 397587
rect 498275 397553 498309 397587
rect 498343 397553 498377 397587
rect 497119 397095 497153 397129
rect 497187 397095 497221 397129
rect 497255 397095 497289 397129
rect 497323 397095 497357 397129
rect 497391 397095 497425 397129
rect 497459 397095 497493 397129
rect 497527 397095 497561 397129
rect 497595 397095 497629 397129
rect 497663 397095 497697 397129
rect 497731 397095 497765 397129
rect 497799 397095 497833 397129
rect 497867 397095 497901 397129
rect 497935 397095 497969 397129
rect 498003 397095 498037 397129
rect 498071 397095 498105 397129
rect 498139 397095 498173 397129
rect 498207 397095 498241 397129
rect 498275 397095 498309 397129
rect 498343 397095 498377 397129
rect 497119 396637 497153 396671
rect 497187 396637 497221 396671
rect 497255 396637 497289 396671
rect 497323 396637 497357 396671
rect 497391 396637 497425 396671
rect 497459 396637 497493 396671
rect 497527 396637 497561 396671
rect 497595 396637 497629 396671
rect 497663 396637 497697 396671
rect 497731 396637 497765 396671
rect 497799 396637 497833 396671
rect 497867 396637 497901 396671
rect 497935 396637 497969 396671
rect 498003 396637 498037 396671
rect 498071 396637 498105 396671
rect 498139 396637 498173 396671
rect 498207 396637 498241 396671
rect 498275 396637 498309 396671
rect 498343 396637 498377 396671
rect 497119 396179 497153 396213
rect 497187 396179 497221 396213
rect 497255 396179 497289 396213
rect 497323 396179 497357 396213
rect 497391 396179 497425 396213
rect 497459 396179 497493 396213
rect 497527 396179 497561 396213
rect 497595 396179 497629 396213
rect 497663 396179 497697 396213
rect 497731 396179 497765 396213
rect 497799 396179 497833 396213
rect 497867 396179 497901 396213
rect 497935 396179 497969 396213
rect 498003 396179 498037 396213
rect 498071 396179 498105 396213
rect 498139 396179 498173 396213
rect 498207 396179 498241 396213
rect 498275 396179 498309 396213
rect 498343 396179 498377 396213
rect 497119 395721 497153 395755
rect 497187 395721 497221 395755
rect 497255 395721 497289 395755
rect 497323 395721 497357 395755
rect 497391 395721 497425 395755
rect 497459 395721 497493 395755
rect 497527 395721 497561 395755
rect 497595 395721 497629 395755
rect 497663 395721 497697 395755
rect 497731 395721 497765 395755
rect 497799 395721 497833 395755
rect 497867 395721 497901 395755
rect 497935 395721 497969 395755
rect 498003 395721 498037 395755
rect 498071 395721 498105 395755
rect 498139 395721 498173 395755
rect 498207 395721 498241 395755
rect 498275 395721 498309 395755
rect 498343 395721 498377 395755
rect 497119 395263 497153 395297
rect 497187 395263 497221 395297
rect 497255 395263 497289 395297
rect 497323 395263 497357 395297
rect 497391 395263 497425 395297
rect 497459 395263 497493 395297
rect 497527 395263 497561 395297
rect 497595 395263 497629 395297
rect 497663 395263 497697 395297
rect 497731 395263 497765 395297
rect 497799 395263 497833 395297
rect 497867 395263 497901 395297
rect 497935 395263 497969 395297
rect 498003 395263 498037 395297
rect 498071 395263 498105 395297
rect 498139 395263 498173 395297
rect 498207 395263 498241 395297
rect 498275 395263 498309 395297
rect 498343 395263 498377 395297
rect 497119 394805 497153 394839
rect 497187 394805 497221 394839
rect 497255 394805 497289 394839
rect 497323 394805 497357 394839
rect 497391 394805 497425 394839
rect 497459 394805 497493 394839
rect 497527 394805 497561 394839
rect 497595 394805 497629 394839
rect 497663 394805 497697 394839
rect 497731 394805 497765 394839
rect 497799 394805 497833 394839
rect 497867 394805 497901 394839
rect 497935 394805 497969 394839
rect 498003 394805 498037 394839
rect 498071 394805 498105 394839
rect 498139 394805 498173 394839
rect 498207 394805 498241 394839
rect 498275 394805 498309 394839
rect 498343 394805 498377 394839
rect 497119 394347 497153 394381
rect 497187 394347 497221 394381
rect 497255 394347 497289 394381
rect 497323 394347 497357 394381
rect 497391 394347 497425 394381
rect 497459 394347 497493 394381
rect 497527 394347 497561 394381
rect 497595 394347 497629 394381
rect 497663 394347 497697 394381
rect 497731 394347 497765 394381
rect 497799 394347 497833 394381
rect 497867 394347 497901 394381
rect 497935 394347 497969 394381
rect 498003 394347 498037 394381
rect 498071 394347 498105 394381
rect 498139 394347 498173 394381
rect 498207 394347 498241 394381
rect 498275 394347 498309 394381
rect 498343 394347 498377 394381
rect 497119 393889 497153 393923
rect 497187 393889 497221 393923
rect 497255 393889 497289 393923
rect 497323 393889 497357 393923
rect 497391 393889 497425 393923
rect 497459 393889 497493 393923
rect 497527 393889 497561 393923
rect 497595 393889 497629 393923
rect 497663 393889 497697 393923
rect 497731 393889 497765 393923
rect 497799 393889 497833 393923
rect 497867 393889 497901 393923
rect 497935 393889 497969 393923
rect 498003 393889 498037 393923
rect 498071 393889 498105 393923
rect 498139 393889 498173 393923
rect 498207 393889 498241 393923
rect 498275 393889 498309 393923
rect 498343 393889 498377 393923
rect 497119 393431 497153 393465
rect 497187 393431 497221 393465
rect 497255 393431 497289 393465
rect 497323 393431 497357 393465
rect 497391 393431 497425 393465
rect 497459 393431 497493 393465
rect 497527 393431 497561 393465
rect 497595 393431 497629 393465
rect 497663 393431 497697 393465
rect 497731 393431 497765 393465
rect 497799 393431 497833 393465
rect 497867 393431 497901 393465
rect 497935 393431 497969 393465
rect 498003 393431 498037 393465
rect 498071 393431 498105 393465
rect 498139 393431 498173 393465
rect 498207 393431 498241 393465
rect 498275 393431 498309 393465
rect 498343 393431 498377 393465
rect 497119 392973 497153 393007
rect 497187 392973 497221 393007
rect 497255 392973 497289 393007
rect 497323 392973 497357 393007
rect 497391 392973 497425 393007
rect 497459 392973 497493 393007
rect 497527 392973 497561 393007
rect 497595 392973 497629 393007
rect 497663 392973 497697 393007
rect 497731 392973 497765 393007
rect 497799 392973 497833 393007
rect 497867 392973 497901 393007
rect 497935 392973 497969 393007
rect 498003 392973 498037 393007
rect 498071 392973 498105 393007
rect 498139 392973 498173 393007
rect 498207 392973 498241 393007
rect 498275 392973 498309 393007
rect 498343 392973 498377 393007
rect 497119 392515 497153 392549
rect 497187 392515 497221 392549
rect 497255 392515 497289 392549
rect 497323 392515 497357 392549
rect 497391 392515 497425 392549
rect 497459 392515 497493 392549
rect 497527 392515 497561 392549
rect 497595 392515 497629 392549
rect 497663 392515 497697 392549
rect 497731 392515 497765 392549
rect 497799 392515 497833 392549
rect 497867 392515 497901 392549
rect 497935 392515 497969 392549
rect 498003 392515 498037 392549
rect 498071 392515 498105 392549
rect 498139 392515 498173 392549
rect 498207 392515 498241 392549
rect 498275 392515 498309 392549
rect 498343 392515 498377 392549
rect 500879 392199 500913 392233
rect 500947 392199 500981 392233
rect 501015 392199 501049 392233
rect 501083 392199 501117 392233
rect 501151 392199 501185 392233
rect 501219 392199 501253 392233
rect 501287 392199 501321 392233
rect 501355 392199 501389 392233
rect 501423 392199 501457 392233
rect 501491 392199 501525 392233
rect 501559 392199 501593 392233
rect 501627 392199 501661 392233
rect 501695 392199 501729 392233
rect 501763 392199 501797 392233
rect 501831 392199 501865 392233
rect 501899 392199 501933 392233
rect 501967 392199 502001 392233
rect 502035 392199 502069 392233
rect 502103 392199 502137 392233
rect 497119 392057 497153 392091
rect 497187 392057 497221 392091
rect 497255 392057 497289 392091
rect 497323 392057 497357 392091
rect 497391 392057 497425 392091
rect 497459 392057 497493 392091
rect 497527 392057 497561 392091
rect 497595 392057 497629 392091
rect 497663 392057 497697 392091
rect 497731 392057 497765 392091
rect 497799 392057 497833 392091
rect 497867 392057 497901 392091
rect 497935 392057 497969 392091
rect 498003 392057 498037 392091
rect 498071 392057 498105 392091
rect 498139 392057 498173 392091
rect 498207 392057 498241 392091
rect 498275 392057 498309 392091
rect 498343 392057 498377 392091
rect 500879 391741 500913 391775
rect 500947 391741 500981 391775
rect 501015 391741 501049 391775
rect 501083 391741 501117 391775
rect 501151 391741 501185 391775
rect 501219 391741 501253 391775
rect 501287 391741 501321 391775
rect 501355 391741 501389 391775
rect 501423 391741 501457 391775
rect 501491 391741 501525 391775
rect 501559 391741 501593 391775
rect 501627 391741 501661 391775
rect 501695 391741 501729 391775
rect 501763 391741 501797 391775
rect 501831 391741 501865 391775
rect 501899 391741 501933 391775
rect 501967 391741 502001 391775
rect 502035 391741 502069 391775
rect 502103 391741 502137 391775
rect 497119 391599 497153 391633
rect 497187 391599 497221 391633
rect 497255 391599 497289 391633
rect 497323 391599 497357 391633
rect 497391 391599 497425 391633
rect 497459 391599 497493 391633
rect 497527 391599 497561 391633
rect 497595 391599 497629 391633
rect 497663 391599 497697 391633
rect 497731 391599 497765 391633
rect 497799 391599 497833 391633
rect 497867 391599 497901 391633
rect 497935 391599 497969 391633
rect 498003 391599 498037 391633
rect 498071 391599 498105 391633
rect 498139 391599 498173 391633
rect 498207 391599 498241 391633
rect 498275 391599 498309 391633
rect 498343 391599 498377 391633
rect 497119 391141 497153 391175
rect 497187 391141 497221 391175
rect 497255 391141 497289 391175
rect 497323 391141 497357 391175
rect 497391 391141 497425 391175
rect 497459 391141 497493 391175
rect 497527 391141 497561 391175
rect 497595 391141 497629 391175
rect 497663 391141 497697 391175
rect 497731 391141 497765 391175
rect 497799 391141 497833 391175
rect 497867 391141 497901 391175
rect 497935 391141 497969 391175
rect 498003 391141 498037 391175
rect 498071 391141 498105 391175
rect 498139 391141 498173 391175
rect 498207 391141 498241 391175
rect 498275 391141 498309 391175
rect 498343 391141 498377 391175
rect 500879 391283 500913 391317
rect 500947 391283 500981 391317
rect 501015 391283 501049 391317
rect 501083 391283 501117 391317
rect 501151 391283 501185 391317
rect 501219 391283 501253 391317
rect 501287 391283 501321 391317
rect 501355 391283 501389 391317
rect 501423 391283 501457 391317
rect 501491 391283 501525 391317
rect 501559 391283 501593 391317
rect 501627 391283 501661 391317
rect 501695 391283 501729 391317
rect 501763 391283 501797 391317
rect 501831 391283 501865 391317
rect 501899 391283 501933 391317
rect 501967 391283 502001 391317
rect 502035 391283 502069 391317
rect 502103 391283 502137 391317
rect 497119 390683 497153 390717
rect 497187 390683 497221 390717
rect 497255 390683 497289 390717
rect 497323 390683 497357 390717
rect 497391 390683 497425 390717
rect 497459 390683 497493 390717
rect 497527 390683 497561 390717
rect 497595 390683 497629 390717
rect 497663 390683 497697 390717
rect 497731 390683 497765 390717
rect 497799 390683 497833 390717
rect 497867 390683 497901 390717
rect 497935 390683 497969 390717
rect 498003 390683 498037 390717
rect 498071 390683 498105 390717
rect 498139 390683 498173 390717
rect 498207 390683 498241 390717
rect 498275 390683 498309 390717
rect 498343 390683 498377 390717
rect 500879 390825 500913 390859
rect 500947 390825 500981 390859
rect 501015 390825 501049 390859
rect 501083 390825 501117 390859
rect 501151 390825 501185 390859
rect 501219 390825 501253 390859
rect 501287 390825 501321 390859
rect 501355 390825 501389 390859
rect 501423 390825 501457 390859
rect 501491 390825 501525 390859
rect 501559 390825 501593 390859
rect 501627 390825 501661 390859
rect 501695 390825 501729 390859
rect 501763 390825 501797 390859
rect 501831 390825 501865 390859
rect 501899 390825 501933 390859
rect 501967 390825 502001 390859
rect 502035 390825 502069 390859
rect 502103 390825 502137 390859
rect 497119 390225 497153 390259
rect 497187 390225 497221 390259
rect 497255 390225 497289 390259
rect 497323 390225 497357 390259
rect 497391 390225 497425 390259
rect 497459 390225 497493 390259
rect 497527 390225 497561 390259
rect 497595 390225 497629 390259
rect 497663 390225 497697 390259
rect 497731 390225 497765 390259
rect 497799 390225 497833 390259
rect 497867 390225 497901 390259
rect 497935 390225 497969 390259
rect 498003 390225 498037 390259
rect 498071 390225 498105 390259
rect 498139 390225 498173 390259
rect 498207 390225 498241 390259
rect 498275 390225 498309 390259
rect 498343 390225 498377 390259
rect 493359 390043 493393 390077
rect 493427 390043 493461 390077
rect 493495 390043 493529 390077
rect 493563 390043 493597 390077
rect 493631 390043 493665 390077
rect 493699 390043 493733 390077
rect 493767 390043 493801 390077
rect 493835 390043 493869 390077
rect 493903 390043 493937 390077
rect 493971 390043 494005 390077
rect 494039 390043 494073 390077
rect 494107 390043 494141 390077
rect 494175 390043 494209 390077
rect 494243 390043 494277 390077
rect 494311 390043 494345 390077
rect 494379 390043 494413 390077
rect 494447 390043 494481 390077
rect 494515 390043 494549 390077
rect 494583 390043 494617 390077
rect 493359 389585 493393 389619
rect 493427 389585 493461 389619
rect 493495 389585 493529 389619
rect 493563 389585 493597 389619
rect 493631 389585 493665 389619
rect 493699 389585 493733 389619
rect 493767 389585 493801 389619
rect 493835 389585 493869 389619
rect 493903 389585 493937 389619
rect 493971 389585 494005 389619
rect 494039 389585 494073 389619
rect 494107 389585 494141 389619
rect 494175 389585 494209 389619
rect 494243 389585 494277 389619
rect 494311 389585 494345 389619
rect 494379 389585 494413 389619
rect 494447 389585 494481 389619
rect 494515 389585 494549 389619
rect 494583 389585 494617 389619
rect 500879 390367 500913 390401
rect 500947 390367 500981 390401
rect 501015 390367 501049 390401
rect 501083 390367 501117 390401
rect 501151 390367 501185 390401
rect 501219 390367 501253 390401
rect 501287 390367 501321 390401
rect 501355 390367 501389 390401
rect 501423 390367 501457 390401
rect 501491 390367 501525 390401
rect 501559 390367 501593 390401
rect 501627 390367 501661 390401
rect 501695 390367 501729 390401
rect 501763 390367 501797 390401
rect 501831 390367 501865 390401
rect 501899 390367 501933 390401
rect 501967 390367 502001 390401
rect 502035 390367 502069 390401
rect 502103 390367 502137 390401
rect 497119 389767 497153 389801
rect 497187 389767 497221 389801
rect 497255 389767 497289 389801
rect 497323 389767 497357 389801
rect 497391 389767 497425 389801
rect 497459 389767 497493 389801
rect 497527 389767 497561 389801
rect 497595 389767 497629 389801
rect 497663 389767 497697 389801
rect 497731 389767 497765 389801
rect 497799 389767 497833 389801
rect 497867 389767 497901 389801
rect 497935 389767 497969 389801
rect 498003 389767 498037 389801
rect 498071 389767 498105 389801
rect 498139 389767 498173 389801
rect 498207 389767 498241 389801
rect 498275 389767 498309 389801
rect 498343 389767 498377 389801
rect 500879 389909 500913 389943
rect 500947 389909 500981 389943
rect 501015 389909 501049 389943
rect 501083 389909 501117 389943
rect 501151 389909 501185 389943
rect 501219 389909 501253 389943
rect 501287 389909 501321 389943
rect 501355 389909 501389 389943
rect 501423 389909 501457 389943
rect 501491 389909 501525 389943
rect 501559 389909 501593 389943
rect 501627 389909 501661 389943
rect 501695 389909 501729 389943
rect 501763 389909 501797 389943
rect 501831 389909 501865 389943
rect 501899 389909 501933 389943
rect 501967 389909 502001 389943
rect 502035 389909 502069 389943
rect 502103 389909 502137 389943
rect 493359 389127 493393 389161
rect 493427 389127 493461 389161
rect 493495 389127 493529 389161
rect 493563 389127 493597 389161
rect 493631 389127 493665 389161
rect 493699 389127 493733 389161
rect 493767 389127 493801 389161
rect 493835 389127 493869 389161
rect 493903 389127 493937 389161
rect 493971 389127 494005 389161
rect 494039 389127 494073 389161
rect 494107 389127 494141 389161
rect 494175 389127 494209 389161
rect 494243 389127 494277 389161
rect 494311 389127 494345 389161
rect 494379 389127 494413 389161
rect 494447 389127 494481 389161
rect 494515 389127 494549 389161
rect 494583 389127 494617 389161
rect 497119 389309 497153 389343
rect 497187 389309 497221 389343
rect 497255 389309 497289 389343
rect 497323 389309 497357 389343
rect 497391 389309 497425 389343
rect 497459 389309 497493 389343
rect 497527 389309 497561 389343
rect 497595 389309 497629 389343
rect 497663 389309 497697 389343
rect 497731 389309 497765 389343
rect 497799 389309 497833 389343
rect 497867 389309 497901 389343
rect 497935 389309 497969 389343
rect 498003 389309 498037 389343
rect 498071 389309 498105 389343
rect 498139 389309 498173 389343
rect 498207 389309 498241 389343
rect 498275 389309 498309 389343
rect 498343 389309 498377 389343
rect 500879 389451 500913 389485
rect 500947 389451 500981 389485
rect 501015 389451 501049 389485
rect 501083 389451 501117 389485
rect 501151 389451 501185 389485
rect 501219 389451 501253 389485
rect 501287 389451 501321 389485
rect 501355 389451 501389 389485
rect 501423 389451 501457 389485
rect 501491 389451 501525 389485
rect 501559 389451 501593 389485
rect 501627 389451 501661 389485
rect 501695 389451 501729 389485
rect 501763 389451 501797 389485
rect 501831 389451 501865 389485
rect 501899 389451 501933 389485
rect 501967 389451 502001 389485
rect 502035 389451 502069 389485
rect 502103 389451 502137 389485
rect 500879 388993 500913 389027
rect 500947 388993 500981 389027
rect 501015 388993 501049 389027
rect 501083 388993 501117 389027
rect 501151 388993 501185 389027
rect 501219 388993 501253 389027
rect 501287 388993 501321 389027
rect 501355 388993 501389 389027
rect 501423 388993 501457 389027
rect 501491 388993 501525 389027
rect 501559 388993 501593 389027
rect 501627 388993 501661 389027
rect 501695 388993 501729 389027
rect 501763 388993 501797 389027
rect 501831 388993 501865 389027
rect 501899 388993 501933 389027
rect 501967 388993 502001 389027
rect 502035 388993 502069 389027
rect 502103 388993 502137 389027
rect 497119 388851 497153 388885
rect 497187 388851 497221 388885
rect 497255 388851 497289 388885
rect 497323 388851 497357 388885
rect 497391 388851 497425 388885
rect 497459 388851 497493 388885
rect 497527 388851 497561 388885
rect 497595 388851 497629 388885
rect 497663 388851 497697 388885
rect 497731 388851 497765 388885
rect 497799 388851 497833 388885
rect 497867 388851 497901 388885
rect 497935 388851 497969 388885
rect 498003 388851 498037 388885
rect 498071 388851 498105 388885
rect 498139 388851 498173 388885
rect 498207 388851 498241 388885
rect 498275 388851 498309 388885
rect 498343 388851 498377 388885
rect 493359 388669 493393 388703
rect 493427 388669 493461 388703
rect 493495 388669 493529 388703
rect 493563 388669 493597 388703
rect 493631 388669 493665 388703
rect 493699 388669 493733 388703
rect 493767 388669 493801 388703
rect 493835 388669 493869 388703
rect 493903 388669 493937 388703
rect 493971 388669 494005 388703
rect 494039 388669 494073 388703
rect 494107 388669 494141 388703
rect 494175 388669 494209 388703
rect 494243 388669 494277 388703
rect 494311 388669 494345 388703
rect 494379 388669 494413 388703
rect 494447 388669 494481 388703
rect 494515 388669 494549 388703
rect 494583 388669 494617 388703
rect 500879 388535 500913 388569
rect 500947 388535 500981 388569
rect 501015 388535 501049 388569
rect 501083 388535 501117 388569
rect 501151 388535 501185 388569
rect 501219 388535 501253 388569
rect 501287 388535 501321 388569
rect 501355 388535 501389 388569
rect 501423 388535 501457 388569
rect 501491 388535 501525 388569
rect 501559 388535 501593 388569
rect 501627 388535 501661 388569
rect 501695 388535 501729 388569
rect 501763 388535 501797 388569
rect 501831 388535 501865 388569
rect 501899 388535 501933 388569
rect 501967 388535 502001 388569
rect 502035 388535 502069 388569
rect 502103 388535 502137 388569
rect 497119 388393 497153 388427
rect 497187 388393 497221 388427
rect 497255 388393 497289 388427
rect 497323 388393 497357 388427
rect 497391 388393 497425 388427
rect 497459 388393 497493 388427
rect 497527 388393 497561 388427
rect 497595 388393 497629 388427
rect 497663 388393 497697 388427
rect 497731 388393 497765 388427
rect 497799 388393 497833 388427
rect 497867 388393 497901 388427
rect 497935 388393 497969 388427
rect 498003 388393 498037 388427
rect 498071 388393 498105 388427
rect 498139 388393 498173 388427
rect 498207 388393 498241 388427
rect 498275 388393 498309 388427
rect 498343 388393 498377 388427
rect 493359 388211 493393 388245
rect 493427 388211 493461 388245
rect 493495 388211 493529 388245
rect 493563 388211 493597 388245
rect 493631 388211 493665 388245
rect 493699 388211 493733 388245
rect 493767 388211 493801 388245
rect 493835 388211 493869 388245
rect 493903 388211 493937 388245
rect 493971 388211 494005 388245
rect 494039 388211 494073 388245
rect 494107 388211 494141 388245
rect 494175 388211 494209 388245
rect 494243 388211 494277 388245
rect 494311 388211 494345 388245
rect 494379 388211 494413 388245
rect 494447 388211 494481 388245
rect 494515 388211 494549 388245
rect 494583 388211 494617 388245
rect 497119 387935 497153 387969
rect 497187 387935 497221 387969
rect 497255 387935 497289 387969
rect 497323 387935 497357 387969
rect 497391 387935 497425 387969
rect 497459 387935 497493 387969
rect 497527 387935 497561 387969
rect 497595 387935 497629 387969
rect 497663 387935 497697 387969
rect 497731 387935 497765 387969
rect 497799 387935 497833 387969
rect 497867 387935 497901 387969
rect 497935 387935 497969 387969
rect 498003 387935 498037 387969
rect 498071 387935 498105 387969
rect 498139 387935 498173 387969
rect 498207 387935 498241 387969
rect 498275 387935 498309 387969
rect 498343 387935 498377 387969
rect 493359 387753 493393 387787
rect 493427 387753 493461 387787
rect 493495 387753 493529 387787
rect 493563 387753 493597 387787
rect 493631 387753 493665 387787
rect 493699 387753 493733 387787
rect 493767 387753 493801 387787
rect 493835 387753 493869 387787
rect 493903 387753 493937 387787
rect 493971 387753 494005 387787
rect 494039 387753 494073 387787
rect 494107 387753 494141 387787
rect 494175 387753 494209 387787
rect 494243 387753 494277 387787
rect 494311 387753 494345 387787
rect 494379 387753 494413 387787
rect 494447 387753 494481 387787
rect 494515 387753 494549 387787
rect 494583 387753 494617 387787
rect 500879 388077 500913 388111
rect 500947 388077 500981 388111
rect 501015 388077 501049 388111
rect 501083 388077 501117 388111
rect 501151 388077 501185 388111
rect 501219 388077 501253 388111
rect 501287 388077 501321 388111
rect 501355 388077 501389 388111
rect 501423 388077 501457 388111
rect 501491 388077 501525 388111
rect 501559 388077 501593 388111
rect 501627 388077 501661 388111
rect 501695 388077 501729 388111
rect 501763 388077 501797 388111
rect 501831 388077 501865 388111
rect 501899 388077 501933 388111
rect 501967 388077 502001 388111
rect 502035 388077 502069 388111
rect 502103 388077 502137 388111
rect 523439 390043 523473 390077
rect 523507 390043 523541 390077
rect 523575 390043 523609 390077
rect 523643 390043 523677 390077
rect 523711 390043 523745 390077
rect 523779 390043 523813 390077
rect 523847 390043 523881 390077
rect 523915 390043 523949 390077
rect 523983 390043 524017 390077
rect 524051 390043 524085 390077
rect 524119 390043 524153 390077
rect 524187 390043 524221 390077
rect 524255 390043 524289 390077
rect 524323 390043 524357 390077
rect 524391 390043 524425 390077
rect 524459 390043 524493 390077
rect 524527 390043 524561 390077
rect 524595 390043 524629 390077
rect 524663 390043 524697 390077
rect 523439 389585 523473 389619
rect 523507 389585 523541 389619
rect 523575 389585 523609 389619
rect 523643 389585 523677 389619
rect 523711 389585 523745 389619
rect 523779 389585 523813 389619
rect 523847 389585 523881 389619
rect 523915 389585 523949 389619
rect 523983 389585 524017 389619
rect 524051 389585 524085 389619
rect 524119 389585 524153 389619
rect 524187 389585 524221 389619
rect 524255 389585 524289 389619
rect 524323 389585 524357 389619
rect 524391 389585 524425 389619
rect 524459 389585 524493 389619
rect 524527 389585 524561 389619
rect 524595 389585 524629 389619
rect 524663 389585 524697 389619
rect 523439 389127 523473 389161
rect 523507 389127 523541 389161
rect 523575 389127 523609 389161
rect 523643 389127 523677 389161
rect 523711 389127 523745 389161
rect 523779 389127 523813 389161
rect 523847 389127 523881 389161
rect 523915 389127 523949 389161
rect 523983 389127 524017 389161
rect 524051 389127 524085 389161
rect 524119 389127 524153 389161
rect 524187 389127 524221 389161
rect 524255 389127 524289 389161
rect 524323 389127 524357 389161
rect 524391 389127 524425 389161
rect 524459 389127 524493 389161
rect 524527 389127 524561 389161
rect 524595 389127 524629 389161
rect 524663 389127 524697 389161
rect 523439 388669 523473 388703
rect 523507 388669 523541 388703
rect 523575 388669 523609 388703
rect 523643 388669 523677 388703
rect 523711 388669 523745 388703
rect 523779 388669 523813 388703
rect 523847 388669 523881 388703
rect 523915 388669 523949 388703
rect 523983 388669 524017 388703
rect 524051 388669 524085 388703
rect 524119 388669 524153 388703
rect 524187 388669 524221 388703
rect 524255 388669 524289 388703
rect 524323 388669 524357 388703
rect 524391 388669 524425 388703
rect 524459 388669 524493 388703
rect 524527 388669 524561 388703
rect 524595 388669 524629 388703
rect 524663 388669 524697 388703
rect 493359 387295 493393 387329
rect 493427 387295 493461 387329
rect 493495 387295 493529 387329
rect 493563 387295 493597 387329
rect 493631 387295 493665 387329
rect 493699 387295 493733 387329
rect 493767 387295 493801 387329
rect 493835 387295 493869 387329
rect 493903 387295 493937 387329
rect 493971 387295 494005 387329
rect 494039 387295 494073 387329
rect 494107 387295 494141 387329
rect 494175 387295 494209 387329
rect 494243 387295 494277 387329
rect 494311 387295 494345 387329
rect 494379 387295 494413 387329
rect 494447 387295 494481 387329
rect 494515 387295 494549 387329
rect 494583 387295 494617 387329
rect 497119 387477 497153 387511
rect 497187 387477 497221 387511
rect 497255 387477 497289 387511
rect 497323 387477 497357 387511
rect 497391 387477 497425 387511
rect 497459 387477 497493 387511
rect 497527 387477 497561 387511
rect 497595 387477 497629 387511
rect 497663 387477 497697 387511
rect 497731 387477 497765 387511
rect 497799 387477 497833 387511
rect 497867 387477 497901 387511
rect 497935 387477 497969 387511
rect 498003 387477 498037 387511
rect 498071 387477 498105 387511
rect 498139 387477 498173 387511
rect 498207 387477 498241 387511
rect 498275 387477 498309 387511
rect 498343 387477 498377 387511
rect 523439 388211 523473 388245
rect 523507 388211 523541 388245
rect 523575 388211 523609 388245
rect 523643 388211 523677 388245
rect 523711 388211 523745 388245
rect 523779 388211 523813 388245
rect 523847 388211 523881 388245
rect 523915 388211 523949 388245
rect 523983 388211 524017 388245
rect 524051 388211 524085 388245
rect 524119 388211 524153 388245
rect 524187 388211 524221 388245
rect 524255 388211 524289 388245
rect 524323 388211 524357 388245
rect 524391 388211 524425 388245
rect 524459 388211 524493 388245
rect 524527 388211 524561 388245
rect 524595 388211 524629 388245
rect 524663 388211 524697 388245
rect 500879 387619 500913 387653
rect 500947 387619 500981 387653
rect 501015 387619 501049 387653
rect 501083 387619 501117 387653
rect 501151 387619 501185 387653
rect 501219 387619 501253 387653
rect 501287 387619 501321 387653
rect 501355 387619 501389 387653
rect 501423 387619 501457 387653
rect 501491 387619 501525 387653
rect 501559 387619 501593 387653
rect 501627 387619 501661 387653
rect 501695 387619 501729 387653
rect 501763 387619 501797 387653
rect 501831 387619 501865 387653
rect 501899 387619 501933 387653
rect 501967 387619 502001 387653
rect 502035 387619 502069 387653
rect 502103 387619 502137 387653
rect 493359 386837 493393 386871
rect 493427 386837 493461 386871
rect 493495 386837 493529 386871
rect 493563 386837 493597 386871
rect 493631 386837 493665 386871
rect 493699 386837 493733 386871
rect 493767 386837 493801 386871
rect 493835 386837 493869 386871
rect 493903 386837 493937 386871
rect 493971 386837 494005 386871
rect 494039 386837 494073 386871
rect 494107 386837 494141 386871
rect 494175 386837 494209 386871
rect 494243 386837 494277 386871
rect 494311 386837 494345 386871
rect 494379 386837 494413 386871
rect 494447 386837 494481 386871
rect 494515 386837 494549 386871
rect 494583 386837 494617 386871
rect 497119 387019 497153 387053
rect 497187 387019 497221 387053
rect 497255 387019 497289 387053
rect 497323 387019 497357 387053
rect 497391 387019 497425 387053
rect 497459 387019 497493 387053
rect 497527 387019 497561 387053
rect 497595 387019 497629 387053
rect 497663 387019 497697 387053
rect 497731 387019 497765 387053
rect 497799 387019 497833 387053
rect 497867 387019 497901 387053
rect 497935 387019 497969 387053
rect 498003 387019 498037 387053
rect 498071 387019 498105 387053
rect 498139 387019 498173 387053
rect 498207 387019 498241 387053
rect 498275 387019 498309 387053
rect 498343 387019 498377 387053
rect 500879 387161 500913 387195
rect 500947 387161 500981 387195
rect 501015 387161 501049 387195
rect 501083 387161 501117 387195
rect 501151 387161 501185 387195
rect 501219 387161 501253 387195
rect 501287 387161 501321 387195
rect 501355 387161 501389 387195
rect 501423 387161 501457 387195
rect 501491 387161 501525 387195
rect 501559 387161 501593 387195
rect 501627 387161 501661 387195
rect 501695 387161 501729 387195
rect 501763 387161 501797 387195
rect 501831 387161 501865 387195
rect 501899 387161 501933 387195
rect 501967 387161 502001 387195
rect 502035 387161 502069 387195
rect 502103 387161 502137 387195
rect 493359 386379 493393 386413
rect 493427 386379 493461 386413
rect 493495 386379 493529 386413
rect 493563 386379 493597 386413
rect 493631 386379 493665 386413
rect 493699 386379 493733 386413
rect 493767 386379 493801 386413
rect 493835 386379 493869 386413
rect 493903 386379 493937 386413
rect 493971 386379 494005 386413
rect 494039 386379 494073 386413
rect 494107 386379 494141 386413
rect 494175 386379 494209 386413
rect 494243 386379 494277 386413
rect 494311 386379 494345 386413
rect 494379 386379 494413 386413
rect 494447 386379 494481 386413
rect 494515 386379 494549 386413
rect 494583 386379 494617 386413
rect 497119 386561 497153 386595
rect 497187 386561 497221 386595
rect 497255 386561 497289 386595
rect 497323 386561 497357 386595
rect 497391 386561 497425 386595
rect 497459 386561 497493 386595
rect 497527 386561 497561 386595
rect 497595 386561 497629 386595
rect 497663 386561 497697 386595
rect 497731 386561 497765 386595
rect 497799 386561 497833 386595
rect 497867 386561 497901 386595
rect 497935 386561 497969 386595
rect 498003 386561 498037 386595
rect 498071 386561 498105 386595
rect 498139 386561 498173 386595
rect 498207 386561 498241 386595
rect 498275 386561 498309 386595
rect 498343 386561 498377 386595
rect 500879 386703 500913 386737
rect 500947 386703 500981 386737
rect 501015 386703 501049 386737
rect 501083 386703 501117 386737
rect 501151 386703 501185 386737
rect 501219 386703 501253 386737
rect 501287 386703 501321 386737
rect 501355 386703 501389 386737
rect 501423 386703 501457 386737
rect 501491 386703 501525 386737
rect 501559 386703 501593 386737
rect 501627 386703 501661 386737
rect 501695 386703 501729 386737
rect 501763 386703 501797 386737
rect 501831 386703 501865 386737
rect 501899 386703 501933 386737
rect 501967 386703 502001 386737
rect 502035 386703 502069 386737
rect 502103 386703 502137 386737
rect 493359 385921 493393 385955
rect 493427 385921 493461 385955
rect 493495 385921 493529 385955
rect 493563 385921 493597 385955
rect 493631 385921 493665 385955
rect 493699 385921 493733 385955
rect 493767 385921 493801 385955
rect 493835 385921 493869 385955
rect 493903 385921 493937 385955
rect 493971 385921 494005 385955
rect 494039 385921 494073 385955
rect 494107 385921 494141 385955
rect 494175 385921 494209 385955
rect 494243 385921 494277 385955
rect 494311 385921 494345 385955
rect 494379 385921 494413 385955
rect 494447 385921 494481 385955
rect 494515 385921 494549 385955
rect 494583 385921 494617 385955
rect 497119 386103 497153 386137
rect 497187 386103 497221 386137
rect 497255 386103 497289 386137
rect 497323 386103 497357 386137
rect 497391 386103 497425 386137
rect 497459 386103 497493 386137
rect 497527 386103 497561 386137
rect 497595 386103 497629 386137
rect 497663 386103 497697 386137
rect 497731 386103 497765 386137
rect 497799 386103 497833 386137
rect 497867 386103 497901 386137
rect 497935 386103 497969 386137
rect 498003 386103 498037 386137
rect 498071 386103 498105 386137
rect 498139 386103 498173 386137
rect 498207 386103 498241 386137
rect 498275 386103 498309 386137
rect 498343 386103 498377 386137
rect 497119 385645 497153 385679
rect 497187 385645 497221 385679
rect 497255 385645 497289 385679
rect 497323 385645 497357 385679
rect 497391 385645 497425 385679
rect 497459 385645 497493 385679
rect 497527 385645 497561 385679
rect 497595 385645 497629 385679
rect 497663 385645 497697 385679
rect 497731 385645 497765 385679
rect 497799 385645 497833 385679
rect 497867 385645 497901 385679
rect 497935 385645 497969 385679
rect 498003 385645 498037 385679
rect 498071 385645 498105 385679
rect 498139 385645 498173 385679
rect 498207 385645 498241 385679
rect 498275 385645 498309 385679
rect 498343 385645 498377 385679
rect 493359 385463 493393 385497
rect 493427 385463 493461 385497
rect 493495 385463 493529 385497
rect 493563 385463 493597 385497
rect 493631 385463 493665 385497
rect 493699 385463 493733 385497
rect 493767 385463 493801 385497
rect 493835 385463 493869 385497
rect 493903 385463 493937 385497
rect 493971 385463 494005 385497
rect 494039 385463 494073 385497
rect 494107 385463 494141 385497
rect 494175 385463 494209 385497
rect 494243 385463 494277 385497
rect 494311 385463 494345 385497
rect 494379 385463 494413 385497
rect 494447 385463 494481 385497
rect 494515 385463 494549 385497
rect 494583 385463 494617 385497
rect 500879 385535 500913 385569
rect 500947 385535 500981 385569
rect 501015 385535 501049 385569
rect 501083 385535 501117 385569
rect 501151 385535 501185 385569
rect 501219 385535 501253 385569
rect 501287 385535 501321 385569
rect 501355 385535 501389 385569
rect 501423 385535 501457 385569
rect 501491 385535 501525 385569
rect 501559 385535 501593 385569
rect 501627 385535 501661 385569
rect 501695 385535 501729 385569
rect 501763 385535 501797 385569
rect 501831 385535 501865 385569
rect 501899 385535 501933 385569
rect 501967 385535 502001 385569
rect 502035 385535 502069 385569
rect 502103 385535 502137 385569
rect 497119 385187 497153 385221
rect 497187 385187 497221 385221
rect 497255 385187 497289 385221
rect 497323 385187 497357 385221
rect 497391 385187 497425 385221
rect 497459 385187 497493 385221
rect 497527 385187 497561 385221
rect 497595 385187 497629 385221
rect 497663 385187 497697 385221
rect 497731 385187 497765 385221
rect 497799 385187 497833 385221
rect 497867 385187 497901 385221
rect 497935 385187 497969 385221
rect 498003 385187 498037 385221
rect 498071 385187 498105 385221
rect 498139 385187 498173 385221
rect 498207 385187 498241 385221
rect 498275 385187 498309 385221
rect 498343 385187 498377 385221
rect 493359 385005 493393 385039
rect 493427 385005 493461 385039
rect 493495 385005 493529 385039
rect 493563 385005 493597 385039
rect 493631 385005 493665 385039
rect 493699 385005 493733 385039
rect 493767 385005 493801 385039
rect 493835 385005 493869 385039
rect 493903 385005 493937 385039
rect 493971 385005 494005 385039
rect 494039 385005 494073 385039
rect 494107 385005 494141 385039
rect 494175 385005 494209 385039
rect 494243 385005 494277 385039
rect 494311 385005 494345 385039
rect 494379 385005 494413 385039
rect 494447 385005 494481 385039
rect 494515 385005 494549 385039
rect 494583 385005 494617 385039
rect 523439 387753 523473 387787
rect 523507 387753 523541 387787
rect 523575 387753 523609 387787
rect 523643 387753 523677 387787
rect 523711 387753 523745 387787
rect 523779 387753 523813 387787
rect 523847 387753 523881 387787
rect 523915 387753 523949 387787
rect 523983 387753 524017 387787
rect 524051 387753 524085 387787
rect 524119 387753 524153 387787
rect 524187 387753 524221 387787
rect 524255 387753 524289 387787
rect 524323 387753 524357 387787
rect 524391 387753 524425 387787
rect 524459 387753 524493 387787
rect 524527 387753 524561 387787
rect 524595 387753 524629 387787
rect 524663 387753 524697 387787
rect 523439 387295 523473 387329
rect 523507 387295 523541 387329
rect 523575 387295 523609 387329
rect 523643 387295 523677 387329
rect 523711 387295 523745 387329
rect 523779 387295 523813 387329
rect 523847 387295 523881 387329
rect 523915 387295 523949 387329
rect 523983 387295 524017 387329
rect 524051 387295 524085 387329
rect 524119 387295 524153 387329
rect 524187 387295 524221 387329
rect 524255 387295 524289 387329
rect 524323 387295 524357 387329
rect 524391 387295 524425 387329
rect 524459 387295 524493 387329
rect 524527 387295 524561 387329
rect 524595 387295 524629 387329
rect 524663 387295 524697 387329
rect 523439 386837 523473 386871
rect 523507 386837 523541 386871
rect 523575 386837 523609 386871
rect 523643 386837 523677 386871
rect 523711 386837 523745 386871
rect 523779 386837 523813 386871
rect 523847 386837 523881 386871
rect 523915 386837 523949 386871
rect 523983 386837 524017 386871
rect 524051 386837 524085 386871
rect 524119 386837 524153 386871
rect 524187 386837 524221 386871
rect 524255 386837 524289 386871
rect 524323 386837 524357 386871
rect 524391 386837 524425 386871
rect 524459 386837 524493 386871
rect 524527 386837 524561 386871
rect 524595 386837 524629 386871
rect 524663 386837 524697 386871
rect 523439 386379 523473 386413
rect 523507 386379 523541 386413
rect 523575 386379 523609 386413
rect 523643 386379 523677 386413
rect 523711 386379 523745 386413
rect 523779 386379 523813 386413
rect 523847 386379 523881 386413
rect 523915 386379 523949 386413
rect 523983 386379 524017 386413
rect 524051 386379 524085 386413
rect 524119 386379 524153 386413
rect 524187 386379 524221 386413
rect 524255 386379 524289 386413
rect 524323 386379 524357 386413
rect 524391 386379 524425 386413
rect 524459 386379 524493 386413
rect 524527 386379 524561 386413
rect 524595 386379 524629 386413
rect 524663 386379 524697 386413
rect 523439 385921 523473 385955
rect 523507 385921 523541 385955
rect 523575 385921 523609 385955
rect 523643 385921 523677 385955
rect 523711 385921 523745 385955
rect 523779 385921 523813 385955
rect 523847 385921 523881 385955
rect 523915 385921 523949 385955
rect 523983 385921 524017 385955
rect 524051 385921 524085 385955
rect 524119 385921 524153 385955
rect 524187 385921 524221 385955
rect 524255 385921 524289 385955
rect 524323 385921 524357 385955
rect 524391 385921 524425 385955
rect 524459 385921 524493 385955
rect 524527 385921 524561 385955
rect 524595 385921 524629 385955
rect 524663 385921 524697 385955
rect 523439 385463 523473 385497
rect 523507 385463 523541 385497
rect 523575 385463 523609 385497
rect 523643 385463 523677 385497
rect 523711 385463 523745 385497
rect 523779 385463 523813 385497
rect 523847 385463 523881 385497
rect 523915 385463 523949 385497
rect 523983 385463 524017 385497
rect 524051 385463 524085 385497
rect 524119 385463 524153 385497
rect 524187 385463 524221 385497
rect 524255 385463 524289 385497
rect 524323 385463 524357 385497
rect 524391 385463 524425 385497
rect 524459 385463 524493 385497
rect 524527 385463 524561 385497
rect 524595 385463 524629 385497
rect 524663 385463 524697 385497
rect 500879 385077 500913 385111
rect 500947 385077 500981 385111
rect 501015 385077 501049 385111
rect 501083 385077 501117 385111
rect 501151 385077 501185 385111
rect 501219 385077 501253 385111
rect 501287 385077 501321 385111
rect 501355 385077 501389 385111
rect 501423 385077 501457 385111
rect 501491 385077 501525 385111
rect 501559 385077 501593 385111
rect 501627 385077 501661 385111
rect 501695 385077 501729 385111
rect 501763 385077 501797 385111
rect 501831 385077 501865 385111
rect 501899 385077 501933 385111
rect 501967 385077 502001 385111
rect 502035 385077 502069 385111
rect 502103 385077 502137 385111
rect 497119 384729 497153 384763
rect 497187 384729 497221 384763
rect 497255 384729 497289 384763
rect 497323 384729 497357 384763
rect 497391 384729 497425 384763
rect 497459 384729 497493 384763
rect 497527 384729 497561 384763
rect 497595 384729 497629 384763
rect 497663 384729 497697 384763
rect 497731 384729 497765 384763
rect 497799 384729 497833 384763
rect 497867 384729 497901 384763
rect 497935 384729 497969 384763
rect 498003 384729 498037 384763
rect 498071 384729 498105 384763
rect 498139 384729 498173 384763
rect 498207 384729 498241 384763
rect 498275 384729 498309 384763
rect 498343 384729 498377 384763
rect 493359 384547 493393 384581
rect 493427 384547 493461 384581
rect 493495 384547 493529 384581
rect 493563 384547 493597 384581
rect 493631 384547 493665 384581
rect 493699 384547 493733 384581
rect 493767 384547 493801 384581
rect 493835 384547 493869 384581
rect 493903 384547 493937 384581
rect 493971 384547 494005 384581
rect 494039 384547 494073 384581
rect 494107 384547 494141 384581
rect 494175 384547 494209 384581
rect 494243 384547 494277 384581
rect 494311 384547 494345 384581
rect 494379 384547 494413 384581
rect 494447 384547 494481 384581
rect 494515 384547 494549 384581
rect 494583 384547 494617 384581
rect 500879 384619 500913 384653
rect 500947 384619 500981 384653
rect 501015 384619 501049 384653
rect 501083 384619 501117 384653
rect 501151 384619 501185 384653
rect 501219 384619 501253 384653
rect 501287 384619 501321 384653
rect 501355 384619 501389 384653
rect 501423 384619 501457 384653
rect 501491 384619 501525 384653
rect 501559 384619 501593 384653
rect 501627 384619 501661 384653
rect 501695 384619 501729 384653
rect 501763 384619 501797 384653
rect 501831 384619 501865 384653
rect 501899 384619 501933 384653
rect 501967 384619 502001 384653
rect 502035 384619 502069 384653
rect 502103 384619 502137 384653
rect 493359 384089 493393 384123
rect 493427 384089 493461 384123
rect 493495 384089 493529 384123
rect 493563 384089 493597 384123
rect 493631 384089 493665 384123
rect 493699 384089 493733 384123
rect 493767 384089 493801 384123
rect 493835 384089 493869 384123
rect 493903 384089 493937 384123
rect 493971 384089 494005 384123
rect 494039 384089 494073 384123
rect 494107 384089 494141 384123
rect 494175 384089 494209 384123
rect 494243 384089 494277 384123
rect 494311 384089 494345 384123
rect 494379 384089 494413 384123
rect 494447 384089 494481 384123
rect 494515 384089 494549 384123
rect 494583 384089 494617 384123
rect 497119 384271 497153 384305
rect 497187 384271 497221 384305
rect 497255 384271 497289 384305
rect 497323 384271 497357 384305
rect 497391 384271 497425 384305
rect 497459 384271 497493 384305
rect 497527 384271 497561 384305
rect 497595 384271 497629 384305
rect 497663 384271 497697 384305
rect 497731 384271 497765 384305
rect 497799 384271 497833 384305
rect 497867 384271 497901 384305
rect 497935 384271 497969 384305
rect 498003 384271 498037 384305
rect 498071 384271 498105 384305
rect 498139 384271 498173 384305
rect 498207 384271 498241 384305
rect 498275 384271 498309 384305
rect 498343 384271 498377 384305
rect 500879 384161 500913 384195
rect 500947 384161 500981 384195
rect 501015 384161 501049 384195
rect 501083 384161 501117 384195
rect 501151 384161 501185 384195
rect 501219 384161 501253 384195
rect 501287 384161 501321 384195
rect 501355 384161 501389 384195
rect 501423 384161 501457 384195
rect 501491 384161 501525 384195
rect 501559 384161 501593 384195
rect 501627 384161 501661 384195
rect 501695 384161 501729 384195
rect 501763 384161 501797 384195
rect 501831 384161 501865 384195
rect 501899 384161 501933 384195
rect 501967 384161 502001 384195
rect 502035 384161 502069 384195
rect 502103 384161 502137 384195
rect 493359 383631 493393 383665
rect 493427 383631 493461 383665
rect 493495 383631 493529 383665
rect 493563 383631 493597 383665
rect 493631 383631 493665 383665
rect 493699 383631 493733 383665
rect 493767 383631 493801 383665
rect 493835 383631 493869 383665
rect 493903 383631 493937 383665
rect 493971 383631 494005 383665
rect 494039 383631 494073 383665
rect 494107 383631 494141 383665
rect 494175 383631 494209 383665
rect 494243 383631 494277 383665
rect 494311 383631 494345 383665
rect 494379 383631 494413 383665
rect 494447 383631 494481 383665
rect 494515 383631 494549 383665
rect 494583 383631 494617 383665
rect 497119 383813 497153 383847
rect 497187 383813 497221 383847
rect 497255 383813 497289 383847
rect 497323 383813 497357 383847
rect 497391 383813 497425 383847
rect 497459 383813 497493 383847
rect 497527 383813 497561 383847
rect 497595 383813 497629 383847
rect 497663 383813 497697 383847
rect 497731 383813 497765 383847
rect 497799 383813 497833 383847
rect 497867 383813 497901 383847
rect 497935 383813 497969 383847
rect 498003 383813 498037 383847
rect 498071 383813 498105 383847
rect 498139 383813 498173 383847
rect 498207 383813 498241 383847
rect 498275 383813 498309 383847
rect 498343 383813 498377 383847
rect 500879 383703 500913 383737
rect 500947 383703 500981 383737
rect 501015 383703 501049 383737
rect 501083 383703 501117 383737
rect 501151 383703 501185 383737
rect 501219 383703 501253 383737
rect 501287 383703 501321 383737
rect 501355 383703 501389 383737
rect 501423 383703 501457 383737
rect 501491 383703 501525 383737
rect 501559 383703 501593 383737
rect 501627 383703 501661 383737
rect 501695 383703 501729 383737
rect 501763 383703 501797 383737
rect 501831 383703 501865 383737
rect 501899 383703 501933 383737
rect 501967 383703 502001 383737
rect 502035 383703 502069 383737
rect 502103 383703 502137 383737
rect 493359 383173 493393 383207
rect 493427 383173 493461 383207
rect 493495 383173 493529 383207
rect 493563 383173 493597 383207
rect 493631 383173 493665 383207
rect 493699 383173 493733 383207
rect 493767 383173 493801 383207
rect 493835 383173 493869 383207
rect 493903 383173 493937 383207
rect 493971 383173 494005 383207
rect 494039 383173 494073 383207
rect 494107 383173 494141 383207
rect 494175 383173 494209 383207
rect 494243 383173 494277 383207
rect 494311 383173 494345 383207
rect 494379 383173 494413 383207
rect 494447 383173 494481 383207
rect 494515 383173 494549 383207
rect 494583 383173 494617 383207
rect 497119 383355 497153 383389
rect 497187 383355 497221 383389
rect 497255 383355 497289 383389
rect 497323 383355 497357 383389
rect 497391 383355 497425 383389
rect 497459 383355 497493 383389
rect 497527 383355 497561 383389
rect 497595 383355 497629 383389
rect 497663 383355 497697 383389
rect 497731 383355 497765 383389
rect 497799 383355 497833 383389
rect 497867 383355 497901 383389
rect 497935 383355 497969 383389
rect 498003 383355 498037 383389
rect 498071 383355 498105 383389
rect 498139 383355 498173 383389
rect 498207 383355 498241 383389
rect 498275 383355 498309 383389
rect 498343 383355 498377 383389
rect 500879 383245 500913 383279
rect 500947 383245 500981 383279
rect 501015 383245 501049 383279
rect 501083 383245 501117 383279
rect 501151 383245 501185 383279
rect 501219 383245 501253 383279
rect 501287 383245 501321 383279
rect 501355 383245 501389 383279
rect 501423 383245 501457 383279
rect 501491 383245 501525 383279
rect 501559 383245 501593 383279
rect 501627 383245 501661 383279
rect 501695 383245 501729 383279
rect 501763 383245 501797 383279
rect 501831 383245 501865 383279
rect 501899 383245 501933 383279
rect 501967 383245 502001 383279
rect 502035 383245 502069 383279
rect 502103 383245 502137 383279
rect 493359 382715 493393 382749
rect 493427 382715 493461 382749
rect 493495 382715 493529 382749
rect 493563 382715 493597 382749
rect 493631 382715 493665 382749
rect 493699 382715 493733 382749
rect 493767 382715 493801 382749
rect 493835 382715 493869 382749
rect 493903 382715 493937 382749
rect 493971 382715 494005 382749
rect 494039 382715 494073 382749
rect 494107 382715 494141 382749
rect 494175 382715 494209 382749
rect 494243 382715 494277 382749
rect 494311 382715 494345 382749
rect 494379 382715 494413 382749
rect 494447 382715 494481 382749
rect 494515 382715 494549 382749
rect 494583 382715 494617 382749
rect 497119 382897 497153 382931
rect 497187 382897 497221 382931
rect 497255 382897 497289 382931
rect 497323 382897 497357 382931
rect 497391 382897 497425 382931
rect 497459 382897 497493 382931
rect 497527 382897 497561 382931
rect 497595 382897 497629 382931
rect 497663 382897 497697 382931
rect 497731 382897 497765 382931
rect 497799 382897 497833 382931
rect 497867 382897 497901 382931
rect 497935 382897 497969 382931
rect 498003 382897 498037 382931
rect 498071 382897 498105 382931
rect 498139 382897 498173 382931
rect 498207 382897 498241 382931
rect 498275 382897 498309 382931
rect 498343 382897 498377 382931
rect 500879 382787 500913 382821
rect 500947 382787 500981 382821
rect 501015 382787 501049 382821
rect 501083 382787 501117 382821
rect 501151 382787 501185 382821
rect 501219 382787 501253 382821
rect 501287 382787 501321 382821
rect 501355 382787 501389 382821
rect 501423 382787 501457 382821
rect 501491 382787 501525 382821
rect 501559 382787 501593 382821
rect 501627 382787 501661 382821
rect 501695 382787 501729 382821
rect 501763 382787 501797 382821
rect 501831 382787 501865 382821
rect 501899 382787 501933 382821
rect 501967 382787 502001 382821
rect 502035 382787 502069 382821
rect 502103 382787 502137 382821
rect 497119 382439 497153 382473
rect 497187 382439 497221 382473
rect 497255 382439 497289 382473
rect 497323 382439 497357 382473
rect 497391 382439 497425 382473
rect 497459 382439 497493 382473
rect 497527 382439 497561 382473
rect 497595 382439 497629 382473
rect 497663 382439 497697 382473
rect 497731 382439 497765 382473
rect 497799 382439 497833 382473
rect 497867 382439 497901 382473
rect 497935 382439 497969 382473
rect 498003 382439 498037 382473
rect 498071 382439 498105 382473
rect 498139 382439 498173 382473
rect 498207 382439 498241 382473
rect 498275 382439 498309 382473
rect 498343 382439 498377 382473
rect 493359 382257 493393 382291
rect 493427 382257 493461 382291
rect 493495 382257 493529 382291
rect 493563 382257 493597 382291
rect 493631 382257 493665 382291
rect 493699 382257 493733 382291
rect 493767 382257 493801 382291
rect 493835 382257 493869 382291
rect 493903 382257 493937 382291
rect 493971 382257 494005 382291
rect 494039 382257 494073 382291
rect 494107 382257 494141 382291
rect 494175 382257 494209 382291
rect 494243 382257 494277 382291
rect 494311 382257 494345 382291
rect 494379 382257 494413 382291
rect 494447 382257 494481 382291
rect 494515 382257 494549 382291
rect 494583 382257 494617 382291
rect 523439 385005 523473 385039
rect 523507 385005 523541 385039
rect 523575 385005 523609 385039
rect 523643 385005 523677 385039
rect 523711 385005 523745 385039
rect 523779 385005 523813 385039
rect 523847 385005 523881 385039
rect 523915 385005 523949 385039
rect 523983 385005 524017 385039
rect 524051 385005 524085 385039
rect 524119 385005 524153 385039
rect 524187 385005 524221 385039
rect 524255 385005 524289 385039
rect 524323 385005 524357 385039
rect 524391 385005 524425 385039
rect 524459 385005 524493 385039
rect 524527 385005 524561 385039
rect 524595 385005 524629 385039
rect 524663 385005 524697 385039
rect 523439 384547 523473 384581
rect 523507 384547 523541 384581
rect 523575 384547 523609 384581
rect 523643 384547 523677 384581
rect 523711 384547 523745 384581
rect 523779 384547 523813 384581
rect 523847 384547 523881 384581
rect 523915 384547 523949 384581
rect 523983 384547 524017 384581
rect 524051 384547 524085 384581
rect 524119 384547 524153 384581
rect 524187 384547 524221 384581
rect 524255 384547 524289 384581
rect 524323 384547 524357 384581
rect 524391 384547 524425 384581
rect 524459 384547 524493 384581
rect 524527 384547 524561 384581
rect 524595 384547 524629 384581
rect 524663 384547 524697 384581
rect 523439 384089 523473 384123
rect 523507 384089 523541 384123
rect 523575 384089 523609 384123
rect 523643 384089 523677 384123
rect 523711 384089 523745 384123
rect 523779 384089 523813 384123
rect 523847 384089 523881 384123
rect 523915 384089 523949 384123
rect 523983 384089 524017 384123
rect 524051 384089 524085 384123
rect 524119 384089 524153 384123
rect 524187 384089 524221 384123
rect 524255 384089 524289 384123
rect 524323 384089 524357 384123
rect 524391 384089 524425 384123
rect 524459 384089 524493 384123
rect 524527 384089 524561 384123
rect 524595 384089 524629 384123
rect 524663 384089 524697 384123
rect 523439 383631 523473 383665
rect 523507 383631 523541 383665
rect 523575 383631 523609 383665
rect 523643 383631 523677 383665
rect 523711 383631 523745 383665
rect 523779 383631 523813 383665
rect 523847 383631 523881 383665
rect 523915 383631 523949 383665
rect 523983 383631 524017 383665
rect 524051 383631 524085 383665
rect 524119 383631 524153 383665
rect 524187 383631 524221 383665
rect 524255 383631 524289 383665
rect 524323 383631 524357 383665
rect 524391 383631 524425 383665
rect 524459 383631 524493 383665
rect 524527 383631 524561 383665
rect 524595 383631 524629 383665
rect 524663 383631 524697 383665
rect 523439 383173 523473 383207
rect 523507 383173 523541 383207
rect 523575 383173 523609 383207
rect 523643 383173 523677 383207
rect 523711 383173 523745 383207
rect 523779 383173 523813 383207
rect 523847 383173 523881 383207
rect 523915 383173 523949 383207
rect 523983 383173 524017 383207
rect 524051 383173 524085 383207
rect 524119 383173 524153 383207
rect 524187 383173 524221 383207
rect 524255 383173 524289 383207
rect 524323 383173 524357 383207
rect 524391 383173 524425 383207
rect 524459 383173 524493 383207
rect 524527 383173 524561 383207
rect 524595 383173 524629 383207
rect 524663 383173 524697 383207
rect 523439 382715 523473 382749
rect 523507 382715 523541 382749
rect 523575 382715 523609 382749
rect 523643 382715 523677 382749
rect 523711 382715 523745 382749
rect 523779 382715 523813 382749
rect 523847 382715 523881 382749
rect 523915 382715 523949 382749
rect 523983 382715 524017 382749
rect 524051 382715 524085 382749
rect 524119 382715 524153 382749
rect 524187 382715 524221 382749
rect 524255 382715 524289 382749
rect 524323 382715 524357 382749
rect 524391 382715 524425 382749
rect 524459 382715 524493 382749
rect 524527 382715 524561 382749
rect 524595 382715 524629 382749
rect 524663 382715 524697 382749
rect 500879 382329 500913 382363
rect 500947 382329 500981 382363
rect 501015 382329 501049 382363
rect 501083 382329 501117 382363
rect 501151 382329 501185 382363
rect 501219 382329 501253 382363
rect 501287 382329 501321 382363
rect 501355 382329 501389 382363
rect 501423 382329 501457 382363
rect 501491 382329 501525 382363
rect 501559 382329 501593 382363
rect 501627 382329 501661 382363
rect 501695 382329 501729 382363
rect 501763 382329 501797 382363
rect 501831 382329 501865 382363
rect 501899 382329 501933 382363
rect 501967 382329 502001 382363
rect 502035 382329 502069 382363
rect 502103 382329 502137 382363
rect 493359 381799 493393 381833
rect 493427 381799 493461 381833
rect 493495 381799 493529 381833
rect 493563 381799 493597 381833
rect 493631 381799 493665 381833
rect 493699 381799 493733 381833
rect 493767 381799 493801 381833
rect 493835 381799 493869 381833
rect 493903 381799 493937 381833
rect 493971 381799 494005 381833
rect 494039 381799 494073 381833
rect 494107 381799 494141 381833
rect 494175 381799 494209 381833
rect 494243 381799 494277 381833
rect 494311 381799 494345 381833
rect 494379 381799 494413 381833
rect 494447 381799 494481 381833
rect 494515 381799 494549 381833
rect 494583 381799 494617 381833
rect 497119 381981 497153 382015
rect 497187 381981 497221 382015
rect 497255 381981 497289 382015
rect 497323 381981 497357 382015
rect 497391 381981 497425 382015
rect 497459 381981 497493 382015
rect 497527 381981 497561 382015
rect 497595 381981 497629 382015
rect 497663 381981 497697 382015
rect 497731 381981 497765 382015
rect 497799 381981 497833 382015
rect 497867 381981 497901 382015
rect 497935 381981 497969 382015
rect 498003 381981 498037 382015
rect 498071 381981 498105 382015
rect 498139 381981 498173 382015
rect 498207 381981 498241 382015
rect 498275 381981 498309 382015
rect 498343 381981 498377 382015
rect 523439 382257 523473 382291
rect 523507 382257 523541 382291
rect 523575 382257 523609 382291
rect 523643 382257 523677 382291
rect 523711 382257 523745 382291
rect 523779 382257 523813 382291
rect 523847 382257 523881 382291
rect 523915 382257 523949 382291
rect 523983 382257 524017 382291
rect 524051 382257 524085 382291
rect 524119 382257 524153 382291
rect 524187 382257 524221 382291
rect 524255 382257 524289 382291
rect 524323 382257 524357 382291
rect 524391 382257 524425 382291
rect 524459 382257 524493 382291
rect 524527 382257 524561 382291
rect 524595 382257 524629 382291
rect 524663 382257 524697 382291
rect 500879 381871 500913 381905
rect 500947 381871 500981 381905
rect 501015 381871 501049 381905
rect 501083 381871 501117 381905
rect 501151 381871 501185 381905
rect 501219 381871 501253 381905
rect 501287 381871 501321 381905
rect 501355 381871 501389 381905
rect 501423 381871 501457 381905
rect 501491 381871 501525 381905
rect 501559 381871 501593 381905
rect 501627 381871 501661 381905
rect 501695 381871 501729 381905
rect 501763 381871 501797 381905
rect 501831 381871 501865 381905
rect 501899 381871 501933 381905
rect 501967 381871 502001 381905
rect 502035 381871 502069 381905
rect 502103 381871 502137 381905
rect 497119 381523 497153 381557
rect 497187 381523 497221 381557
rect 497255 381523 497289 381557
rect 497323 381523 497357 381557
rect 497391 381523 497425 381557
rect 497459 381523 497493 381557
rect 497527 381523 497561 381557
rect 497595 381523 497629 381557
rect 497663 381523 497697 381557
rect 497731 381523 497765 381557
rect 497799 381523 497833 381557
rect 497867 381523 497901 381557
rect 497935 381523 497969 381557
rect 498003 381523 498037 381557
rect 498071 381523 498105 381557
rect 498139 381523 498173 381557
rect 498207 381523 498241 381557
rect 498275 381523 498309 381557
rect 498343 381523 498377 381557
rect 493359 381341 493393 381375
rect 493427 381341 493461 381375
rect 493495 381341 493529 381375
rect 493563 381341 493597 381375
rect 493631 381341 493665 381375
rect 493699 381341 493733 381375
rect 493767 381341 493801 381375
rect 493835 381341 493869 381375
rect 493903 381341 493937 381375
rect 493971 381341 494005 381375
rect 494039 381341 494073 381375
rect 494107 381341 494141 381375
rect 494175 381341 494209 381375
rect 494243 381341 494277 381375
rect 494311 381341 494345 381375
rect 494379 381341 494413 381375
rect 494447 381341 494481 381375
rect 494515 381341 494549 381375
rect 494583 381341 494617 381375
rect 523439 381799 523473 381833
rect 523507 381799 523541 381833
rect 523575 381799 523609 381833
rect 523643 381799 523677 381833
rect 523711 381799 523745 381833
rect 523779 381799 523813 381833
rect 523847 381799 523881 381833
rect 523915 381799 523949 381833
rect 523983 381799 524017 381833
rect 524051 381799 524085 381833
rect 524119 381799 524153 381833
rect 524187 381799 524221 381833
rect 524255 381799 524289 381833
rect 524323 381799 524357 381833
rect 524391 381799 524425 381833
rect 524459 381799 524493 381833
rect 524527 381799 524561 381833
rect 524595 381799 524629 381833
rect 524663 381799 524697 381833
rect 500879 381413 500913 381447
rect 500947 381413 500981 381447
rect 501015 381413 501049 381447
rect 501083 381413 501117 381447
rect 501151 381413 501185 381447
rect 501219 381413 501253 381447
rect 501287 381413 501321 381447
rect 501355 381413 501389 381447
rect 501423 381413 501457 381447
rect 501491 381413 501525 381447
rect 501559 381413 501593 381447
rect 501627 381413 501661 381447
rect 501695 381413 501729 381447
rect 501763 381413 501797 381447
rect 501831 381413 501865 381447
rect 501899 381413 501933 381447
rect 501967 381413 502001 381447
rect 502035 381413 502069 381447
rect 502103 381413 502137 381447
rect 493359 380883 493393 380917
rect 493427 380883 493461 380917
rect 493495 380883 493529 380917
rect 493563 380883 493597 380917
rect 493631 380883 493665 380917
rect 493699 380883 493733 380917
rect 493767 380883 493801 380917
rect 493835 380883 493869 380917
rect 493903 380883 493937 380917
rect 493971 380883 494005 380917
rect 494039 380883 494073 380917
rect 494107 380883 494141 380917
rect 494175 380883 494209 380917
rect 494243 380883 494277 380917
rect 494311 380883 494345 380917
rect 494379 380883 494413 380917
rect 494447 380883 494481 380917
rect 494515 380883 494549 380917
rect 494583 380883 494617 380917
rect 497119 381065 497153 381099
rect 497187 381065 497221 381099
rect 497255 381065 497289 381099
rect 497323 381065 497357 381099
rect 497391 381065 497425 381099
rect 497459 381065 497493 381099
rect 497527 381065 497561 381099
rect 497595 381065 497629 381099
rect 497663 381065 497697 381099
rect 497731 381065 497765 381099
rect 497799 381065 497833 381099
rect 497867 381065 497901 381099
rect 497935 381065 497969 381099
rect 498003 381065 498037 381099
rect 498071 381065 498105 381099
rect 498139 381065 498173 381099
rect 498207 381065 498241 381099
rect 498275 381065 498309 381099
rect 498343 381065 498377 381099
rect 493359 380425 493393 380459
rect 493427 380425 493461 380459
rect 493495 380425 493529 380459
rect 493563 380425 493597 380459
rect 493631 380425 493665 380459
rect 493699 380425 493733 380459
rect 493767 380425 493801 380459
rect 493835 380425 493869 380459
rect 493903 380425 493937 380459
rect 493971 380425 494005 380459
rect 494039 380425 494073 380459
rect 494107 380425 494141 380459
rect 494175 380425 494209 380459
rect 494243 380425 494277 380459
rect 494311 380425 494345 380459
rect 494379 380425 494413 380459
rect 494447 380425 494481 380459
rect 494515 380425 494549 380459
rect 494583 380425 494617 380459
rect 500879 380955 500913 380989
rect 500947 380955 500981 380989
rect 501015 380955 501049 380989
rect 501083 380955 501117 380989
rect 501151 380955 501185 380989
rect 501219 380955 501253 380989
rect 501287 380955 501321 380989
rect 501355 380955 501389 380989
rect 501423 380955 501457 380989
rect 501491 380955 501525 380989
rect 501559 380955 501593 380989
rect 501627 380955 501661 380989
rect 501695 380955 501729 380989
rect 501763 380955 501797 380989
rect 501831 380955 501865 380989
rect 501899 380955 501933 380989
rect 501967 380955 502001 380989
rect 502035 380955 502069 380989
rect 502103 380955 502137 380989
rect 497119 380607 497153 380641
rect 497187 380607 497221 380641
rect 497255 380607 497289 380641
rect 497323 380607 497357 380641
rect 497391 380607 497425 380641
rect 497459 380607 497493 380641
rect 497527 380607 497561 380641
rect 497595 380607 497629 380641
rect 497663 380607 497697 380641
rect 497731 380607 497765 380641
rect 497799 380607 497833 380641
rect 497867 380607 497901 380641
rect 497935 380607 497969 380641
rect 498003 380607 498037 380641
rect 498071 380607 498105 380641
rect 498139 380607 498173 380641
rect 498207 380607 498241 380641
rect 498275 380607 498309 380641
rect 498343 380607 498377 380641
rect 500879 380497 500913 380531
rect 500947 380497 500981 380531
rect 501015 380497 501049 380531
rect 501083 380497 501117 380531
rect 501151 380497 501185 380531
rect 501219 380497 501253 380531
rect 501287 380497 501321 380531
rect 501355 380497 501389 380531
rect 501423 380497 501457 380531
rect 501491 380497 501525 380531
rect 501559 380497 501593 380531
rect 501627 380497 501661 380531
rect 501695 380497 501729 380531
rect 501763 380497 501797 380531
rect 501831 380497 501865 380531
rect 501899 380497 501933 380531
rect 501967 380497 502001 380531
rect 502035 380497 502069 380531
rect 502103 380497 502137 380531
rect 493359 379967 493393 380001
rect 493427 379967 493461 380001
rect 493495 379967 493529 380001
rect 493563 379967 493597 380001
rect 493631 379967 493665 380001
rect 493699 379967 493733 380001
rect 493767 379967 493801 380001
rect 493835 379967 493869 380001
rect 493903 379967 493937 380001
rect 493971 379967 494005 380001
rect 494039 379967 494073 380001
rect 494107 379967 494141 380001
rect 494175 379967 494209 380001
rect 494243 379967 494277 380001
rect 494311 379967 494345 380001
rect 494379 379967 494413 380001
rect 494447 379967 494481 380001
rect 494515 379967 494549 380001
rect 494583 379967 494617 380001
rect 497119 380149 497153 380183
rect 497187 380149 497221 380183
rect 497255 380149 497289 380183
rect 497323 380149 497357 380183
rect 497391 380149 497425 380183
rect 497459 380149 497493 380183
rect 497527 380149 497561 380183
rect 497595 380149 497629 380183
rect 497663 380149 497697 380183
rect 497731 380149 497765 380183
rect 497799 380149 497833 380183
rect 497867 380149 497901 380183
rect 497935 380149 497969 380183
rect 498003 380149 498037 380183
rect 498071 380149 498105 380183
rect 498139 380149 498173 380183
rect 498207 380149 498241 380183
rect 498275 380149 498309 380183
rect 498343 380149 498377 380183
rect 500879 380039 500913 380073
rect 500947 380039 500981 380073
rect 501015 380039 501049 380073
rect 501083 380039 501117 380073
rect 501151 380039 501185 380073
rect 501219 380039 501253 380073
rect 501287 380039 501321 380073
rect 501355 380039 501389 380073
rect 501423 380039 501457 380073
rect 501491 380039 501525 380073
rect 501559 380039 501593 380073
rect 501627 380039 501661 380073
rect 501695 380039 501729 380073
rect 501763 380039 501797 380073
rect 501831 380039 501865 380073
rect 501899 380039 501933 380073
rect 501967 380039 502001 380073
rect 502035 380039 502069 380073
rect 502103 380039 502137 380073
rect 493359 379509 493393 379543
rect 493427 379509 493461 379543
rect 493495 379509 493529 379543
rect 493563 379509 493597 379543
rect 493631 379509 493665 379543
rect 493699 379509 493733 379543
rect 493767 379509 493801 379543
rect 493835 379509 493869 379543
rect 493903 379509 493937 379543
rect 493971 379509 494005 379543
rect 494039 379509 494073 379543
rect 494107 379509 494141 379543
rect 494175 379509 494209 379543
rect 494243 379509 494277 379543
rect 494311 379509 494345 379543
rect 494379 379509 494413 379543
rect 494447 379509 494481 379543
rect 494515 379509 494549 379543
rect 494583 379509 494617 379543
rect 497119 379691 497153 379725
rect 497187 379691 497221 379725
rect 497255 379691 497289 379725
rect 497323 379691 497357 379725
rect 497391 379691 497425 379725
rect 497459 379691 497493 379725
rect 497527 379691 497561 379725
rect 497595 379691 497629 379725
rect 497663 379691 497697 379725
rect 497731 379691 497765 379725
rect 497799 379691 497833 379725
rect 497867 379691 497901 379725
rect 497935 379691 497969 379725
rect 498003 379691 498037 379725
rect 498071 379691 498105 379725
rect 498139 379691 498173 379725
rect 498207 379691 498241 379725
rect 498275 379691 498309 379725
rect 498343 379691 498377 379725
rect 523439 381341 523473 381375
rect 523507 381341 523541 381375
rect 523575 381341 523609 381375
rect 523643 381341 523677 381375
rect 523711 381341 523745 381375
rect 523779 381341 523813 381375
rect 523847 381341 523881 381375
rect 523915 381341 523949 381375
rect 523983 381341 524017 381375
rect 524051 381341 524085 381375
rect 524119 381341 524153 381375
rect 524187 381341 524221 381375
rect 524255 381341 524289 381375
rect 524323 381341 524357 381375
rect 524391 381341 524425 381375
rect 524459 381341 524493 381375
rect 524527 381341 524561 381375
rect 524595 381341 524629 381375
rect 524663 381341 524697 381375
rect 523439 380883 523473 380917
rect 523507 380883 523541 380917
rect 523575 380883 523609 380917
rect 523643 380883 523677 380917
rect 523711 380883 523745 380917
rect 523779 380883 523813 380917
rect 523847 380883 523881 380917
rect 523915 380883 523949 380917
rect 523983 380883 524017 380917
rect 524051 380883 524085 380917
rect 524119 380883 524153 380917
rect 524187 380883 524221 380917
rect 524255 380883 524289 380917
rect 524323 380883 524357 380917
rect 524391 380883 524425 380917
rect 524459 380883 524493 380917
rect 524527 380883 524561 380917
rect 524595 380883 524629 380917
rect 524663 380883 524697 380917
rect 523439 380425 523473 380459
rect 523507 380425 523541 380459
rect 523575 380425 523609 380459
rect 523643 380425 523677 380459
rect 523711 380425 523745 380459
rect 523779 380425 523813 380459
rect 523847 380425 523881 380459
rect 523915 380425 523949 380459
rect 523983 380425 524017 380459
rect 524051 380425 524085 380459
rect 524119 380425 524153 380459
rect 524187 380425 524221 380459
rect 524255 380425 524289 380459
rect 524323 380425 524357 380459
rect 524391 380425 524425 380459
rect 524459 380425 524493 380459
rect 524527 380425 524561 380459
rect 524595 380425 524629 380459
rect 524663 380425 524697 380459
rect 523439 379967 523473 380001
rect 523507 379967 523541 380001
rect 523575 379967 523609 380001
rect 523643 379967 523677 380001
rect 523711 379967 523745 380001
rect 523779 379967 523813 380001
rect 523847 379967 523881 380001
rect 523915 379967 523949 380001
rect 523983 379967 524017 380001
rect 524051 379967 524085 380001
rect 524119 379967 524153 380001
rect 524187 379967 524221 380001
rect 524255 379967 524289 380001
rect 524323 379967 524357 380001
rect 524391 379967 524425 380001
rect 524459 379967 524493 380001
rect 524527 379967 524561 380001
rect 524595 379967 524629 380001
rect 524663 379967 524697 380001
rect 523439 379509 523473 379543
rect 523507 379509 523541 379543
rect 523575 379509 523609 379543
rect 523643 379509 523677 379543
rect 523711 379509 523745 379543
rect 523779 379509 523813 379543
rect 523847 379509 523881 379543
rect 523915 379509 523949 379543
rect 523983 379509 524017 379543
rect 524051 379509 524085 379543
rect 524119 379509 524153 379543
rect 524187 379509 524221 379543
rect 524255 379509 524289 379543
rect 524323 379509 524357 379543
rect 524391 379509 524425 379543
rect 524459 379509 524493 379543
rect 524527 379509 524561 379543
rect 524595 379509 524629 379543
rect 524663 379509 524697 379543
rect 497119 379233 497153 379267
rect 497187 379233 497221 379267
rect 497255 379233 497289 379267
rect 497323 379233 497357 379267
rect 497391 379233 497425 379267
rect 497459 379233 497493 379267
rect 497527 379233 497561 379267
rect 497595 379233 497629 379267
rect 497663 379233 497697 379267
rect 497731 379233 497765 379267
rect 497799 379233 497833 379267
rect 497867 379233 497901 379267
rect 497935 379233 497969 379267
rect 498003 379233 498037 379267
rect 498071 379233 498105 379267
rect 498139 379233 498173 379267
rect 498207 379233 498241 379267
rect 498275 379233 498309 379267
rect 498343 379233 498377 379267
rect 493359 379051 493393 379085
rect 493427 379051 493461 379085
rect 493495 379051 493529 379085
rect 493563 379051 493597 379085
rect 493631 379051 493665 379085
rect 493699 379051 493733 379085
rect 493767 379051 493801 379085
rect 493835 379051 493869 379085
rect 493903 379051 493937 379085
rect 493971 379051 494005 379085
rect 494039 379051 494073 379085
rect 494107 379051 494141 379085
rect 494175 379051 494209 379085
rect 494243 379051 494277 379085
rect 494311 379051 494345 379085
rect 494379 379051 494413 379085
rect 494447 379051 494481 379085
rect 494515 379051 494549 379085
rect 494583 379051 494617 379085
rect 523439 379051 523473 379085
rect 523507 379051 523541 379085
rect 523575 379051 523609 379085
rect 523643 379051 523677 379085
rect 523711 379051 523745 379085
rect 523779 379051 523813 379085
rect 523847 379051 523881 379085
rect 523915 379051 523949 379085
rect 523983 379051 524017 379085
rect 524051 379051 524085 379085
rect 524119 379051 524153 379085
rect 524187 379051 524221 379085
rect 524255 379051 524289 379085
rect 524323 379051 524357 379085
rect 524391 379051 524425 379085
rect 524459 379051 524493 379085
rect 524527 379051 524561 379085
rect 524595 379051 524629 379085
rect 524663 379051 524697 379085
rect 497119 378775 497153 378809
rect 497187 378775 497221 378809
rect 497255 378775 497289 378809
rect 497323 378775 497357 378809
rect 497391 378775 497425 378809
rect 497459 378775 497493 378809
rect 497527 378775 497561 378809
rect 497595 378775 497629 378809
rect 497663 378775 497697 378809
rect 497731 378775 497765 378809
rect 497799 378775 497833 378809
rect 497867 378775 497901 378809
rect 497935 378775 497969 378809
rect 498003 378775 498037 378809
rect 498071 378775 498105 378809
rect 498139 378775 498173 378809
rect 498207 378775 498241 378809
rect 498275 378775 498309 378809
rect 498343 378775 498377 378809
rect 493359 378593 493393 378627
rect 493427 378593 493461 378627
rect 493495 378593 493529 378627
rect 493563 378593 493597 378627
rect 493631 378593 493665 378627
rect 493699 378593 493733 378627
rect 493767 378593 493801 378627
rect 493835 378593 493869 378627
rect 493903 378593 493937 378627
rect 493971 378593 494005 378627
rect 494039 378593 494073 378627
rect 494107 378593 494141 378627
rect 494175 378593 494209 378627
rect 494243 378593 494277 378627
rect 494311 378593 494345 378627
rect 494379 378593 494413 378627
rect 494447 378593 494481 378627
rect 494515 378593 494549 378627
rect 494583 378593 494617 378627
rect 523439 378593 523473 378627
rect 523507 378593 523541 378627
rect 523575 378593 523609 378627
rect 523643 378593 523677 378627
rect 523711 378593 523745 378627
rect 523779 378593 523813 378627
rect 523847 378593 523881 378627
rect 523915 378593 523949 378627
rect 523983 378593 524017 378627
rect 524051 378593 524085 378627
rect 524119 378593 524153 378627
rect 524187 378593 524221 378627
rect 524255 378593 524289 378627
rect 524323 378593 524357 378627
rect 524391 378593 524425 378627
rect 524459 378593 524493 378627
rect 524527 378593 524561 378627
rect 524595 378593 524629 378627
rect 524663 378593 524697 378627
rect 493359 378135 493393 378169
rect 493427 378135 493461 378169
rect 493495 378135 493529 378169
rect 493563 378135 493597 378169
rect 493631 378135 493665 378169
rect 493699 378135 493733 378169
rect 493767 378135 493801 378169
rect 493835 378135 493869 378169
rect 493903 378135 493937 378169
rect 493971 378135 494005 378169
rect 494039 378135 494073 378169
rect 494107 378135 494141 378169
rect 494175 378135 494209 378169
rect 494243 378135 494277 378169
rect 494311 378135 494345 378169
rect 494379 378135 494413 378169
rect 494447 378135 494481 378169
rect 494515 378135 494549 378169
rect 494583 378135 494617 378169
rect 497119 378317 497153 378351
rect 497187 378317 497221 378351
rect 497255 378317 497289 378351
rect 497323 378317 497357 378351
rect 497391 378317 497425 378351
rect 497459 378317 497493 378351
rect 497527 378317 497561 378351
rect 497595 378317 497629 378351
rect 497663 378317 497697 378351
rect 497731 378317 497765 378351
rect 497799 378317 497833 378351
rect 497867 378317 497901 378351
rect 497935 378317 497969 378351
rect 498003 378317 498037 378351
rect 498071 378317 498105 378351
rect 498139 378317 498173 378351
rect 498207 378317 498241 378351
rect 498275 378317 498309 378351
rect 498343 378317 498377 378351
rect 493359 377677 493393 377711
rect 493427 377677 493461 377711
rect 493495 377677 493529 377711
rect 493563 377677 493597 377711
rect 493631 377677 493665 377711
rect 493699 377677 493733 377711
rect 493767 377677 493801 377711
rect 493835 377677 493869 377711
rect 493903 377677 493937 377711
rect 493971 377677 494005 377711
rect 494039 377677 494073 377711
rect 494107 377677 494141 377711
rect 494175 377677 494209 377711
rect 494243 377677 494277 377711
rect 494311 377677 494345 377711
rect 494379 377677 494413 377711
rect 494447 377677 494481 377711
rect 494515 377677 494549 377711
rect 494583 377677 494617 377711
rect 523439 378135 523473 378169
rect 523507 378135 523541 378169
rect 523575 378135 523609 378169
rect 523643 378135 523677 378169
rect 523711 378135 523745 378169
rect 523779 378135 523813 378169
rect 523847 378135 523881 378169
rect 523915 378135 523949 378169
rect 523983 378135 524017 378169
rect 524051 378135 524085 378169
rect 524119 378135 524153 378169
rect 524187 378135 524221 378169
rect 524255 378135 524289 378169
rect 524323 378135 524357 378169
rect 524391 378135 524425 378169
rect 524459 378135 524493 378169
rect 524527 378135 524561 378169
rect 524595 378135 524629 378169
rect 524663 378135 524697 378169
rect 497119 377859 497153 377893
rect 497187 377859 497221 377893
rect 497255 377859 497289 377893
rect 497323 377859 497357 377893
rect 497391 377859 497425 377893
rect 497459 377859 497493 377893
rect 497527 377859 497561 377893
rect 497595 377859 497629 377893
rect 497663 377859 497697 377893
rect 497731 377859 497765 377893
rect 497799 377859 497833 377893
rect 497867 377859 497901 377893
rect 497935 377859 497969 377893
rect 498003 377859 498037 377893
rect 498071 377859 498105 377893
rect 498139 377859 498173 377893
rect 498207 377859 498241 377893
rect 498275 377859 498309 377893
rect 498343 377859 498377 377893
rect 493359 377219 493393 377253
rect 493427 377219 493461 377253
rect 493495 377219 493529 377253
rect 493563 377219 493597 377253
rect 493631 377219 493665 377253
rect 493699 377219 493733 377253
rect 493767 377219 493801 377253
rect 493835 377219 493869 377253
rect 493903 377219 493937 377253
rect 493971 377219 494005 377253
rect 494039 377219 494073 377253
rect 494107 377219 494141 377253
rect 494175 377219 494209 377253
rect 494243 377219 494277 377253
rect 494311 377219 494345 377253
rect 494379 377219 494413 377253
rect 494447 377219 494481 377253
rect 494515 377219 494549 377253
rect 494583 377219 494617 377253
rect 497119 377401 497153 377435
rect 497187 377401 497221 377435
rect 497255 377401 497289 377435
rect 497323 377401 497357 377435
rect 497391 377401 497425 377435
rect 497459 377401 497493 377435
rect 497527 377401 497561 377435
rect 497595 377401 497629 377435
rect 497663 377401 497697 377435
rect 497731 377401 497765 377435
rect 497799 377401 497833 377435
rect 497867 377401 497901 377435
rect 497935 377401 497969 377435
rect 498003 377401 498037 377435
rect 498071 377401 498105 377435
rect 498139 377401 498173 377435
rect 498207 377401 498241 377435
rect 498275 377401 498309 377435
rect 498343 377401 498377 377435
rect 493359 376761 493393 376795
rect 493427 376761 493461 376795
rect 493495 376761 493529 376795
rect 493563 376761 493597 376795
rect 493631 376761 493665 376795
rect 493699 376761 493733 376795
rect 493767 376761 493801 376795
rect 493835 376761 493869 376795
rect 493903 376761 493937 376795
rect 493971 376761 494005 376795
rect 494039 376761 494073 376795
rect 494107 376761 494141 376795
rect 494175 376761 494209 376795
rect 494243 376761 494277 376795
rect 494311 376761 494345 376795
rect 494379 376761 494413 376795
rect 494447 376761 494481 376795
rect 494515 376761 494549 376795
rect 494583 376761 494617 376795
rect 523439 377677 523473 377711
rect 523507 377677 523541 377711
rect 523575 377677 523609 377711
rect 523643 377677 523677 377711
rect 523711 377677 523745 377711
rect 523779 377677 523813 377711
rect 523847 377677 523881 377711
rect 523915 377677 523949 377711
rect 523983 377677 524017 377711
rect 524051 377677 524085 377711
rect 524119 377677 524153 377711
rect 524187 377677 524221 377711
rect 524255 377677 524289 377711
rect 524323 377677 524357 377711
rect 524391 377677 524425 377711
rect 524459 377677 524493 377711
rect 524527 377677 524561 377711
rect 524595 377677 524629 377711
rect 524663 377677 524697 377711
rect 504639 377401 504673 377435
rect 504707 377401 504741 377435
rect 504775 377401 504809 377435
rect 504843 377401 504877 377435
rect 504911 377401 504945 377435
rect 504979 377401 505013 377435
rect 505047 377401 505081 377435
rect 505115 377401 505149 377435
rect 505183 377401 505217 377435
rect 505251 377401 505285 377435
rect 505319 377401 505353 377435
rect 505387 377401 505421 377435
rect 505455 377401 505489 377435
rect 505523 377401 505557 377435
rect 505591 377401 505625 377435
rect 505659 377401 505693 377435
rect 505727 377401 505761 377435
rect 505795 377401 505829 377435
rect 505863 377401 505897 377435
rect 497119 376943 497153 376977
rect 497187 376943 497221 376977
rect 497255 376943 497289 376977
rect 497323 376943 497357 376977
rect 497391 376943 497425 376977
rect 497459 376943 497493 376977
rect 497527 376943 497561 376977
rect 497595 376943 497629 376977
rect 497663 376943 497697 376977
rect 497731 376943 497765 376977
rect 497799 376943 497833 376977
rect 497867 376943 497901 376977
rect 497935 376943 497969 376977
rect 498003 376943 498037 376977
rect 498071 376943 498105 376977
rect 498139 376943 498173 376977
rect 498207 376943 498241 376977
rect 498275 376943 498309 376977
rect 498343 376943 498377 376977
rect 493359 376303 493393 376337
rect 493427 376303 493461 376337
rect 493495 376303 493529 376337
rect 493563 376303 493597 376337
rect 493631 376303 493665 376337
rect 493699 376303 493733 376337
rect 493767 376303 493801 376337
rect 493835 376303 493869 376337
rect 493903 376303 493937 376337
rect 493971 376303 494005 376337
rect 494039 376303 494073 376337
rect 494107 376303 494141 376337
rect 494175 376303 494209 376337
rect 494243 376303 494277 376337
rect 494311 376303 494345 376337
rect 494379 376303 494413 376337
rect 494447 376303 494481 376337
rect 494515 376303 494549 376337
rect 494583 376303 494617 376337
rect 512159 377401 512193 377435
rect 512227 377401 512261 377435
rect 512295 377401 512329 377435
rect 512363 377401 512397 377435
rect 512431 377401 512465 377435
rect 512499 377401 512533 377435
rect 512567 377401 512601 377435
rect 512635 377401 512669 377435
rect 512703 377401 512737 377435
rect 512771 377401 512805 377435
rect 512839 377401 512873 377435
rect 512907 377401 512941 377435
rect 512975 377401 513009 377435
rect 513043 377401 513077 377435
rect 513111 377401 513145 377435
rect 513179 377401 513213 377435
rect 513247 377401 513281 377435
rect 513315 377401 513349 377435
rect 513383 377401 513417 377435
rect 504639 376943 504673 376977
rect 504707 376943 504741 376977
rect 504775 376943 504809 376977
rect 504843 376943 504877 376977
rect 504911 376943 504945 376977
rect 504979 376943 505013 376977
rect 505047 376943 505081 376977
rect 505115 376943 505149 376977
rect 505183 376943 505217 376977
rect 505251 376943 505285 376977
rect 505319 376943 505353 376977
rect 505387 376943 505421 376977
rect 505455 376943 505489 376977
rect 505523 376943 505557 376977
rect 505591 376943 505625 376977
rect 505659 376943 505693 376977
rect 505727 376943 505761 376977
rect 505795 376943 505829 376977
rect 505863 376943 505897 376977
rect 497119 376485 497153 376519
rect 497187 376485 497221 376519
rect 497255 376485 497289 376519
rect 497323 376485 497357 376519
rect 497391 376485 497425 376519
rect 497459 376485 497493 376519
rect 497527 376485 497561 376519
rect 497595 376485 497629 376519
rect 497663 376485 497697 376519
rect 497731 376485 497765 376519
rect 497799 376485 497833 376519
rect 497867 376485 497901 376519
rect 497935 376485 497969 376519
rect 498003 376485 498037 376519
rect 498071 376485 498105 376519
rect 498139 376485 498173 376519
rect 498207 376485 498241 376519
rect 498275 376485 498309 376519
rect 498343 376485 498377 376519
rect 512159 376943 512193 376977
rect 512227 376943 512261 376977
rect 512295 376943 512329 376977
rect 512363 376943 512397 376977
rect 512431 376943 512465 376977
rect 512499 376943 512533 376977
rect 512567 376943 512601 376977
rect 512635 376943 512669 376977
rect 512703 376943 512737 376977
rect 512771 376943 512805 376977
rect 512839 376943 512873 376977
rect 512907 376943 512941 376977
rect 512975 376943 513009 376977
rect 513043 376943 513077 376977
rect 513111 376943 513145 376977
rect 513179 376943 513213 376977
rect 513247 376943 513281 376977
rect 513315 376943 513349 376977
rect 513383 376943 513417 376977
rect 504639 376485 504673 376519
rect 504707 376485 504741 376519
rect 504775 376485 504809 376519
rect 504843 376485 504877 376519
rect 504911 376485 504945 376519
rect 504979 376485 505013 376519
rect 505047 376485 505081 376519
rect 505115 376485 505149 376519
rect 505183 376485 505217 376519
rect 505251 376485 505285 376519
rect 505319 376485 505353 376519
rect 505387 376485 505421 376519
rect 505455 376485 505489 376519
rect 505523 376485 505557 376519
rect 505591 376485 505625 376519
rect 505659 376485 505693 376519
rect 505727 376485 505761 376519
rect 505795 376485 505829 376519
rect 505863 376485 505897 376519
rect 497119 376027 497153 376061
rect 497187 376027 497221 376061
rect 497255 376027 497289 376061
rect 497323 376027 497357 376061
rect 497391 376027 497425 376061
rect 497459 376027 497493 376061
rect 497527 376027 497561 376061
rect 497595 376027 497629 376061
rect 497663 376027 497697 376061
rect 497731 376027 497765 376061
rect 497799 376027 497833 376061
rect 497867 376027 497901 376061
rect 497935 376027 497969 376061
rect 498003 376027 498037 376061
rect 498071 376027 498105 376061
rect 498139 376027 498173 376061
rect 498207 376027 498241 376061
rect 498275 376027 498309 376061
rect 498343 376027 498377 376061
rect 493359 375845 493393 375879
rect 493427 375845 493461 375879
rect 493495 375845 493529 375879
rect 493563 375845 493597 375879
rect 493631 375845 493665 375879
rect 493699 375845 493733 375879
rect 493767 375845 493801 375879
rect 493835 375845 493869 375879
rect 493903 375845 493937 375879
rect 493971 375845 494005 375879
rect 494039 375845 494073 375879
rect 494107 375845 494141 375879
rect 494175 375845 494209 375879
rect 494243 375845 494277 375879
rect 494311 375845 494345 375879
rect 494379 375845 494413 375879
rect 494447 375845 494481 375879
rect 494515 375845 494549 375879
rect 494583 375845 494617 375879
rect 512159 376485 512193 376519
rect 512227 376485 512261 376519
rect 512295 376485 512329 376519
rect 512363 376485 512397 376519
rect 512431 376485 512465 376519
rect 512499 376485 512533 376519
rect 512567 376485 512601 376519
rect 512635 376485 512669 376519
rect 512703 376485 512737 376519
rect 512771 376485 512805 376519
rect 512839 376485 512873 376519
rect 512907 376485 512941 376519
rect 512975 376485 513009 376519
rect 513043 376485 513077 376519
rect 513111 376485 513145 376519
rect 513179 376485 513213 376519
rect 513247 376485 513281 376519
rect 513315 376485 513349 376519
rect 513383 376485 513417 376519
rect 504639 376027 504673 376061
rect 504707 376027 504741 376061
rect 504775 376027 504809 376061
rect 504843 376027 504877 376061
rect 504911 376027 504945 376061
rect 504979 376027 505013 376061
rect 505047 376027 505081 376061
rect 505115 376027 505149 376061
rect 505183 376027 505217 376061
rect 505251 376027 505285 376061
rect 505319 376027 505353 376061
rect 505387 376027 505421 376061
rect 505455 376027 505489 376061
rect 505523 376027 505557 376061
rect 505591 376027 505625 376061
rect 505659 376027 505693 376061
rect 505727 376027 505761 376061
rect 505795 376027 505829 376061
rect 505863 376027 505897 376061
rect 497119 375569 497153 375603
rect 497187 375569 497221 375603
rect 497255 375569 497289 375603
rect 497323 375569 497357 375603
rect 497391 375569 497425 375603
rect 497459 375569 497493 375603
rect 497527 375569 497561 375603
rect 497595 375569 497629 375603
rect 497663 375569 497697 375603
rect 497731 375569 497765 375603
rect 497799 375569 497833 375603
rect 497867 375569 497901 375603
rect 497935 375569 497969 375603
rect 498003 375569 498037 375603
rect 498071 375569 498105 375603
rect 498139 375569 498173 375603
rect 498207 375569 498241 375603
rect 498275 375569 498309 375603
rect 498343 375569 498377 375603
rect 493359 375387 493393 375421
rect 493427 375387 493461 375421
rect 493495 375387 493529 375421
rect 493563 375387 493597 375421
rect 493631 375387 493665 375421
rect 493699 375387 493733 375421
rect 493767 375387 493801 375421
rect 493835 375387 493869 375421
rect 493903 375387 493937 375421
rect 493971 375387 494005 375421
rect 494039 375387 494073 375421
rect 494107 375387 494141 375421
rect 494175 375387 494209 375421
rect 494243 375387 494277 375421
rect 494311 375387 494345 375421
rect 494379 375387 494413 375421
rect 494447 375387 494481 375421
rect 494515 375387 494549 375421
rect 494583 375387 494617 375421
rect 512159 376027 512193 376061
rect 512227 376027 512261 376061
rect 512295 376027 512329 376061
rect 512363 376027 512397 376061
rect 512431 376027 512465 376061
rect 512499 376027 512533 376061
rect 512567 376027 512601 376061
rect 512635 376027 512669 376061
rect 512703 376027 512737 376061
rect 512771 376027 512805 376061
rect 512839 376027 512873 376061
rect 512907 376027 512941 376061
rect 512975 376027 513009 376061
rect 513043 376027 513077 376061
rect 513111 376027 513145 376061
rect 513179 376027 513213 376061
rect 513247 376027 513281 376061
rect 513315 376027 513349 376061
rect 513383 376027 513417 376061
rect 504639 375569 504673 375603
rect 504707 375569 504741 375603
rect 504775 375569 504809 375603
rect 504843 375569 504877 375603
rect 504911 375569 504945 375603
rect 504979 375569 505013 375603
rect 505047 375569 505081 375603
rect 505115 375569 505149 375603
rect 505183 375569 505217 375603
rect 505251 375569 505285 375603
rect 505319 375569 505353 375603
rect 505387 375569 505421 375603
rect 505455 375569 505489 375603
rect 505523 375569 505557 375603
rect 505591 375569 505625 375603
rect 505659 375569 505693 375603
rect 505727 375569 505761 375603
rect 505795 375569 505829 375603
rect 505863 375569 505897 375603
rect 493359 374929 493393 374963
rect 493427 374929 493461 374963
rect 493495 374929 493529 374963
rect 493563 374929 493597 374963
rect 493631 374929 493665 374963
rect 493699 374929 493733 374963
rect 493767 374929 493801 374963
rect 493835 374929 493869 374963
rect 493903 374929 493937 374963
rect 493971 374929 494005 374963
rect 494039 374929 494073 374963
rect 494107 374929 494141 374963
rect 494175 374929 494209 374963
rect 494243 374929 494277 374963
rect 494311 374929 494345 374963
rect 494379 374929 494413 374963
rect 494447 374929 494481 374963
rect 494515 374929 494549 374963
rect 494583 374929 494617 374963
rect 497119 375111 497153 375145
rect 497187 375111 497221 375145
rect 497255 375111 497289 375145
rect 497323 375111 497357 375145
rect 497391 375111 497425 375145
rect 497459 375111 497493 375145
rect 497527 375111 497561 375145
rect 497595 375111 497629 375145
rect 497663 375111 497697 375145
rect 497731 375111 497765 375145
rect 497799 375111 497833 375145
rect 497867 375111 497901 375145
rect 497935 375111 497969 375145
rect 498003 375111 498037 375145
rect 498071 375111 498105 375145
rect 498139 375111 498173 375145
rect 498207 375111 498241 375145
rect 498275 375111 498309 375145
rect 498343 375111 498377 375145
rect 493359 374471 493393 374505
rect 493427 374471 493461 374505
rect 493495 374471 493529 374505
rect 493563 374471 493597 374505
rect 493631 374471 493665 374505
rect 493699 374471 493733 374505
rect 493767 374471 493801 374505
rect 493835 374471 493869 374505
rect 493903 374471 493937 374505
rect 493971 374471 494005 374505
rect 494039 374471 494073 374505
rect 494107 374471 494141 374505
rect 494175 374471 494209 374505
rect 494243 374471 494277 374505
rect 494311 374471 494345 374505
rect 494379 374471 494413 374505
rect 494447 374471 494481 374505
rect 494515 374471 494549 374505
rect 494583 374471 494617 374505
rect 512159 375569 512193 375603
rect 512227 375569 512261 375603
rect 512295 375569 512329 375603
rect 512363 375569 512397 375603
rect 512431 375569 512465 375603
rect 512499 375569 512533 375603
rect 512567 375569 512601 375603
rect 512635 375569 512669 375603
rect 512703 375569 512737 375603
rect 512771 375569 512805 375603
rect 512839 375569 512873 375603
rect 512907 375569 512941 375603
rect 512975 375569 513009 375603
rect 513043 375569 513077 375603
rect 513111 375569 513145 375603
rect 513179 375569 513213 375603
rect 513247 375569 513281 375603
rect 513315 375569 513349 375603
rect 513383 375569 513417 375603
rect 504639 375111 504673 375145
rect 504707 375111 504741 375145
rect 504775 375111 504809 375145
rect 504843 375111 504877 375145
rect 504911 375111 504945 375145
rect 504979 375111 505013 375145
rect 505047 375111 505081 375145
rect 505115 375111 505149 375145
rect 505183 375111 505217 375145
rect 505251 375111 505285 375145
rect 505319 375111 505353 375145
rect 505387 375111 505421 375145
rect 505455 375111 505489 375145
rect 505523 375111 505557 375145
rect 505591 375111 505625 375145
rect 505659 375111 505693 375145
rect 505727 375111 505761 375145
rect 505795 375111 505829 375145
rect 505863 375111 505897 375145
rect 497119 374653 497153 374687
rect 497187 374653 497221 374687
rect 497255 374653 497289 374687
rect 497323 374653 497357 374687
rect 497391 374653 497425 374687
rect 497459 374653 497493 374687
rect 497527 374653 497561 374687
rect 497595 374653 497629 374687
rect 497663 374653 497697 374687
rect 497731 374653 497765 374687
rect 497799 374653 497833 374687
rect 497867 374653 497901 374687
rect 497935 374653 497969 374687
rect 498003 374653 498037 374687
rect 498071 374653 498105 374687
rect 498139 374653 498173 374687
rect 498207 374653 498241 374687
rect 498275 374653 498309 374687
rect 498343 374653 498377 374687
rect 493359 374013 493393 374047
rect 493427 374013 493461 374047
rect 493495 374013 493529 374047
rect 493563 374013 493597 374047
rect 493631 374013 493665 374047
rect 493699 374013 493733 374047
rect 493767 374013 493801 374047
rect 493835 374013 493869 374047
rect 493903 374013 493937 374047
rect 493971 374013 494005 374047
rect 494039 374013 494073 374047
rect 494107 374013 494141 374047
rect 494175 374013 494209 374047
rect 494243 374013 494277 374047
rect 494311 374013 494345 374047
rect 494379 374013 494413 374047
rect 494447 374013 494481 374047
rect 494515 374013 494549 374047
rect 494583 374013 494617 374047
rect 497119 374195 497153 374229
rect 497187 374195 497221 374229
rect 497255 374195 497289 374229
rect 497323 374195 497357 374229
rect 497391 374195 497425 374229
rect 497459 374195 497493 374229
rect 497527 374195 497561 374229
rect 497595 374195 497629 374229
rect 497663 374195 497697 374229
rect 497731 374195 497765 374229
rect 497799 374195 497833 374229
rect 497867 374195 497901 374229
rect 497935 374195 497969 374229
rect 498003 374195 498037 374229
rect 498071 374195 498105 374229
rect 498139 374195 498173 374229
rect 498207 374195 498241 374229
rect 498275 374195 498309 374229
rect 498343 374195 498377 374229
rect 493359 373555 493393 373589
rect 493427 373555 493461 373589
rect 493495 373555 493529 373589
rect 493563 373555 493597 373589
rect 493631 373555 493665 373589
rect 493699 373555 493733 373589
rect 493767 373555 493801 373589
rect 493835 373555 493869 373589
rect 493903 373555 493937 373589
rect 493971 373555 494005 373589
rect 494039 373555 494073 373589
rect 494107 373555 494141 373589
rect 494175 373555 494209 373589
rect 494243 373555 494277 373589
rect 494311 373555 494345 373589
rect 494379 373555 494413 373589
rect 494447 373555 494481 373589
rect 494515 373555 494549 373589
rect 494583 373555 494617 373589
rect 512159 375111 512193 375145
rect 512227 375111 512261 375145
rect 512295 375111 512329 375145
rect 512363 375111 512397 375145
rect 512431 375111 512465 375145
rect 512499 375111 512533 375145
rect 512567 375111 512601 375145
rect 512635 375111 512669 375145
rect 512703 375111 512737 375145
rect 512771 375111 512805 375145
rect 512839 375111 512873 375145
rect 512907 375111 512941 375145
rect 512975 375111 513009 375145
rect 513043 375111 513077 375145
rect 513111 375111 513145 375145
rect 513179 375111 513213 375145
rect 513247 375111 513281 375145
rect 513315 375111 513349 375145
rect 513383 375111 513417 375145
rect 504639 374653 504673 374687
rect 504707 374653 504741 374687
rect 504775 374653 504809 374687
rect 504843 374653 504877 374687
rect 504911 374653 504945 374687
rect 504979 374653 505013 374687
rect 505047 374653 505081 374687
rect 505115 374653 505149 374687
rect 505183 374653 505217 374687
rect 505251 374653 505285 374687
rect 505319 374653 505353 374687
rect 505387 374653 505421 374687
rect 505455 374653 505489 374687
rect 505523 374653 505557 374687
rect 505591 374653 505625 374687
rect 505659 374653 505693 374687
rect 505727 374653 505761 374687
rect 505795 374653 505829 374687
rect 505863 374653 505897 374687
rect 497119 373737 497153 373771
rect 497187 373737 497221 373771
rect 497255 373737 497289 373771
rect 497323 373737 497357 373771
rect 497391 373737 497425 373771
rect 497459 373737 497493 373771
rect 497527 373737 497561 373771
rect 497595 373737 497629 373771
rect 497663 373737 497697 373771
rect 497731 373737 497765 373771
rect 497799 373737 497833 373771
rect 497867 373737 497901 373771
rect 497935 373737 497969 373771
rect 498003 373737 498037 373771
rect 498071 373737 498105 373771
rect 498139 373737 498173 373771
rect 498207 373737 498241 373771
rect 498275 373737 498309 373771
rect 498343 373737 498377 373771
rect 523439 377219 523473 377253
rect 523507 377219 523541 377253
rect 523575 377219 523609 377253
rect 523643 377219 523677 377253
rect 523711 377219 523745 377253
rect 523779 377219 523813 377253
rect 523847 377219 523881 377253
rect 523915 377219 523949 377253
rect 523983 377219 524017 377253
rect 524051 377219 524085 377253
rect 524119 377219 524153 377253
rect 524187 377219 524221 377253
rect 524255 377219 524289 377253
rect 524323 377219 524357 377253
rect 524391 377219 524425 377253
rect 524459 377219 524493 377253
rect 524527 377219 524561 377253
rect 524595 377219 524629 377253
rect 524663 377219 524697 377253
rect 523439 376761 523473 376795
rect 523507 376761 523541 376795
rect 523575 376761 523609 376795
rect 523643 376761 523677 376795
rect 523711 376761 523745 376795
rect 523779 376761 523813 376795
rect 523847 376761 523881 376795
rect 523915 376761 523949 376795
rect 523983 376761 524017 376795
rect 524051 376761 524085 376795
rect 524119 376761 524153 376795
rect 524187 376761 524221 376795
rect 524255 376761 524289 376795
rect 524323 376761 524357 376795
rect 524391 376761 524425 376795
rect 524459 376761 524493 376795
rect 524527 376761 524561 376795
rect 524595 376761 524629 376795
rect 524663 376761 524697 376795
rect 523439 376303 523473 376337
rect 523507 376303 523541 376337
rect 523575 376303 523609 376337
rect 523643 376303 523677 376337
rect 523711 376303 523745 376337
rect 523779 376303 523813 376337
rect 523847 376303 523881 376337
rect 523915 376303 523949 376337
rect 523983 376303 524017 376337
rect 524051 376303 524085 376337
rect 524119 376303 524153 376337
rect 524187 376303 524221 376337
rect 524255 376303 524289 376337
rect 524323 376303 524357 376337
rect 524391 376303 524425 376337
rect 524459 376303 524493 376337
rect 524527 376303 524561 376337
rect 524595 376303 524629 376337
rect 524663 376303 524697 376337
rect 523439 375845 523473 375879
rect 523507 375845 523541 375879
rect 523575 375845 523609 375879
rect 523643 375845 523677 375879
rect 523711 375845 523745 375879
rect 523779 375845 523813 375879
rect 523847 375845 523881 375879
rect 523915 375845 523949 375879
rect 523983 375845 524017 375879
rect 524051 375845 524085 375879
rect 524119 375845 524153 375879
rect 524187 375845 524221 375879
rect 524255 375845 524289 375879
rect 524323 375845 524357 375879
rect 524391 375845 524425 375879
rect 524459 375845 524493 375879
rect 524527 375845 524561 375879
rect 524595 375845 524629 375879
rect 524663 375845 524697 375879
rect 523439 375387 523473 375421
rect 523507 375387 523541 375421
rect 523575 375387 523609 375421
rect 523643 375387 523677 375421
rect 523711 375387 523745 375421
rect 523779 375387 523813 375421
rect 523847 375387 523881 375421
rect 523915 375387 523949 375421
rect 523983 375387 524017 375421
rect 524051 375387 524085 375421
rect 524119 375387 524153 375421
rect 524187 375387 524221 375421
rect 524255 375387 524289 375421
rect 524323 375387 524357 375421
rect 524391 375387 524425 375421
rect 524459 375387 524493 375421
rect 524527 375387 524561 375421
rect 524595 375387 524629 375421
rect 524663 375387 524697 375421
rect 523439 374929 523473 374963
rect 523507 374929 523541 374963
rect 523575 374929 523609 374963
rect 523643 374929 523677 374963
rect 523711 374929 523745 374963
rect 523779 374929 523813 374963
rect 523847 374929 523881 374963
rect 523915 374929 523949 374963
rect 523983 374929 524017 374963
rect 524051 374929 524085 374963
rect 524119 374929 524153 374963
rect 524187 374929 524221 374963
rect 524255 374929 524289 374963
rect 524323 374929 524357 374963
rect 524391 374929 524425 374963
rect 524459 374929 524493 374963
rect 524527 374929 524561 374963
rect 524595 374929 524629 374963
rect 524663 374929 524697 374963
rect 512159 374653 512193 374687
rect 512227 374653 512261 374687
rect 512295 374653 512329 374687
rect 512363 374653 512397 374687
rect 512431 374653 512465 374687
rect 512499 374653 512533 374687
rect 512567 374653 512601 374687
rect 512635 374653 512669 374687
rect 512703 374653 512737 374687
rect 512771 374653 512805 374687
rect 512839 374653 512873 374687
rect 512907 374653 512941 374687
rect 512975 374653 513009 374687
rect 513043 374653 513077 374687
rect 513111 374653 513145 374687
rect 513179 374653 513213 374687
rect 513247 374653 513281 374687
rect 513315 374653 513349 374687
rect 513383 374653 513417 374687
rect 493359 373097 493393 373131
rect 493427 373097 493461 373131
rect 493495 373097 493529 373131
rect 493563 373097 493597 373131
rect 493631 373097 493665 373131
rect 493699 373097 493733 373131
rect 493767 373097 493801 373131
rect 493835 373097 493869 373131
rect 493903 373097 493937 373131
rect 493971 373097 494005 373131
rect 494039 373097 494073 373131
rect 494107 373097 494141 373131
rect 494175 373097 494209 373131
rect 494243 373097 494277 373131
rect 494311 373097 494345 373131
rect 494379 373097 494413 373131
rect 494447 373097 494481 373131
rect 494515 373097 494549 373131
rect 494583 373097 494617 373131
rect 497119 373279 497153 373313
rect 497187 373279 497221 373313
rect 497255 373279 497289 373313
rect 497323 373279 497357 373313
rect 497391 373279 497425 373313
rect 497459 373279 497493 373313
rect 497527 373279 497561 373313
rect 497595 373279 497629 373313
rect 497663 373279 497697 373313
rect 497731 373279 497765 373313
rect 497799 373279 497833 373313
rect 497867 373279 497901 373313
rect 497935 373279 497969 373313
rect 498003 373279 498037 373313
rect 498071 373279 498105 373313
rect 498139 373279 498173 373313
rect 498207 373279 498241 373313
rect 498275 373279 498309 373313
rect 498343 373279 498377 373313
rect 497119 372821 497153 372855
rect 497187 372821 497221 372855
rect 497255 372821 497289 372855
rect 497323 372821 497357 372855
rect 497391 372821 497425 372855
rect 497459 372821 497493 372855
rect 497527 372821 497561 372855
rect 497595 372821 497629 372855
rect 497663 372821 497697 372855
rect 497731 372821 497765 372855
rect 497799 372821 497833 372855
rect 497867 372821 497901 372855
rect 497935 372821 497969 372855
rect 498003 372821 498037 372855
rect 498071 372821 498105 372855
rect 498139 372821 498173 372855
rect 498207 372821 498241 372855
rect 498275 372821 498309 372855
rect 498343 372821 498377 372855
rect 493359 372639 493393 372673
rect 493427 372639 493461 372673
rect 493495 372639 493529 372673
rect 493563 372639 493597 372673
rect 493631 372639 493665 372673
rect 493699 372639 493733 372673
rect 493767 372639 493801 372673
rect 493835 372639 493869 372673
rect 493903 372639 493937 372673
rect 493971 372639 494005 372673
rect 494039 372639 494073 372673
rect 494107 372639 494141 372673
rect 494175 372639 494209 372673
rect 494243 372639 494277 372673
rect 494311 372639 494345 372673
rect 494379 372639 494413 372673
rect 494447 372639 494481 372673
rect 494515 372639 494549 372673
rect 494583 372639 494617 372673
rect 497119 372363 497153 372397
rect 497187 372363 497221 372397
rect 497255 372363 497289 372397
rect 497323 372363 497357 372397
rect 497391 372363 497425 372397
rect 497459 372363 497493 372397
rect 497527 372363 497561 372397
rect 497595 372363 497629 372397
rect 497663 372363 497697 372397
rect 497731 372363 497765 372397
rect 497799 372363 497833 372397
rect 497867 372363 497901 372397
rect 497935 372363 497969 372397
rect 498003 372363 498037 372397
rect 498071 372363 498105 372397
rect 498139 372363 498173 372397
rect 498207 372363 498241 372397
rect 498275 372363 498309 372397
rect 498343 372363 498377 372397
rect 493359 372181 493393 372215
rect 493427 372181 493461 372215
rect 493495 372181 493529 372215
rect 493563 372181 493597 372215
rect 493631 372181 493665 372215
rect 493699 372181 493733 372215
rect 493767 372181 493801 372215
rect 493835 372181 493869 372215
rect 493903 372181 493937 372215
rect 493971 372181 494005 372215
rect 494039 372181 494073 372215
rect 494107 372181 494141 372215
rect 494175 372181 494209 372215
rect 494243 372181 494277 372215
rect 494311 372181 494345 372215
rect 494379 372181 494413 372215
rect 494447 372181 494481 372215
rect 494515 372181 494549 372215
rect 494583 372181 494617 372215
rect 501280 372752 501314 372786
rect 501370 372752 501404 372786
rect 501460 372752 501494 372786
rect 501550 372752 501584 372786
rect 501640 372752 501674 372786
rect 501730 372752 501764 372786
rect 501820 372752 501854 372786
rect 501280 372662 501314 372696
rect 501370 372662 501404 372696
rect 501460 372662 501494 372696
rect 501550 372662 501584 372696
rect 501640 372662 501674 372696
rect 501730 372662 501764 372696
rect 501820 372662 501854 372696
rect 501280 372572 501314 372606
rect 501370 372572 501404 372606
rect 501460 372572 501494 372606
rect 501550 372572 501584 372606
rect 501640 372572 501674 372606
rect 501730 372572 501764 372606
rect 501820 372572 501854 372606
rect 501280 372482 501314 372516
rect 501370 372482 501404 372516
rect 501460 372482 501494 372516
rect 501550 372482 501584 372516
rect 501640 372482 501674 372516
rect 501730 372482 501764 372516
rect 501820 372482 501854 372516
rect 501280 372392 501314 372426
rect 501370 372392 501404 372426
rect 501460 372392 501494 372426
rect 501550 372392 501584 372426
rect 501640 372392 501674 372426
rect 501730 372392 501764 372426
rect 501820 372392 501854 372426
rect 501280 372302 501314 372336
rect 501370 372302 501404 372336
rect 501460 372302 501494 372336
rect 501550 372302 501584 372336
rect 501640 372302 501674 372336
rect 501730 372302 501764 372336
rect 501820 372302 501854 372336
rect 501280 372212 501314 372246
rect 501370 372212 501404 372246
rect 501460 372212 501494 372246
rect 501550 372212 501584 372246
rect 501640 372212 501674 372246
rect 501730 372212 501764 372246
rect 501820 372212 501854 372246
rect 493359 371723 493393 371757
rect 493427 371723 493461 371757
rect 493495 371723 493529 371757
rect 493563 371723 493597 371757
rect 493631 371723 493665 371757
rect 493699 371723 493733 371757
rect 493767 371723 493801 371757
rect 493835 371723 493869 371757
rect 493903 371723 493937 371757
rect 493971 371723 494005 371757
rect 494039 371723 494073 371757
rect 494107 371723 494141 371757
rect 494175 371723 494209 371757
rect 494243 371723 494277 371757
rect 494311 371723 494345 371757
rect 494379 371723 494413 371757
rect 494447 371723 494481 371757
rect 494515 371723 494549 371757
rect 494583 371723 494617 371757
rect 493359 371265 493393 371299
rect 493427 371265 493461 371299
rect 493495 371265 493529 371299
rect 493563 371265 493597 371299
rect 493631 371265 493665 371299
rect 493699 371265 493733 371299
rect 493767 371265 493801 371299
rect 493835 371265 493869 371299
rect 493903 371265 493937 371299
rect 493971 371265 494005 371299
rect 494039 371265 494073 371299
rect 494107 371265 494141 371299
rect 494175 371265 494209 371299
rect 494243 371265 494277 371299
rect 494311 371265 494345 371299
rect 494379 371265 494413 371299
rect 494447 371265 494481 371299
rect 494515 371265 494549 371299
rect 494583 371265 494617 371299
rect 493359 370807 493393 370841
rect 493427 370807 493461 370841
rect 493495 370807 493529 370841
rect 493563 370807 493597 370841
rect 493631 370807 493665 370841
rect 493699 370807 493733 370841
rect 493767 370807 493801 370841
rect 493835 370807 493869 370841
rect 493903 370807 493937 370841
rect 493971 370807 494005 370841
rect 494039 370807 494073 370841
rect 494107 370807 494141 370841
rect 494175 370807 494209 370841
rect 494243 370807 494277 370841
rect 494311 370807 494345 370841
rect 494379 370807 494413 370841
rect 494447 370807 494481 370841
rect 494515 370807 494549 370841
rect 494583 370807 494617 370841
rect 493359 370349 493393 370383
rect 493427 370349 493461 370383
rect 493495 370349 493529 370383
rect 493563 370349 493597 370383
rect 493631 370349 493665 370383
rect 493699 370349 493733 370383
rect 493767 370349 493801 370383
rect 493835 370349 493869 370383
rect 493903 370349 493937 370383
rect 493971 370349 494005 370383
rect 494039 370349 494073 370383
rect 494107 370349 494141 370383
rect 494175 370349 494209 370383
rect 494243 370349 494277 370383
rect 494311 370349 494345 370383
rect 494379 370349 494413 370383
rect 494447 370349 494481 370383
rect 494515 370349 494549 370383
rect 494583 370349 494617 370383
rect 493359 369891 493393 369925
rect 493427 369891 493461 369925
rect 493495 369891 493529 369925
rect 493563 369891 493597 369925
rect 493631 369891 493665 369925
rect 493699 369891 493733 369925
rect 493767 369891 493801 369925
rect 493835 369891 493869 369925
rect 493903 369891 493937 369925
rect 493971 369891 494005 369925
rect 494039 369891 494073 369925
rect 494107 369891 494141 369925
rect 494175 369891 494209 369925
rect 494243 369891 494277 369925
rect 494311 369891 494345 369925
rect 494379 369891 494413 369925
rect 494447 369891 494481 369925
rect 494515 369891 494549 369925
rect 494583 369891 494617 369925
rect 493359 369433 493393 369467
rect 493427 369433 493461 369467
rect 493495 369433 493529 369467
rect 493563 369433 493597 369467
rect 493631 369433 493665 369467
rect 493699 369433 493733 369467
rect 493767 369433 493801 369467
rect 493835 369433 493869 369467
rect 493903 369433 493937 369467
rect 493971 369433 494005 369467
rect 494039 369433 494073 369467
rect 494107 369433 494141 369467
rect 494175 369433 494209 369467
rect 494243 369433 494277 369467
rect 494311 369433 494345 369467
rect 494379 369433 494413 369467
rect 494447 369433 494481 369467
rect 494515 369433 494549 369467
rect 494583 369433 494617 369467
rect 493359 368975 493393 369009
rect 493427 368975 493461 369009
rect 493495 368975 493529 369009
rect 493563 368975 493597 369009
rect 493631 368975 493665 369009
rect 493699 368975 493733 369009
rect 493767 368975 493801 369009
rect 493835 368975 493869 369009
rect 493903 368975 493937 369009
rect 493971 368975 494005 369009
rect 494039 368975 494073 369009
rect 494107 368975 494141 369009
rect 494175 368975 494209 369009
rect 494243 368975 494277 369009
rect 494311 368975 494345 369009
rect 494379 368975 494413 369009
rect 494447 368975 494481 369009
rect 494515 368975 494549 369009
rect 494583 368975 494617 369009
rect 493359 368517 493393 368551
rect 493427 368517 493461 368551
rect 493495 368517 493529 368551
rect 493563 368517 493597 368551
rect 493631 368517 493665 368551
rect 493699 368517 493733 368551
rect 493767 368517 493801 368551
rect 493835 368517 493869 368551
rect 493903 368517 493937 368551
rect 493971 368517 494005 368551
rect 494039 368517 494073 368551
rect 494107 368517 494141 368551
rect 494175 368517 494209 368551
rect 494243 368517 494277 368551
rect 494311 368517 494345 368551
rect 494379 368517 494413 368551
rect 494447 368517 494481 368551
rect 494515 368517 494549 368551
rect 494583 368517 494617 368551
rect 493359 368059 493393 368093
rect 493427 368059 493461 368093
rect 493495 368059 493529 368093
rect 493563 368059 493597 368093
rect 493631 368059 493665 368093
rect 493699 368059 493733 368093
rect 493767 368059 493801 368093
rect 493835 368059 493869 368093
rect 493903 368059 493937 368093
rect 493971 368059 494005 368093
rect 494039 368059 494073 368093
rect 494107 368059 494141 368093
rect 494175 368059 494209 368093
rect 494243 368059 494277 368093
rect 494311 368059 494345 368093
rect 494379 368059 494413 368093
rect 494447 368059 494481 368093
rect 494515 368059 494549 368093
rect 494583 368059 494617 368093
rect 493359 367601 493393 367635
rect 493427 367601 493461 367635
rect 493495 367601 493529 367635
rect 493563 367601 493597 367635
rect 493631 367601 493665 367635
rect 493699 367601 493733 367635
rect 493767 367601 493801 367635
rect 493835 367601 493869 367635
rect 493903 367601 493937 367635
rect 493971 367601 494005 367635
rect 494039 367601 494073 367635
rect 494107 367601 494141 367635
rect 494175 367601 494209 367635
rect 494243 367601 494277 367635
rect 494311 367601 494345 367635
rect 494379 367601 494413 367635
rect 494447 367601 494481 367635
rect 494515 367601 494549 367635
rect 494583 367601 494617 367635
rect 493359 367143 493393 367177
rect 493427 367143 493461 367177
rect 493495 367143 493529 367177
rect 493563 367143 493597 367177
rect 493631 367143 493665 367177
rect 493699 367143 493733 367177
rect 493767 367143 493801 367177
rect 493835 367143 493869 367177
rect 493903 367143 493937 367177
rect 493971 367143 494005 367177
rect 494039 367143 494073 367177
rect 494107 367143 494141 367177
rect 494175 367143 494209 367177
rect 494243 367143 494277 367177
rect 494311 367143 494345 367177
rect 494379 367143 494413 367177
rect 494447 367143 494481 367177
rect 494515 367143 494549 367177
rect 494583 367143 494617 367177
rect 493359 366685 493393 366719
rect 493427 366685 493461 366719
rect 493495 366685 493529 366719
rect 493563 366685 493597 366719
rect 493631 366685 493665 366719
rect 493699 366685 493733 366719
rect 493767 366685 493801 366719
rect 493835 366685 493869 366719
rect 493903 366685 493937 366719
rect 493971 366685 494005 366719
rect 494039 366685 494073 366719
rect 494107 366685 494141 366719
rect 494175 366685 494209 366719
rect 494243 366685 494277 366719
rect 494311 366685 494345 366719
rect 494379 366685 494413 366719
rect 494447 366685 494481 366719
rect 494515 366685 494549 366719
rect 494583 366685 494617 366719
rect 493359 366227 493393 366261
rect 493427 366227 493461 366261
rect 493495 366227 493529 366261
rect 493563 366227 493597 366261
rect 493631 366227 493665 366261
rect 493699 366227 493733 366261
rect 493767 366227 493801 366261
rect 493835 366227 493869 366261
rect 493903 366227 493937 366261
rect 493971 366227 494005 366261
rect 494039 366227 494073 366261
rect 494107 366227 494141 366261
rect 494175 366227 494209 366261
rect 494243 366227 494277 366261
rect 494311 366227 494345 366261
rect 494379 366227 494413 366261
rect 494447 366227 494481 366261
rect 494515 366227 494549 366261
rect 494583 366227 494617 366261
rect 493359 365769 493393 365803
rect 493427 365769 493461 365803
rect 493495 365769 493529 365803
rect 493563 365769 493597 365803
rect 493631 365769 493665 365803
rect 493699 365769 493733 365803
rect 493767 365769 493801 365803
rect 493835 365769 493869 365803
rect 493903 365769 493937 365803
rect 493971 365769 494005 365803
rect 494039 365769 494073 365803
rect 494107 365769 494141 365803
rect 494175 365769 494209 365803
rect 494243 365769 494277 365803
rect 494311 365769 494345 365803
rect 494379 365769 494413 365803
rect 494447 365769 494481 365803
rect 494515 365769 494549 365803
rect 494583 365769 494617 365803
rect 493359 365311 493393 365345
rect 493427 365311 493461 365345
rect 493495 365311 493529 365345
rect 493563 365311 493597 365345
rect 493631 365311 493665 365345
rect 493699 365311 493733 365345
rect 493767 365311 493801 365345
rect 493835 365311 493869 365345
rect 493903 365311 493937 365345
rect 493971 365311 494005 365345
rect 494039 365311 494073 365345
rect 494107 365311 494141 365345
rect 494175 365311 494209 365345
rect 494243 365311 494277 365345
rect 494311 365311 494345 365345
rect 494379 365311 494413 365345
rect 494447 365311 494481 365345
rect 494515 365311 494549 365345
rect 494583 365311 494617 365345
rect 493359 364853 493393 364887
rect 493427 364853 493461 364887
rect 493495 364853 493529 364887
rect 493563 364853 493597 364887
rect 493631 364853 493665 364887
rect 493699 364853 493733 364887
rect 493767 364853 493801 364887
rect 493835 364853 493869 364887
rect 493903 364853 493937 364887
rect 493971 364853 494005 364887
rect 494039 364853 494073 364887
rect 494107 364853 494141 364887
rect 494175 364853 494209 364887
rect 494243 364853 494277 364887
rect 494311 364853 494345 364887
rect 494379 364853 494413 364887
rect 494447 364853 494481 364887
rect 494515 364853 494549 364887
rect 494583 364853 494617 364887
rect 493359 364395 493393 364429
rect 493427 364395 493461 364429
rect 493495 364395 493529 364429
rect 493563 364395 493597 364429
rect 493631 364395 493665 364429
rect 493699 364395 493733 364429
rect 493767 364395 493801 364429
rect 493835 364395 493869 364429
rect 493903 364395 493937 364429
rect 493971 364395 494005 364429
rect 494039 364395 494073 364429
rect 494107 364395 494141 364429
rect 494175 364395 494209 364429
rect 494243 364395 494277 364429
rect 494311 364395 494345 364429
rect 494379 364395 494413 364429
rect 494447 364395 494481 364429
rect 494515 364395 494549 364429
rect 494583 364395 494617 364429
rect 493359 363937 493393 363971
rect 493427 363937 493461 363971
rect 493495 363937 493529 363971
rect 493563 363937 493597 363971
rect 493631 363937 493665 363971
rect 493699 363937 493733 363971
rect 493767 363937 493801 363971
rect 493835 363937 493869 363971
rect 493903 363937 493937 363971
rect 493971 363937 494005 363971
rect 494039 363937 494073 363971
rect 494107 363937 494141 363971
rect 494175 363937 494209 363971
rect 494243 363937 494277 363971
rect 494311 363937 494345 363971
rect 494379 363937 494413 363971
rect 494447 363937 494481 363971
rect 494515 363937 494549 363971
rect 494583 363937 494617 363971
rect 493359 363479 493393 363513
rect 493427 363479 493461 363513
rect 493495 363479 493529 363513
rect 493563 363479 493597 363513
rect 493631 363479 493665 363513
rect 493699 363479 493733 363513
rect 493767 363479 493801 363513
rect 493835 363479 493869 363513
rect 493903 363479 493937 363513
rect 493971 363479 494005 363513
rect 494039 363479 494073 363513
rect 494107 363479 494141 363513
rect 494175 363479 494209 363513
rect 494243 363479 494277 363513
rect 494311 363479 494345 363513
rect 494379 363479 494413 363513
rect 494447 363479 494481 363513
rect 494515 363479 494549 363513
rect 494583 363479 494617 363513
rect 493359 363021 493393 363055
rect 493427 363021 493461 363055
rect 493495 363021 493529 363055
rect 493563 363021 493597 363055
rect 493631 363021 493665 363055
rect 493699 363021 493733 363055
rect 493767 363021 493801 363055
rect 493835 363021 493869 363055
rect 493903 363021 493937 363055
rect 493971 363021 494005 363055
rect 494039 363021 494073 363055
rect 494107 363021 494141 363055
rect 494175 363021 494209 363055
rect 494243 363021 494277 363055
rect 494311 363021 494345 363055
rect 494379 363021 494413 363055
rect 494447 363021 494481 363055
rect 494515 363021 494549 363055
rect 494583 363021 494617 363055
rect 493359 362563 493393 362597
rect 493427 362563 493461 362597
rect 493495 362563 493529 362597
rect 493563 362563 493597 362597
rect 493631 362563 493665 362597
rect 493699 362563 493733 362597
rect 493767 362563 493801 362597
rect 493835 362563 493869 362597
rect 493903 362563 493937 362597
rect 493971 362563 494005 362597
rect 494039 362563 494073 362597
rect 494107 362563 494141 362597
rect 494175 362563 494209 362597
rect 494243 362563 494277 362597
rect 494311 362563 494345 362597
rect 494379 362563 494413 362597
rect 494447 362563 494481 362597
rect 494515 362563 494549 362597
rect 494583 362563 494617 362597
rect 497520 371576 497554 371610
rect 497610 371576 497644 371610
rect 497700 371576 497734 371610
rect 497790 371576 497824 371610
rect 497880 371576 497914 371610
rect 497970 371576 498004 371610
rect 498060 371576 498094 371610
rect 497520 371486 497554 371520
rect 497610 371486 497644 371520
rect 497700 371486 497734 371520
rect 497790 371486 497824 371520
rect 497880 371486 497914 371520
rect 497970 371486 498004 371520
rect 498060 371486 498094 371520
rect 497520 371396 497554 371430
rect 497610 371396 497644 371430
rect 497700 371396 497734 371430
rect 497790 371396 497824 371430
rect 497880 371396 497914 371430
rect 497970 371396 498004 371430
rect 498060 371396 498094 371430
rect 497520 371306 497554 371340
rect 497610 371306 497644 371340
rect 497700 371306 497734 371340
rect 497790 371306 497824 371340
rect 497880 371306 497914 371340
rect 497970 371306 498004 371340
rect 498060 371306 498094 371340
rect 497520 371216 497554 371250
rect 497610 371216 497644 371250
rect 497700 371216 497734 371250
rect 497790 371216 497824 371250
rect 497880 371216 497914 371250
rect 497970 371216 498004 371250
rect 498060 371216 498094 371250
rect 497520 371126 497554 371160
rect 497610 371126 497644 371160
rect 497700 371126 497734 371160
rect 497790 371126 497824 371160
rect 497880 371126 497914 371160
rect 497970 371126 498004 371160
rect 498060 371126 498094 371160
rect 497520 371036 497554 371070
rect 497610 371036 497644 371070
rect 497700 371036 497734 371070
rect 497790 371036 497824 371070
rect 497880 371036 497914 371070
rect 497970 371036 498004 371070
rect 498060 371036 498094 371070
rect 497520 370236 497554 370270
rect 497610 370236 497644 370270
rect 497700 370236 497734 370270
rect 497790 370236 497824 370270
rect 497880 370236 497914 370270
rect 497970 370236 498004 370270
rect 498060 370236 498094 370270
rect 497520 370146 497554 370180
rect 497610 370146 497644 370180
rect 497700 370146 497734 370180
rect 497790 370146 497824 370180
rect 497880 370146 497914 370180
rect 497970 370146 498004 370180
rect 498060 370146 498094 370180
rect 497520 370056 497554 370090
rect 497610 370056 497644 370090
rect 497700 370056 497734 370090
rect 497790 370056 497824 370090
rect 497880 370056 497914 370090
rect 497970 370056 498004 370090
rect 498060 370056 498094 370090
rect 497520 369966 497554 370000
rect 497610 369966 497644 370000
rect 497700 369966 497734 370000
rect 497790 369966 497824 370000
rect 497880 369966 497914 370000
rect 497970 369966 498004 370000
rect 498060 369966 498094 370000
rect 497520 369876 497554 369910
rect 497610 369876 497644 369910
rect 497700 369876 497734 369910
rect 497790 369876 497824 369910
rect 497880 369876 497914 369910
rect 497970 369876 498004 369910
rect 498060 369876 498094 369910
rect 497520 369786 497554 369820
rect 497610 369786 497644 369820
rect 497700 369786 497734 369820
rect 497790 369786 497824 369820
rect 497880 369786 497914 369820
rect 497970 369786 498004 369820
rect 498060 369786 498094 369820
rect 497520 369696 497554 369730
rect 497610 369696 497644 369730
rect 497700 369696 497734 369730
rect 497790 369696 497824 369730
rect 497880 369696 497914 369730
rect 497970 369696 498004 369730
rect 498060 369696 498094 369730
rect 497520 368896 497554 368930
rect 497610 368896 497644 368930
rect 497700 368896 497734 368930
rect 497790 368896 497824 368930
rect 497880 368896 497914 368930
rect 497970 368896 498004 368930
rect 498060 368896 498094 368930
rect 497520 368806 497554 368840
rect 497610 368806 497644 368840
rect 497700 368806 497734 368840
rect 497790 368806 497824 368840
rect 497880 368806 497914 368840
rect 497970 368806 498004 368840
rect 498060 368806 498094 368840
rect 497520 368716 497554 368750
rect 497610 368716 497644 368750
rect 497700 368716 497734 368750
rect 497790 368716 497824 368750
rect 497880 368716 497914 368750
rect 497970 368716 498004 368750
rect 498060 368716 498094 368750
rect 497520 368626 497554 368660
rect 497610 368626 497644 368660
rect 497700 368626 497734 368660
rect 497790 368626 497824 368660
rect 497880 368626 497914 368660
rect 497970 368626 498004 368660
rect 498060 368626 498094 368660
rect 497520 368536 497554 368570
rect 497610 368536 497644 368570
rect 497700 368536 497734 368570
rect 497790 368536 497824 368570
rect 497880 368536 497914 368570
rect 497970 368536 498004 368570
rect 498060 368536 498094 368570
rect 497520 368446 497554 368480
rect 497610 368446 497644 368480
rect 497700 368446 497734 368480
rect 497790 368446 497824 368480
rect 497880 368446 497914 368480
rect 497970 368446 498004 368480
rect 498060 368446 498094 368480
rect 497520 368356 497554 368390
rect 497610 368356 497644 368390
rect 497700 368356 497734 368390
rect 497790 368356 497824 368390
rect 497880 368356 497914 368390
rect 497970 368356 498004 368390
rect 498060 368356 498094 368390
rect 497520 367556 497554 367590
rect 497610 367556 497644 367590
rect 497700 367556 497734 367590
rect 497790 367556 497824 367590
rect 497880 367556 497914 367590
rect 497970 367556 498004 367590
rect 498060 367556 498094 367590
rect 497520 367466 497554 367500
rect 497610 367466 497644 367500
rect 497700 367466 497734 367500
rect 497790 367466 497824 367500
rect 497880 367466 497914 367500
rect 497970 367466 498004 367500
rect 498060 367466 498094 367500
rect 497520 367376 497554 367410
rect 497610 367376 497644 367410
rect 497700 367376 497734 367410
rect 497790 367376 497824 367410
rect 497880 367376 497914 367410
rect 497970 367376 498004 367410
rect 498060 367376 498094 367410
rect 497520 367286 497554 367320
rect 497610 367286 497644 367320
rect 497700 367286 497734 367320
rect 497790 367286 497824 367320
rect 497880 367286 497914 367320
rect 497970 367286 498004 367320
rect 498060 367286 498094 367320
rect 497520 367196 497554 367230
rect 497610 367196 497644 367230
rect 497700 367196 497734 367230
rect 497790 367196 497824 367230
rect 497880 367196 497914 367230
rect 497970 367196 498004 367230
rect 498060 367196 498094 367230
rect 497520 367106 497554 367140
rect 497610 367106 497644 367140
rect 497700 367106 497734 367140
rect 497790 367106 497824 367140
rect 497880 367106 497914 367140
rect 497970 367106 498004 367140
rect 498060 367106 498094 367140
rect 497520 367016 497554 367050
rect 497610 367016 497644 367050
rect 497700 367016 497734 367050
rect 497790 367016 497824 367050
rect 497880 367016 497914 367050
rect 497970 367016 498004 367050
rect 498060 367016 498094 367050
rect 497520 366216 497554 366250
rect 497610 366216 497644 366250
rect 497700 366216 497734 366250
rect 497790 366216 497824 366250
rect 497880 366216 497914 366250
rect 497970 366216 498004 366250
rect 498060 366216 498094 366250
rect 497520 366126 497554 366160
rect 497610 366126 497644 366160
rect 497700 366126 497734 366160
rect 497790 366126 497824 366160
rect 497880 366126 497914 366160
rect 497970 366126 498004 366160
rect 498060 366126 498094 366160
rect 497520 366036 497554 366070
rect 497610 366036 497644 366070
rect 497700 366036 497734 366070
rect 497790 366036 497824 366070
rect 497880 366036 497914 366070
rect 497970 366036 498004 366070
rect 498060 366036 498094 366070
rect 497520 365946 497554 365980
rect 497610 365946 497644 365980
rect 497700 365946 497734 365980
rect 497790 365946 497824 365980
rect 497880 365946 497914 365980
rect 497970 365946 498004 365980
rect 498060 365946 498094 365980
rect 497520 365856 497554 365890
rect 497610 365856 497644 365890
rect 497700 365856 497734 365890
rect 497790 365856 497824 365890
rect 497880 365856 497914 365890
rect 497970 365856 498004 365890
rect 498060 365856 498094 365890
rect 497520 365766 497554 365800
rect 497610 365766 497644 365800
rect 497700 365766 497734 365800
rect 497790 365766 497824 365800
rect 497880 365766 497914 365800
rect 497970 365766 498004 365800
rect 498060 365766 498094 365800
rect 497520 365676 497554 365710
rect 497610 365676 497644 365710
rect 497700 365676 497734 365710
rect 497790 365676 497824 365710
rect 497880 365676 497914 365710
rect 497970 365676 498004 365710
rect 498060 365676 498094 365710
rect 497520 364876 497554 364910
rect 497610 364876 497644 364910
rect 497700 364876 497734 364910
rect 497790 364876 497824 364910
rect 497880 364876 497914 364910
rect 497970 364876 498004 364910
rect 498060 364876 498094 364910
rect 497520 364786 497554 364820
rect 497610 364786 497644 364820
rect 497700 364786 497734 364820
rect 497790 364786 497824 364820
rect 497880 364786 497914 364820
rect 497970 364786 498004 364820
rect 498060 364786 498094 364820
rect 497520 364696 497554 364730
rect 497610 364696 497644 364730
rect 497700 364696 497734 364730
rect 497790 364696 497824 364730
rect 497880 364696 497914 364730
rect 497970 364696 498004 364730
rect 498060 364696 498094 364730
rect 497520 364606 497554 364640
rect 497610 364606 497644 364640
rect 497700 364606 497734 364640
rect 497790 364606 497824 364640
rect 497880 364606 497914 364640
rect 497970 364606 498004 364640
rect 498060 364606 498094 364640
rect 497520 364516 497554 364550
rect 497610 364516 497644 364550
rect 497700 364516 497734 364550
rect 497790 364516 497824 364550
rect 497880 364516 497914 364550
rect 497970 364516 498004 364550
rect 498060 364516 498094 364550
rect 497520 364426 497554 364460
rect 497610 364426 497644 364460
rect 497700 364426 497734 364460
rect 497790 364426 497824 364460
rect 497880 364426 497914 364460
rect 497970 364426 498004 364460
rect 498060 364426 498094 364460
rect 497520 364336 497554 364370
rect 497610 364336 497644 364370
rect 497700 364336 497734 364370
rect 497790 364336 497824 364370
rect 497880 364336 497914 364370
rect 497970 364336 498004 364370
rect 498060 364336 498094 364370
rect 497520 363536 497554 363570
rect 497610 363536 497644 363570
rect 497700 363536 497734 363570
rect 497790 363536 497824 363570
rect 497880 363536 497914 363570
rect 497970 363536 498004 363570
rect 498060 363536 498094 363570
rect 497520 363446 497554 363480
rect 497610 363446 497644 363480
rect 497700 363446 497734 363480
rect 497790 363446 497824 363480
rect 497880 363446 497914 363480
rect 497970 363446 498004 363480
rect 498060 363446 498094 363480
rect 497520 363356 497554 363390
rect 497610 363356 497644 363390
rect 497700 363356 497734 363390
rect 497790 363356 497824 363390
rect 497880 363356 497914 363390
rect 497970 363356 498004 363390
rect 498060 363356 498094 363390
rect 497520 363266 497554 363300
rect 497610 363266 497644 363300
rect 497700 363266 497734 363300
rect 497790 363266 497824 363300
rect 497880 363266 497914 363300
rect 497970 363266 498004 363300
rect 498060 363266 498094 363300
rect 497520 363176 497554 363210
rect 497610 363176 497644 363210
rect 497700 363176 497734 363210
rect 497790 363176 497824 363210
rect 497880 363176 497914 363210
rect 497970 363176 498004 363210
rect 498060 363176 498094 363210
rect 497520 363086 497554 363120
rect 497610 363086 497644 363120
rect 497700 363086 497734 363120
rect 497790 363086 497824 363120
rect 497880 363086 497914 363120
rect 497970 363086 498004 363120
rect 498060 363086 498094 363120
rect 497520 362996 497554 363030
rect 497610 362996 497644 363030
rect 497700 362996 497734 363030
rect 497790 362996 497824 363030
rect 497880 362996 497914 363030
rect 497970 362996 498004 363030
rect 498060 362996 498094 363030
rect 501280 371412 501314 371446
rect 501370 371412 501404 371446
rect 501460 371412 501494 371446
rect 501550 371412 501584 371446
rect 501640 371412 501674 371446
rect 501730 371412 501764 371446
rect 501820 371412 501854 371446
rect 501280 371322 501314 371356
rect 501370 371322 501404 371356
rect 501460 371322 501494 371356
rect 501550 371322 501584 371356
rect 501640 371322 501674 371356
rect 501730 371322 501764 371356
rect 501820 371322 501854 371356
rect 501280 371232 501314 371266
rect 501370 371232 501404 371266
rect 501460 371232 501494 371266
rect 501550 371232 501584 371266
rect 501640 371232 501674 371266
rect 501730 371232 501764 371266
rect 501820 371232 501854 371266
rect 501280 371142 501314 371176
rect 501370 371142 501404 371176
rect 501460 371142 501494 371176
rect 501550 371142 501584 371176
rect 501640 371142 501674 371176
rect 501730 371142 501764 371176
rect 501820 371142 501854 371176
rect 501280 371052 501314 371086
rect 501370 371052 501404 371086
rect 501460 371052 501494 371086
rect 501550 371052 501584 371086
rect 501640 371052 501674 371086
rect 501730 371052 501764 371086
rect 501820 371052 501854 371086
rect 501280 370962 501314 370996
rect 501370 370962 501404 370996
rect 501460 370962 501494 370996
rect 501550 370962 501584 370996
rect 501640 370962 501674 370996
rect 501730 370962 501764 370996
rect 501820 370962 501854 370996
rect 501280 370872 501314 370906
rect 501370 370872 501404 370906
rect 501460 370872 501494 370906
rect 501550 370872 501584 370906
rect 501640 370872 501674 370906
rect 501730 370872 501764 370906
rect 501820 370872 501854 370906
rect 501280 370072 501314 370106
rect 501370 370072 501404 370106
rect 501460 370072 501494 370106
rect 501550 370072 501584 370106
rect 501640 370072 501674 370106
rect 501730 370072 501764 370106
rect 501820 370072 501854 370106
rect 501280 369982 501314 370016
rect 501370 369982 501404 370016
rect 501460 369982 501494 370016
rect 501550 369982 501584 370016
rect 501640 369982 501674 370016
rect 501730 369982 501764 370016
rect 501820 369982 501854 370016
rect 501280 369892 501314 369926
rect 501370 369892 501404 369926
rect 501460 369892 501494 369926
rect 501550 369892 501584 369926
rect 501640 369892 501674 369926
rect 501730 369892 501764 369926
rect 501820 369892 501854 369926
rect 501280 369802 501314 369836
rect 501370 369802 501404 369836
rect 501460 369802 501494 369836
rect 501550 369802 501584 369836
rect 501640 369802 501674 369836
rect 501730 369802 501764 369836
rect 501820 369802 501854 369836
rect 501280 369712 501314 369746
rect 501370 369712 501404 369746
rect 501460 369712 501494 369746
rect 501550 369712 501584 369746
rect 501640 369712 501674 369746
rect 501730 369712 501764 369746
rect 501820 369712 501854 369746
rect 501280 369622 501314 369656
rect 501370 369622 501404 369656
rect 501460 369622 501494 369656
rect 501550 369622 501584 369656
rect 501640 369622 501674 369656
rect 501730 369622 501764 369656
rect 501820 369622 501854 369656
rect 501280 369532 501314 369566
rect 501370 369532 501404 369566
rect 501460 369532 501494 369566
rect 501550 369532 501584 369566
rect 501640 369532 501674 369566
rect 501730 369532 501764 369566
rect 501820 369532 501854 369566
rect 501280 368732 501314 368766
rect 501370 368732 501404 368766
rect 501460 368732 501494 368766
rect 501550 368732 501584 368766
rect 501640 368732 501674 368766
rect 501730 368732 501764 368766
rect 501820 368732 501854 368766
rect 501280 368642 501314 368676
rect 501370 368642 501404 368676
rect 501460 368642 501494 368676
rect 501550 368642 501584 368676
rect 501640 368642 501674 368676
rect 501730 368642 501764 368676
rect 501820 368642 501854 368676
rect 501280 368552 501314 368586
rect 501370 368552 501404 368586
rect 501460 368552 501494 368586
rect 501550 368552 501584 368586
rect 501640 368552 501674 368586
rect 501730 368552 501764 368586
rect 501820 368552 501854 368586
rect 501280 368462 501314 368496
rect 501370 368462 501404 368496
rect 501460 368462 501494 368496
rect 501550 368462 501584 368496
rect 501640 368462 501674 368496
rect 501730 368462 501764 368496
rect 501820 368462 501854 368496
rect 501280 368372 501314 368406
rect 501370 368372 501404 368406
rect 501460 368372 501494 368406
rect 501550 368372 501584 368406
rect 501640 368372 501674 368406
rect 501730 368372 501764 368406
rect 501820 368372 501854 368406
rect 501280 368282 501314 368316
rect 501370 368282 501404 368316
rect 501460 368282 501494 368316
rect 501550 368282 501584 368316
rect 501640 368282 501674 368316
rect 501730 368282 501764 368316
rect 501820 368282 501854 368316
rect 501280 368192 501314 368226
rect 501370 368192 501404 368226
rect 501460 368192 501494 368226
rect 501550 368192 501584 368226
rect 501640 368192 501674 368226
rect 501730 368192 501764 368226
rect 501820 368192 501854 368226
rect 501280 367392 501314 367426
rect 501370 367392 501404 367426
rect 501460 367392 501494 367426
rect 501550 367392 501584 367426
rect 501640 367392 501674 367426
rect 501730 367392 501764 367426
rect 501820 367392 501854 367426
rect 501280 367302 501314 367336
rect 501370 367302 501404 367336
rect 501460 367302 501494 367336
rect 501550 367302 501584 367336
rect 501640 367302 501674 367336
rect 501730 367302 501764 367336
rect 501820 367302 501854 367336
rect 501280 367212 501314 367246
rect 501370 367212 501404 367246
rect 501460 367212 501494 367246
rect 501550 367212 501584 367246
rect 501640 367212 501674 367246
rect 501730 367212 501764 367246
rect 501820 367212 501854 367246
rect 501280 367122 501314 367156
rect 501370 367122 501404 367156
rect 501460 367122 501494 367156
rect 501550 367122 501584 367156
rect 501640 367122 501674 367156
rect 501730 367122 501764 367156
rect 501820 367122 501854 367156
rect 501280 367032 501314 367066
rect 501370 367032 501404 367066
rect 501460 367032 501494 367066
rect 501550 367032 501584 367066
rect 501640 367032 501674 367066
rect 501730 367032 501764 367066
rect 501820 367032 501854 367066
rect 501280 366942 501314 366976
rect 501370 366942 501404 366976
rect 501460 366942 501494 366976
rect 501550 366942 501584 366976
rect 501640 366942 501674 366976
rect 501730 366942 501764 366976
rect 501820 366942 501854 366976
rect 501280 366852 501314 366886
rect 501370 366852 501404 366886
rect 501460 366852 501494 366886
rect 501550 366852 501584 366886
rect 501640 366852 501674 366886
rect 501730 366852 501764 366886
rect 501820 366852 501854 366886
rect 501280 366052 501314 366086
rect 501370 366052 501404 366086
rect 501460 366052 501494 366086
rect 501550 366052 501584 366086
rect 501640 366052 501674 366086
rect 501730 366052 501764 366086
rect 501820 366052 501854 366086
rect 501280 365962 501314 365996
rect 501370 365962 501404 365996
rect 501460 365962 501494 365996
rect 501550 365962 501584 365996
rect 501640 365962 501674 365996
rect 501730 365962 501764 365996
rect 501820 365962 501854 365996
rect 501280 365872 501314 365906
rect 501370 365872 501404 365906
rect 501460 365872 501494 365906
rect 501550 365872 501584 365906
rect 501640 365872 501674 365906
rect 501730 365872 501764 365906
rect 501820 365872 501854 365906
rect 501280 365782 501314 365816
rect 501370 365782 501404 365816
rect 501460 365782 501494 365816
rect 501550 365782 501584 365816
rect 501640 365782 501674 365816
rect 501730 365782 501764 365816
rect 501820 365782 501854 365816
rect 501280 365692 501314 365726
rect 501370 365692 501404 365726
rect 501460 365692 501494 365726
rect 501550 365692 501584 365726
rect 501640 365692 501674 365726
rect 501730 365692 501764 365726
rect 501820 365692 501854 365726
rect 501280 365602 501314 365636
rect 501370 365602 501404 365636
rect 501460 365602 501494 365636
rect 501550 365602 501584 365636
rect 501640 365602 501674 365636
rect 501730 365602 501764 365636
rect 501820 365602 501854 365636
rect 501280 365512 501314 365546
rect 501370 365512 501404 365546
rect 501460 365512 501494 365546
rect 501550 365512 501584 365546
rect 501640 365512 501674 365546
rect 501730 365512 501764 365546
rect 501820 365512 501854 365546
rect 501280 364712 501314 364746
rect 501370 364712 501404 364746
rect 501460 364712 501494 364746
rect 501550 364712 501584 364746
rect 501640 364712 501674 364746
rect 501730 364712 501764 364746
rect 501820 364712 501854 364746
rect 501280 364622 501314 364656
rect 501370 364622 501404 364656
rect 501460 364622 501494 364656
rect 501550 364622 501584 364656
rect 501640 364622 501674 364656
rect 501730 364622 501764 364656
rect 501820 364622 501854 364656
rect 501280 364532 501314 364566
rect 501370 364532 501404 364566
rect 501460 364532 501494 364566
rect 501550 364532 501584 364566
rect 501640 364532 501674 364566
rect 501730 364532 501764 364566
rect 501820 364532 501854 364566
rect 501280 364442 501314 364476
rect 501370 364442 501404 364476
rect 501460 364442 501494 364476
rect 501550 364442 501584 364476
rect 501640 364442 501674 364476
rect 501730 364442 501764 364476
rect 501820 364442 501854 364476
rect 501280 364352 501314 364386
rect 501370 364352 501404 364386
rect 501460 364352 501494 364386
rect 501550 364352 501584 364386
rect 501640 364352 501674 364386
rect 501730 364352 501764 364386
rect 501820 364352 501854 364386
rect 501280 364262 501314 364296
rect 501370 364262 501404 364296
rect 501460 364262 501494 364296
rect 501550 364262 501584 364296
rect 501640 364262 501674 364296
rect 501730 364262 501764 364296
rect 501820 364262 501854 364296
rect 501280 364172 501314 364206
rect 501370 364172 501404 364206
rect 501460 364172 501494 364206
rect 501550 364172 501584 364206
rect 501640 364172 501674 364206
rect 501730 364172 501764 364206
rect 501820 364172 501854 364206
rect 501280 363372 501314 363406
rect 501370 363372 501404 363406
rect 501460 363372 501494 363406
rect 501550 363372 501584 363406
rect 501640 363372 501674 363406
rect 501730 363372 501764 363406
rect 501820 363372 501854 363406
rect 501280 363282 501314 363316
rect 501370 363282 501404 363316
rect 501460 363282 501494 363316
rect 501550 363282 501584 363316
rect 501640 363282 501674 363316
rect 501730 363282 501764 363316
rect 501820 363282 501854 363316
rect 501280 363192 501314 363226
rect 501370 363192 501404 363226
rect 501460 363192 501494 363226
rect 501550 363192 501584 363226
rect 501640 363192 501674 363226
rect 501730 363192 501764 363226
rect 501820 363192 501854 363226
rect 501280 363102 501314 363136
rect 501370 363102 501404 363136
rect 501460 363102 501494 363136
rect 501550 363102 501584 363136
rect 501640 363102 501674 363136
rect 501730 363102 501764 363136
rect 501820 363102 501854 363136
rect 501280 363012 501314 363046
rect 501370 363012 501404 363046
rect 501460 363012 501494 363046
rect 501550 363012 501584 363046
rect 501640 363012 501674 363046
rect 501730 363012 501764 363046
rect 501820 363012 501854 363046
rect 501280 362922 501314 362956
rect 501370 362922 501404 362956
rect 501460 362922 501494 362956
rect 501550 362922 501584 362956
rect 501640 362922 501674 362956
rect 501730 362922 501764 362956
rect 501820 362922 501854 362956
rect 501280 362832 501314 362866
rect 501370 362832 501404 362866
rect 501460 362832 501494 362866
rect 501550 362832 501584 362866
rect 501640 362832 501674 362866
rect 501730 362832 501764 362866
rect 501820 362832 501854 362866
rect 505040 372752 505074 372786
rect 505130 372752 505164 372786
rect 505220 372752 505254 372786
rect 505310 372752 505344 372786
rect 505400 372752 505434 372786
rect 505490 372752 505524 372786
rect 505580 372752 505614 372786
rect 505040 372662 505074 372696
rect 505130 372662 505164 372696
rect 505220 372662 505254 372696
rect 505310 372662 505344 372696
rect 505400 372662 505434 372696
rect 505490 372662 505524 372696
rect 505580 372662 505614 372696
rect 505040 372572 505074 372606
rect 505130 372572 505164 372606
rect 505220 372572 505254 372606
rect 505310 372572 505344 372606
rect 505400 372572 505434 372606
rect 505490 372572 505524 372606
rect 505580 372572 505614 372606
rect 505040 372482 505074 372516
rect 505130 372482 505164 372516
rect 505220 372482 505254 372516
rect 505310 372482 505344 372516
rect 505400 372482 505434 372516
rect 505490 372482 505524 372516
rect 505580 372482 505614 372516
rect 505040 372392 505074 372426
rect 505130 372392 505164 372426
rect 505220 372392 505254 372426
rect 505310 372392 505344 372426
rect 505400 372392 505434 372426
rect 505490 372392 505524 372426
rect 505580 372392 505614 372426
rect 505040 372302 505074 372336
rect 505130 372302 505164 372336
rect 505220 372302 505254 372336
rect 505310 372302 505344 372336
rect 505400 372302 505434 372336
rect 505490 372302 505524 372336
rect 505580 372302 505614 372336
rect 505040 372212 505074 372246
rect 505130 372212 505164 372246
rect 505220 372212 505254 372246
rect 505310 372212 505344 372246
rect 505400 372212 505434 372246
rect 505490 372212 505524 372246
rect 505580 372212 505614 372246
rect 505040 371412 505074 371446
rect 505130 371412 505164 371446
rect 505220 371412 505254 371446
rect 505310 371412 505344 371446
rect 505400 371412 505434 371446
rect 505490 371412 505524 371446
rect 505580 371412 505614 371446
rect 505040 371322 505074 371356
rect 505130 371322 505164 371356
rect 505220 371322 505254 371356
rect 505310 371322 505344 371356
rect 505400 371322 505434 371356
rect 505490 371322 505524 371356
rect 505580 371322 505614 371356
rect 505040 371232 505074 371266
rect 505130 371232 505164 371266
rect 505220 371232 505254 371266
rect 505310 371232 505344 371266
rect 505400 371232 505434 371266
rect 505490 371232 505524 371266
rect 505580 371232 505614 371266
rect 505040 371142 505074 371176
rect 505130 371142 505164 371176
rect 505220 371142 505254 371176
rect 505310 371142 505344 371176
rect 505400 371142 505434 371176
rect 505490 371142 505524 371176
rect 505580 371142 505614 371176
rect 505040 371052 505074 371086
rect 505130 371052 505164 371086
rect 505220 371052 505254 371086
rect 505310 371052 505344 371086
rect 505400 371052 505434 371086
rect 505490 371052 505524 371086
rect 505580 371052 505614 371086
rect 505040 370962 505074 370996
rect 505130 370962 505164 370996
rect 505220 370962 505254 370996
rect 505310 370962 505344 370996
rect 505400 370962 505434 370996
rect 505490 370962 505524 370996
rect 505580 370962 505614 370996
rect 505040 370872 505074 370906
rect 505130 370872 505164 370906
rect 505220 370872 505254 370906
rect 505310 370872 505344 370906
rect 505400 370872 505434 370906
rect 505490 370872 505524 370906
rect 505580 370872 505614 370906
rect 505040 370072 505074 370106
rect 505130 370072 505164 370106
rect 505220 370072 505254 370106
rect 505310 370072 505344 370106
rect 505400 370072 505434 370106
rect 505490 370072 505524 370106
rect 505580 370072 505614 370106
rect 505040 369982 505074 370016
rect 505130 369982 505164 370016
rect 505220 369982 505254 370016
rect 505310 369982 505344 370016
rect 505400 369982 505434 370016
rect 505490 369982 505524 370016
rect 505580 369982 505614 370016
rect 505040 369892 505074 369926
rect 505130 369892 505164 369926
rect 505220 369892 505254 369926
rect 505310 369892 505344 369926
rect 505400 369892 505434 369926
rect 505490 369892 505524 369926
rect 505580 369892 505614 369926
rect 505040 369802 505074 369836
rect 505130 369802 505164 369836
rect 505220 369802 505254 369836
rect 505310 369802 505344 369836
rect 505400 369802 505434 369836
rect 505490 369802 505524 369836
rect 505580 369802 505614 369836
rect 505040 369712 505074 369746
rect 505130 369712 505164 369746
rect 505220 369712 505254 369746
rect 505310 369712 505344 369746
rect 505400 369712 505434 369746
rect 505490 369712 505524 369746
rect 505580 369712 505614 369746
rect 505040 369622 505074 369656
rect 505130 369622 505164 369656
rect 505220 369622 505254 369656
rect 505310 369622 505344 369656
rect 505400 369622 505434 369656
rect 505490 369622 505524 369656
rect 505580 369622 505614 369656
rect 505040 369532 505074 369566
rect 505130 369532 505164 369566
rect 505220 369532 505254 369566
rect 505310 369532 505344 369566
rect 505400 369532 505434 369566
rect 505490 369532 505524 369566
rect 505580 369532 505614 369566
rect 505040 368732 505074 368766
rect 505130 368732 505164 368766
rect 505220 368732 505254 368766
rect 505310 368732 505344 368766
rect 505400 368732 505434 368766
rect 505490 368732 505524 368766
rect 505580 368732 505614 368766
rect 505040 368642 505074 368676
rect 505130 368642 505164 368676
rect 505220 368642 505254 368676
rect 505310 368642 505344 368676
rect 505400 368642 505434 368676
rect 505490 368642 505524 368676
rect 505580 368642 505614 368676
rect 505040 368552 505074 368586
rect 505130 368552 505164 368586
rect 505220 368552 505254 368586
rect 505310 368552 505344 368586
rect 505400 368552 505434 368586
rect 505490 368552 505524 368586
rect 505580 368552 505614 368586
rect 505040 368462 505074 368496
rect 505130 368462 505164 368496
rect 505220 368462 505254 368496
rect 505310 368462 505344 368496
rect 505400 368462 505434 368496
rect 505490 368462 505524 368496
rect 505580 368462 505614 368496
rect 505040 368372 505074 368406
rect 505130 368372 505164 368406
rect 505220 368372 505254 368406
rect 505310 368372 505344 368406
rect 505400 368372 505434 368406
rect 505490 368372 505524 368406
rect 505580 368372 505614 368406
rect 505040 368282 505074 368316
rect 505130 368282 505164 368316
rect 505220 368282 505254 368316
rect 505310 368282 505344 368316
rect 505400 368282 505434 368316
rect 505490 368282 505524 368316
rect 505580 368282 505614 368316
rect 505040 368192 505074 368226
rect 505130 368192 505164 368226
rect 505220 368192 505254 368226
rect 505310 368192 505344 368226
rect 505400 368192 505434 368226
rect 505490 368192 505524 368226
rect 505580 368192 505614 368226
rect 505040 367392 505074 367426
rect 505130 367392 505164 367426
rect 505220 367392 505254 367426
rect 505310 367392 505344 367426
rect 505400 367392 505434 367426
rect 505490 367392 505524 367426
rect 505580 367392 505614 367426
rect 505040 367302 505074 367336
rect 505130 367302 505164 367336
rect 505220 367302 505254 367336
rect 505310 367302 505344 367336
rect 505400 367302 505434 367336
rect 505490 367302 505524 367336
rect 505580 367302 505614 367336
rect 505040 367212 505074 367246
rect 505130 367212 505164 367246
rect 505220 367212 505254 367246
rect 505310 367212 505344 367246
rect 505400 367212 505434 367246
rect 505490 367212 505524 367246
rect 505580 367212 505614 367246
rect 505040 367122 505074 367156
rect 505130 367122 505164 367156
rect 505220 367122 505254 367156
rect 505310 367122 505344 367156
rect 505400 367122 505434 367156
rect 505490 367122 505524 367156
rect 505580 367122 505614 367156
rect 505040 367032 505074 367066
rect 505130 367032 505164 367066
rect 505220 367032 505254 367066
rect 505310 367032 505344 367066
rect 505400 367032 505434 367066
rect 505490 367032 505524 367066
rect 505580 367032 505614 367066
rect 505040 366942 505074 366976
rect 505130 366942 505164 366976
rect 505220 366942 505254 366976
rect 505310 366942 505344 366976
rect 505400 366942 505434 366976
rect 505490 366942 505524 366976
rect 505580 366942 505614 366976
rect 505040 366852 505074 366886
rect 505130 366852 505164 366886
rect 505220 366852 505254 366886
rect 505310 366852 505344 366886
rect 505400 366852 505434 366886
rect 505490 366852 505524 366886
rect 505580 366852 505614 366886
rect 505040 366052 505074 366086
rect 505130 366052 505164 366086
rect 505220 366052 505254 366086
rect 505310 366052 505344 366086
rect 505400 366052 505434 366086
rect 505490 366052 505524 366086
rect 505580 366052 505614 366086
rect 505040 365962 505074 365996
rect 505130 365962 505164 365996
rect 505220 365962 505254 365996
rect 505310 365962 505344 365996
rect 505400 365962 505434 365996
rect 505490 365962 505524 365996
rect 505580 365962 505614 365996
rect 505040 365872 505074 365906
rect 505130 365872 505164 365906
rect 505220 365872 505254 365906
rect 505310 365872 505344 365906
rect 505400 365872 505434 365906
rect 505490 365872 505524 365906
rect 505580 365872 505614 365906
rect 505040 365782 505074 365816
rect 505130 365782 505164 365816
rect 505220 365782 505254 365816
rect 505310 365782 505344 365816
rect 505400 365782 505434 365816
rect 505490 365782 505524 365816
rect 505580 365782 505614 365816
rect 505040 365692 505074 365726
rect 505130 365692 505164 365726
rect 505220 365692 505254 365726
rect 505310 365692 505344 365726
rect 505400 365692 505434 365726
rect 505490 365692 505524 365726
rect 505580 365692 505614 365726
rect 505040 365602 505074 365636
rect 505130 365602 505164 365636
rect 505220 365602 505254 365636
rect 505310 365602 505344 365636
rect 505400 365602 505434 365636
rect 505490 365602 505524 365636
rect 505580 365602 505614 365636
rect 505040 365512 505074 365546
rect 505130 365512 505164 365546
rect 505220 365512 505254 365546
rect 505310 365512 505344 365546
rect 505400 365512 505434 365546
rect 505490 365512 505524 365546
rect 505580 365512 505614 365546
rect 505040 364712 505074 364746
rect 505130 364712 505164 364746
rect 505220 364712 505254 364746
rect 505310 364712 505344 364746
rect 505400 364712 505434 364746
rect 505490 364712 505524 364746
rect 505580 364712 505614 364746
rect 505040 364622 505074 364656
rect 505130 364622 505164 364656
rect 505220 364622 505254 364656
rect 505310 364622 505344 364656
rect 505400 364622 505434 364656
rect 505490 364622 505524 364656
rect 505580 364622 505614 364656
rect 505040 364532 505074 364566
rect 505130 364532 505164 364566
rect 505220 364532 505254 364566
rect 505310 364532 505344 364566
rect 505400 364532 505434 364566
rect 505490 364532 505524 364566
rect 505580 364532 505614 364566
rect 505040 364442 505074 364476
rect 505130 364442 505164 364476
rect 505220 364442 505254 364476
rect 505310 364442 505344 364476
rect 505400 364442 505434 364476
rect 505490 364442 505524 364476
rect 505580 364442 505614 364476
rect 505040 364352 505074 364386
rect 505130 364352 505164 364386
rect 505220 364352 505254 364386
rect 505310 364352 505344 364386
rect 505400 364352 505434 364386
rect 505490 364352 505524 364386
rect 505580 364352 505614 364386
rect 505040 364262 505074 364296
rect 505130 364262 505164 364296
rect 505220 364262 505254 364296
rect 505310 364262 505344 364296
rect 505400 364262 505434 364296
rect 505490 364262 505524 364296
rect 505580 364262 505614 364296
rect 505040 364172 505074 364206
rect 505130 364172 505164 364206
rect 505220 364172 505254 364206
rect 505310 364172 505344 364206
rect 505400 364172 505434 364206
rect 505490 364172 505524 364206
rect 505580 364172 505614 364206
rect 505040 363372 505074 363406
rect 505130 363372 505164 363406
rect 505220 363372 505254 363406
rect 505310 363372 505344 363406
rect 505400 363372 505434 363406
rect 505490 363372 505524 363406
rect 505580 363372 505614 363406
rect 505040 363282 505074 363316
rect 505130 363282 505164 363316
rect 505220 363282 505254 363316
rect 505310 363282 505344 363316
rect 505400 363282 505434 363316
rect 505490 363282 505524 363316
rect 505580 363282 505614 363316
rect 505040 363192 505074 363226
rect 505130 363192 505164 363226
rect 505220 363192 505254 363226
rect 505310 363192 505344 363226
rect 505400 363192 505434 363226
rect 505490 363192 505524 363226
rect 505580 363192 505614 363226
rect 505040 363102 505074 363136
rect 505130 363102 505164 363136
rect 505220 363102 505254 363136
rect 505310 363102 505344 363136
rect 505400 363102 505434 363136
rect 505490 363102 505524 363136
rect 505580 363102 505614 363136
rect 505040 363012 505074 363046
rect 505130 363012 505164 363046
rect 505220 363012 505254 363046
rect 505310 363012 505344 363046
rect 505400 363012 505434 363046
rect 505490 363012 505524 363046
rect 505580 363012 505614 363046
rect 505040 362922 505074 362956
rect 505130 362922 505164 362956
rect 505220 362922 505254 362956
rect 505310 362922 505344 362956
rect 505400 362922 505434 362956
rect 505490 362922 505524 362956
rect 505580 362922 505614 362956
rect 505040 362832 505074 362866
rect 505130 362832 505164 362866
rect 505220 362832 505254 362866
rect 505310 362832 505344 362866
rect 505400 362832 505434 362866
rect 505490 362832 505524 362866
rect 505580 362832 505614 362866
rect 508800 372752 508834 372786
rect 508890 372752 508924 372786
rect 508980 372752 509014 372786
rect 509070 372752 509104 372786
rect 509160 372752 509194 372786
rect 509250 372752 509284 372786
rect 509340 372752 509374 372786
rect 508800 372662 508834 372696
rect 508890 372662 508924 372696
rect 508980 372662 509014 372696
rect 509070 372662 509104 372696
rect 509160 372662 509194 372696
rect 509250 372662 509284 372696
rect 509340 372662 509374 372696
rect 508800 372572 508834 372606
rect 508890 372572 508924 372606
rect 508980 372572 509014 372606
rect 509070 372572 509104 372606
rect 509160 372572 509194 372606
rect 509250 372572 509284 372606
rect 509340 372572 509374 372606
rect 508800 372482 508834 372516
rect 508890 372482 508924 372516
rect 508980 372482 509014 372516
rect 509070 372482 509104 372516
rect 509160 372482 509194 372516
rect 509250 372482 509284 372516
rect 509340 372482 509374 372516
rect 508800 372392 508834 372426
rect 508890 372392 508924 372426
rect 508980 372392 509014 372426
rect 509070 372392 509104 372426
rect 509160 372392 509194 372426
rect 509250 372392 509284 372426
rect 509340 372392 509374 372426
rect 508800 372302 508834 372336
rect 508890 372302 508924 372336
rect 508980 372302 509014 372336
rect 509070 372302 509104 372336
rect 509160 372302 509194 372336
rect 509250 372302 509284 372336
rect 509340 372302 509374 372336
rect 508800 372212 508834 372246
rect 508890 372212 508924 372246
rect 508980 372212 509014 372246
rect 509070 372212 509104 372246
rect 509160 372212 509194 372246
rect 509250 372212 509284 372246
rect 509340 372212 509374 372246
rect 508800 371412 508834 371446
rect 508890 371412 508924 371446
rect 508980 371412 509014 371446
rect 509070 371412 509104 371446
rect 509160 371412 509194 371446
rect 509250 371412 509284 371446
rect 509340 371412 509374 371446
rect 508800 371322 508834 371356
rect 508890 371322 508924 371356
rect 508980 371322 509014 371356
rect 509070 371322 509104 371356
rect 509160 371322 509194 371356
rect 509250 371322 509284 371356
rect 509340 371322 509374 371356
rect 508800 371232 508834 371266
rect 508890 371232 508924 371266
rect 508980 371232 509014 371266
rect 509070 371232 509104 371266
rect 509160 371232 509194 371266
rect 509250 371232 509284 371266
rect 509340 371232 509374 371266
rect 508800 371142 508834 371176
rect 508890 371142 508924 371176
rect 508980 371142 509014 371176
rect 509070 371142 509104 371176
rect 509160 371142 509194 371176
rect 509250 371142 509284 371176
rect 509340 371142 509374 371176
rect 508800 371052 508834 371086
rect 508890 371052 508924 371086
rect 508980 371052 509014 371086
rect 509070 371052 509104 371086
rect 509160 371052 509194 371086
rect 509250 371052 509284 371086
rect 509340 371052 509374 371086
rect 508800 370962 508834 370996
rect 508890 370962 508924 370996
rect 508980 370962 509014 370996
rect 509070 370962 509104 370996
rect 509160 370962 509194 370996
rect 509250 370962 509284 370996
rect 509340 370962 509374 370996
rect 508800 370872 508834 370906
rect 508890 370872 508924 370906
rect 508980 370872 509014 370906
rect 509070 370872 509104 370906
rect 509160 370872 509194 370906
rect 509250 370872 509284 370906
rect 509340 370872 509374 370906
rect 508800 370072 508834 370106
rect 508890 370072 508924 370106
rect 508980 370072 509014 370106
rect 509070 370072 509104 370106
rect 509160 370072 509194 370106
rect 509250 370072 509284 370106
rect 509340 370072 509374 370106
rect 508800 369982 508834 370016
rect 508890 369982 508924 370016
rect 508980 369982 509014 370016
rect 509070 369982 509104 370016
rect 509160 369982 509194 370016
rect 509250 369982 509284 370016
rect 509340 369982 509374 370016
rect 508800 369892 508834 369926
rect 508890 369892 508924 369926
rect 508980 369892 509014 369926
rect 509070 369892 509104 369926
rect 509160 369892 509194 369926
rect 509250 369892 509284 369926
rect 509340 369892 509374 369926
rect 508800 369802 508834 369836
rect 508890 369802 508924 369836
rect 508980 369802 509014 369836
rect 509070 369802 509104 369836
rect 509160 369802 509194 369836
rect 509250 369802 509284 369836
rect 509340 369802 509374 369836
rect 508800 369712 508834 369746
rect 508890 369712 508924 369746
rect 508980 369712 509014 369746
rect 509070 369712 509104 369746
rect 509160 369712 509194 369746
rect 509250 369712 509284 369746
rect 509340 369712 509374 369746
rect 508800 369622 508834 369656
rect 508890 369622 508924 369656
rect 508980 369622 509014 369656
rect 509070 369622 509104 369656
rect 509160 369622 509194 369656
rect 509250 369622 509284 369656
rect 509340 369622 509374 369656
rect 508800 369532 508834 369566
rect 508890 369532 508924 369566
rect 508980 369532 509014 369566
rect 509070 369532 509104 369566
rect 509160 369532 509194 369566
rect 509250 369532 509284 369566
rect 509340 369532 509374 369566
rect 508800 368732 508834 368766
rect 508890 368732 508924 368766
rect 508980 368732 509014 368766
rect 509070 368732 509104 368766
rect 509160 368732 509194 368766
rect 509250 368732 509284 368766
rect 509340 368732 509374 368766
rect 508800 368642 508834 368676
rect 508890 368642 508924 368676
rect 508980 368642 509014 368676
rect 509070 368642 509104 368676
rect 509160 368642 509194 368676
rect 509250 368642 509284 368676
rect 509340 368642 509374 368676
rect 508800 368552 508834 368586
rect 508890 368552 508924 368586
rect 508980 368552 509014 368586
rect 509070 368552 509104 368586
rect 509160 368552 509194 368586
rect 509250 368552 509284 368586
rect 509340 368552 509374 368586
rect 508800 368462 508834 368496
rect 508890 368462 508924 368496
rect 508980 368462 509014 368496
rect 509070 368462 509104 368496
rect 509160 368462 509194 368496
rect 509250 368462 509284 368496
rect 509340 368462 509374 368496
rect 508800 368372 508834 368406
rect 508890 368372 508924 368406
rect 508980 368372 509014 368406
rect 509070 368372 509104 368406
rect 509160 368372 509194 368406
rect 509250 368372 509284 368406
rect 509340 368372 509374 368406
rect 508800 368282 508834 368316
rect 508890 368282 508924 368316
rect 508980 368282 509014 368316
rect 509070 368282 509104 368316
rect 509160 368282 509194 368316
rect 509250 368282 509284 368316
rect 509340 368282 509374 368316
rect 508800 368192 508834 368226
rect 508890 368192 508924 368226
rect 508980 368192 509014 368226
rect 509070 368192 509104 368226
rect 509160 368192 509194 368226
rect 509250 368192 509284 368226
rect 509340 368192 509374 368226
rect 508800 367392 508834 367426
rect 508890 367392 508924 367426
rect 508980 367392 509014 367426
rect 509070 367392 509104 367426
rect 509160 367392 509194 367426
rect 509250 367392 509284 367426
rect 509340 367392 509374 367426
rect 508800 367302 508834 367336
rect 508890 367302 508924 367336
rect 508980 367302 509014 367336
rect 509070 367302 509104 367336
rect 509160 367302 509194 367336
rect 509250 367302 509284 367336
rect 509340 367302 509374 367336
rect 508800 367212 508834 367246
rect 508890 367212 508924 367246
rect 508980 367212 509014 367246
rect 509070 367212 509104 367246
rect 509160 367212 509194 367246
rect 509250 367212 509284 367246
rect 509340 367212 509374 367246
rect 508800 367122 508834 367156
rect 508890 367122 508924 367156
rect 508980 367122 509014 367156
rect 509070 367122 509104 367156
rect 509160 367122 509194 367156
rect 509250 367122 509284 367156
rect 509340 367122 509374 367156
rect 508800 367032 508834 367066
rect 508890 367032 508924 367066
rect 508980 367032 509014 367066
rect 509070 367032 509104 367066
rect 509160 367032 509194 367066
rect 509250 367032 509284 367066
rect 509340 367032 509374 367066
rect 508800 366942 508834 366976
rect 508890 366942 508924 366976
rect 508980 366942 509014 366976
rect 509070 366942 509104 366976
rect 509160 366942 509194 366976
rect 509250 366942 509284 366976
rect 509340 366942 509374 366976
rect 508800 366852 508834 366886
rect 508890 366852 508924 366886
rect 508980 366852 509014 366886
rect 509070 366852 509104 366886
rect 509160 366852 509194 366886
rect 509250 366852 509284 366886
rect 509340 366852 509374 366886
rect 508800 366052 508834 366086
rect 508890 366052 508924 366086
rect 508980 366052 509014 366086
rect 509070 366052 509104 366086
rect 509160 366052 509194 366086
rect 509250 366052 509284 366086
rect 509340 366052 509374 366086
rect 508800 365962 508834 365996
rect 508890 365962 508924 365996
rect 508980 365962 509014 365996
rect 509070 365962 509104 365996
rect 509160 365962 509194 365996
rect 509250 365962 509284 365996
rect 509340 365962 509374 365996
rect 508800 365872 508834 365906
rect 508890 365872 508924 365906
rect 508980 365872 509014 365906
rect 509070 365872 509104 365906
rect 509160 365872 509194 365906
rect 509250 365872 509284 365906
rect 509340 365872 509374 365906
rect 508800 365782 508834 365816
rect 508890 365782 508924 365816
rect 508980 365782 509014 365816
rect 509070 365782 509104 365816
rect 509160 365782 509194 365816
rect 509250 365782 509284 365816
rect 509340 365782 509374 365816
rect 508800 365692 508834 365726
rect 508890 365692 508924 365726
rect 508980 365692 509014 365726
rect 509070 365692 509104 365726
rect 509160 365692 509194 365726
rect 509250 365692 509284 365726
rect 509340 365692 509374 365726
rect 508800 365602 508834 365636
rect 508890 365602 508924 365636
rect 508980 365602 509014 365636
rect 509070 365602 509104 365636
rect 509160 365602 509194 365636
rect 509250 365602 509284 365636
rect 509340 365602 509374 365636
rect 508800 365512 508834 365546
rect 508890 365512 508924 365546
rect 508980 365512 509014 365546
rect 509070 365512 509104 365546
rect 509160 365512 509194 365546
rect 509250 365512 509284 365546
rect 509340 365512 509374 365546
rect 508800 364712 508834 364746
rect 508890 364712 508924 364746
rect 508980 364712 509014 364746
rect 509070 364712 509104 364746
rect 509160 364712 509194 364746
rect 509250 364712 509284 364746
rect 509340 364712 509374 364746
rect 508800 364622 508834 364656
rect 508890 364622 508924 364656
rect 508980 364622 509014 364656
rect 509070 364622 509104 364656
rect 509160 364622 509194 364656
rect 509250 364622 509284 364656
rect 509340 364622 509374 364656
rect 508800 364532 508834 364566
rect 508890 364532 508924 364566
rect 508980 364532 509014 364566
rect 509070 364532 509104 364566
rect 509160 364532 509194 364566
rect 509250 364532 509284 364566
rect 509340 364532 509374 364566
rect 508800 364442 508834 364476
rect 508890 364442 508924 364476
rect 508980 364442 509014 364476
rect 509070 364442 509104 364476
rect 509160 364442 509194 364476
rect 509250 364442 509284 364476
rect 509340 364442 509374 364476
rect 508800 364352 508834 364386
rect 508890 364352 508924 364386
rect 508980 364352 509014 364386
rect 509070 364352 509104 364386
rect 509160 364352 509194 364386
rect 509250 364352 509284 364386
rect 509340 364352 509374 364386
rect 508800 364262 508834 364296
rect 508890 364262 508924 364296
rect 508980 364262 509014 364296
rect 509070 364262 509104 364296
rect 509160 364262 509194 364296
rect 509250 364262 509284 364296
rect 509340 364262 509374 364296
rect 508800 364172 508834 364206
rect 508890 364172 508924 364206
rect 508980 364172 509014 364206
rect 509070 364172 509104 364206
rect 509160 364172 509194 364206
rect 509250 364172 509284 364206
rect 509340 364172 509374 364206
rect 508800 363372 508834 363406
rect 508890 363372 508924 363406
rect 508980 363372 509014 363406
rect 509070 363372 509104 363406
rect 509160 363372 509194 363406
rect 509250 363372 509284 363406
rect 509340 363372 509374 363406
rect 508800 363282 508834 363316
rect 508890 363282 508924 363316
rect 508980 363282 509014 363316
rect 509070 363282 509104 363316
rect 509160 363282 509194 363316
rect 509250 363282 509284 363316
rect 509340 363282 509374 363316
rect 508800 363192 508834 363226
rect 508890 363192 508924 363226
rect 508980 363192 509014 363226
rect 509070 363192 509104 363226
rect 509160 363192 509194 363226
rect 509250 363192 509284 363226
rect 509340 363192 509374 363226
rect 508800 363102 508834 363136
rect 508890 363102 508924 363136
rect 508980 363102 509014 363136
rect 509070 363102 509104 363136
rect 509160 363102 509194 363136
rect 509250 363102 509284 363136
rect 509340 363102 509374 363136
rect 508800 363012 508834 363046
rect 508890 363012 508924 363046
rect 508980 363012 509014 363046
rect 509070 363012 509104 363046
rect 509160 363012 509194 363046
rect 509250 363012 509284 363046
rect 509340 363012 509374 363046
rect 508800 362922 508834 362956
rect 508890 362922 508924 362956
rect 508980 362922 509014 362956
rect 509070 362922 509104 362956
rect 509160 362922 509194 362956
rect 509250 362922 509284 362956
rect 509340 362922 509374 362956
rect 508800 362832 508834 362866
rect 508890 362832 508924 362866
rect 508980 362832 509014 362866
rect 509070 362832 509104 362866
rect 509160 362832 509194 362866
rect 509250 362832 509284 362866
rect 509340 362832 509374 362866
rect 512560 372752 512594 372786
rect 512650 372752 512684 372786
rect 512740 372752 512774 372786
rect 512830 372752 512864 372786
rect 512920 372752 512954 372786
rect 513010 372752 513044 372786
rect 513100 372752 513134 372786
rect 512560 372662 512594 372696
rect 512650 372662 512684 372696
rect 512740 372662 512774 372696
rect 512830 372662 512864 372696
rect 512920 372662 512954 372696
rect 513010 372662 513044 372696
rect 513100 372662 513134 372696
rect 512560 372572 512594 372606
rect 512650 372572 512684 372606
rect 512740 372572 512774 372606
rect 512830 372572 512864 372606
rect 512920 372572 512954 372606
rect 513010 372572 513044 372606
rect 513100 372572 513134 372606
rect 512560 372482 512594 372516
rect 512650 372482 512684 372516
rect 512740 372482 512774 372516
rect 512830 372482 512864 372516
rect 512920 372482 512954 372516
rect 513010 372482 513044 372516
rect 513100 372482 513134 372516
rect 512560 372392 512594 372426
rect 512650 372392 512684 372426
rect 512740 372392 512774 372426
rect 512830 372392 512864 372426
rect 512920 372392 512954 372426
rect 513010 372392 513044 372426
rect 513100 372392 513134 372426
rect 512560 372302 512594 372336
rect 512650 372302 512684 372336
rect 512740 372302 512774 372336
rect 512830 372302 512864 372336
rect 512920 372302 512954 372336
rect 513010 372302 513044 372336
rect 513100 372302 513134 372336
rect 512560 372212 512594 372246
rect 512650 372212 512684 372246
rect 512740 372212 512774 372246
rect 512830 372212 512864 372246
rect 512920 372212 512954 372246
rect 513010 372212 513044 372246
rect 513100 372212 513134 372246
rect 523439 374471 523473 374505
rect 523507 374471 523541 374505
rect 523575 374471 523609 374505
rect 523643 374471 523677 374505
rect 523711 374471 523745 374505
rect 523779 374471 523813 374505
rect 523847 374471 523881 374505
rect 523915 374471 523949 374505
rect 523983 374471 524017 374505
rect 524051 374471 524085 374505
rect 524119 374471 524153 374505
rect 524187 374471 524221 374505
rect 524255 374471 524289 374505
rect 524323 374471 524357 374505
rect 524391 374471 524425 374505
rect 524459 374471 524493 374505
rect 524527 374471 524561 374505
rect 524595 374471 524629 374505
rect 524663 374471 524697 374505
rect 523439 374013 523473 374047
rect 523507 374013 523541 374047
rect 523575 374013 523609 374047
rect 523643 374013 523677 374047
rect 523711 374013 523745 374047
rect 523779 374013 523813 374047
rect 523847 374013 523881 374047
rect 523915 374013 523949 374047
rect 523983 374013 524017 374047
rect 524051 374013 524085 374047
rect 524119 374013 524153 374047
rect 524187 374013 524221 374047
rect 524255 374013 524289 374047
rect 524323 374013 524357 374047
rect 524391 374013 524425 374047
rect 524459 374013 524493 374047
rect 524527 374013 524561 374047
rect 524595 374013 524629 374047
rect 524663 374013 524697 374047
rect 523439 373555 523473 373589
rect 523507 373555 523541 373589
rect 523575 373555 523609 373589
rect 523643 373555 523677 373589
rect 523711 373555 523745 373589
rect 523779 373555 523813 373589
rect 523847 373555 523881 373589
rect 523915 373555 523949 373589
rect 523983 373555 524017 373589
rect 524051 373555 524085 373589
rect 524119 373555 524153 373589
rect 524187 373555 524221 373589
rect 524255 373555 524289 373589
rect 524323 373555 524357 373589
rect 524391 373555 524425 373589
rect 524459 373555 524493 373589
rect 524527 373555 524561 373589
rect 524595 373555 524629 373589
rect 524663 373555 524697 373589
rect 523439 373097 523473 373131
rect 523507 373097 523541 373131
rect 523575 373097 523609 373131
rect 523643 373097 523677 373131
rect 523711 373097 523745 373131
rect 523779 373097 523813 373131
rect 523847 373097 523881 373131
rect 523915 373097 523949 373131
rect 523983 373097 524017 373131
rect 524051 373097 524085 373131
rect 524119 373097 524153 373131
rect 524187 373097 524221 373131
rect 524255 373097 524289 373131
rect 524323 373097 524357 373131
rect 524391 373097 524425 373131
rect 524459 373097 524493 373131
rect 524527 373097 524561 373131
rect 524595 373097 524629 373131
rect 524663 373097 524697 373131
rect 523439 372639 523473 372673
rect 523507 372639 523541 372673
rect 523575 372639 523609 372673
rect 523643 372639 523677 372673
rect 523711 372639 523745 372673
rect 523779 372639 523813 372673
rect 523847 372639 523881 372673
rect 523915 372639 523949 372673
rect 523983 372639 524017 372673
rect 524051 372639 524085 372673
rect 524119 372639 524153 372673
rect 524187 372639 524221 372673
rect 524255 372639 524289 372673
rect 524323 372639 524357 372673
rect 524391 372639 524425 372673
rect 524459 372639 524493 372673
rect 524527 372639 524561 372673
rect 524595 372639 524629 372673
rect 524663 372639 524697 372673
rect 523439 372181 523473 372215
rect 523507 372181 523541 372215
rect 523575 372181 523609 372215
rect 523643 372181 523677 372215
rect 523711 372181 523745 372215
rect 523779 372181 523813 372215
rect 523847 372181 523881 372215
rect 523915 372181 523949 372215
rect 523983 372181 524017 372215
rect 524051 372181 524085 372215
rect 524119 372181 524153 372215
rect 524187 372181 524221 372215
rect 524255 372181 524289 372215
rect 524323 372181 524357 372215
rect 524391 372181 524425 372215
rect 524459 372181 524493 372215
rect 524527 372181 524561 372215
rect 524595 372181 524629 372215
rect 524663 372181 524697 372215
rect 512560 371412 512594 371446
rect 512650 371412 512684 371446
rect 512740 371412 512774 371446
rect 512830 371412 512864 371446
rect 512920 371412 512954 371446
rect 513010 371412 513044 371446
rect 513100 371412 513134 371446
rect 512560 371322 512594 371356
rect 512650 371322 512684 371356
rect 512740 371322 512774 371356
rect 512830 371322 512864 371356
rect 512920 371322 512954 371356
rect 513010 371322 513044 371356
rect 513100 371322 513134 371356
rect 512560 371232 512594 371266
rect 512650 371232 512684 371266
rect 512740 371232 512774 371266
rect 512830 371232 512864 371266
rect 512920 371232 512954 371266
rect 513010 371232 513044 371266
rect 513100 371232 513134 371266
rect 512560 371142 512594 371176
rect 512650 371142 512684 371176
rect 512740 371142 512774 371176
rect 512830 371142 512864 371176
rect 512920 371142 512954 371176
rect 513010 371142 513044 371176
rect 513100 371142 513134 371176
rect 512560 371052 512594 371086
rect 512650 371052 512684 371086
rect 512740 371052 512774 371086
rect 512830 371052 512864 371086
rect 512920 371052 512954 371086
rect 513010 371052 513044 371086
rect 513100 371052 513134 371086
rect 512560 370962 512594 370996
rect 512650 370962 512684 370996
rect 512740 370962 512774 370996
rect 512830 370962 512864 370996
rect 512920 370962 512954 370996
rect 513010 370962 513044 370996
rect 513100 370962 513134 370996
rect 512560 370872 512594 370906
rect 512650 370872 512684 370906
rect 512740 370872 512774 370906
rect 512830 370872 512864 370906
rect 512920 370872 512954 370906
rect 513010 370872 513044 370906
rect 513100 370872 513134 370906
rect 512560 370072 512594 370106
rect 512650 370072 512684 370106
rect 512740 370072 512774 370106
rect 512830 370072 512864 370106
rect 512920 370072 512954 370106
rect 513010 370072 513044 370106
rect 513100 370072 513134 370106
rect 512560 369982 512594 370016
rect 512650 369982 512684 370016
rect 512740 369982 512774 370016
rect 512830 369982 512864 370016
rect 512920 369982 512954 370016
rect 513010 369982 513044 370016
rect 513100 369982 513134 370016
rect 512560 369892 512594 369926
rect 512650 369892 512684 369926
rect 512740 369892 512774 369926
rect 512830 369892 512864 369926
rect 512920 369892 512954 369926
rect 513010 369892 513044 369926
rect 513100 369892 513134 369926
rect 512560 369802 512594 369836
rect 512650 369802 512684 369836
rect 512740 369802 512774 369836
rect 512830 369802 512864 369836
rect 512920 369802 512954 369836
rect 513010 369802 513044 369836
rect 513100 369802 513134 369836
rect 512560 369712 512594 369746
rect 512650 369712 512684 369746
rect 512740 369712 512774 369746
rect 512830 369712 512864 369746
rect 512920 369712 512954 369746
rect 513010 369712 513044 369746
rect 513100 369712 513134 369746
rect 512560 369622 512594 369656
rect 512650 369622 512684 369656
rect 512740 369622 512774 369656
rect 512830 369622 512864 369656
rect 512920 369622 512954 369656
rect 513010 369622 513044 369656
rect 513100 369622 513134 369656
rect 512560 369532 512594 369566
rect 512650 369532 512684 369566
rect 512740 369532 512774 369566
rect 512830 369532 512864 369566
rect 512920 369532 512954 369566
rect 513010 369532 513044 369566
rect 513100 369532 513134 369566
rect 523439 371723 523473 371757
rect 523507 371723 523541 371757
rect 523575 371723 523609 371757
rect 523643 371723 523677 371757
rect 523711 371723 523745 371757
rect 523779 371723 523813 371757
rect 523847 371723 523881 371757
rect 523915 371723 523949 371757
rect 523983 371723 524017 371757
rect 524051 371723 524085 371757
rect 524119 371723 524153 371757
rect 524187 371723 524221 371757
rect 524255 371723 524289 371757
rect 524323 371723 524357 371757
rect 524391 371723 524425 371757
rect 524459 371723 524493 371757
rect 524527 371723 524561 371757
rect 524595 371723 524629 371757
rect 524663 371723 524697 371757
rect 523439 371265 523473 371299
rect 523507 371265 523541 371299
rect 523575 371265 523609 371299
rect 523643 371265 523677 371299
rect 523711 371265 523745 371299
rect 523779 371265 523813 371299
rect 523847 371265 523881 371299
rect 523915 371265 523949 371299
rect 523983 371265 524017 371299
rect 524051 371265 524085 371299
rect 524119 371265 524153 371299
rect 524187 371265 524221 371299
rect 524255 371265 524289 371299
rect 524323 371265 524357 371299
rect 524391 371265 524425 371299
rect 524459 371265 524493 371299
rect 524527 371265 524561 371299
rect 524595 371265 524629 371299
rect 524663 371265 524697 371299
rect 523439 370807 523473 370841
rect 523507 370807 523541 370841
rect 523575 370807 523609 370841
rect 523643 370807 523677 370841
rect 523711 370807 523745 370841
rect 523779 370807 523813 370841
rect 523847 370807 523881 370841
rect 523915 370807 523949 370841
rect 523983 370807 524017 370841
rect 524051 370807 524085 370841
rect 524119 370807 524153 370841
rect 524187 370807 524221 370841
rect 524255 370807 524289 370841
rect 524323 370807 524357 370841
rect 524391 370807 524425 370841
rect 524459 370807 524493 370841
rect 524527 370807 524561 370841
rect 524595 370807 524629 370841
rect 524663 370807 524697 370841
rect 523439 370349 523473 370383
rect 523507 370349 523541 370383
rect 523575 370349 523609 370383
rect 523643 370349 523677 370383
rect 523711 370349 523745 370383
rect 523779 370349 523813 370383
rect 523847 370349 523881 370383
rect 523915 370349 523949 370383
rect 523983 370349 524017 370383
rect 524051 370349 524085 370383
rect 524119 370349 524153 370383
rect 524187 370349 524221 370383
rect 524255 370349 524289 370383
rect 524323 370349 524357 370383
rect 524391 370349 524425 370383
rect 524459 370349 524493 370383
rect 524527 370349 524561 370383
rect 524595 370349 524629 370383
rect 524663 370349 524697 370383
rect 523439 369891 523473 369925
rect 523507 369891 523541 369925
rect 523575 369891 523609 369925
rect 523643 369891 523677 369925
rect 523711 369891 523745 369925
rect 523779 369891 523813 369925
rect 523847 369891 523881 369925
rect 523915 369891 523949 369925
rect 523983 369891 524017 369925
rect 524051 369891 524085 369925
rect 524119 369891 524153 369925
rect 524187 369891 524221 369925
rect 524255 369891 524289 369925
rect 524323 369891 524357 369925
rect 524391 369891 524425 369925
rect 524459 369891 524493 369925
rect 524527 369891 524561 369925
rect 524595 369891 524629 369925
rect 524663 369891 524697 369925
rect 523439 369433 523473 369467
rect 523507 369433 523541 369467
rect 523575 369433 523609 369467
rect 523643 369433 523677 369467
rect 523711 369433 523745 369467
rect 523779 369433 523813 369467
rect 523847 369433 523881 369467
rect 523915 369433 523949 369467
rect 523983 369433 524017 369467
rect 524051 369433 524085 369467
rect 524119 369433 524153 369467
rect 524187 369433 524221 369467
rect 524255 369433 524289 369467
rect 524323 369433 524357 369467
rect 524391 369433 524425 369467
rect 524459 369433 524493 369467
rect 524527 369433 524561 369467
rect 524595 369433 524629 369467
rect 524663 369433 524697 369467
rect 512560 368732 512594 368766
rect 512650 368732 512684 368766
rect 512740 368732 512774 368766
rect 512830 368732 512864 368766
rect 512920 368732 512954 368766
rect 513010 368732 513044 368766
rect 513100 368732 513134 368766
rect 512560 368642 512594 368676
rect 512650 368642 512684 368676
rect 512740 368642 512774 368676
rect 512830 368642 512864 368676
rect 512920 368642 512954 368676
rect 513010 368642 513044 368676
rect 513100 368642 513134 368676
rect 512560 368552 512594 368586
rect 512650 368552 512684 368586
rect 512740 368552 512774 368586
rect 512830 368552 512864 368586
rect 512920 368552 512954 368586
rect 513010 368552 513044 368586
rect 513100 368552 513134 368586
rect 512560 368462 512594 368496
rect 512650 368462 512684 368496
rect 512740 368462 512774 368496
rect 512830 368462 512864 368496
rect 512920 368462 512954 368496
rect 513010 368462 513044 368496
rect 513100 368462 513134 368496
rect 512560 368372 512594 368406
rect 512650 368372 512684 368406
rect 512740 368372 512774 368406
rect 512830 368372 512864 368406
rect 512920 368372 512954 368406
rect 513010 368372 513044 368406
rect 513100 368372 513134 368406
rect 512560 368282 512594 368316
rect 512650 368282 512684 368316
rect 512740 368282 512774 368316
rect 512830 368282 512864 368316
rect 512920 368282 512954 368316
rect 513010 368282 513044 368316
rect 513100 368282 513134 368316
rect 512560 368192 512594 368226
rect 512650 368192 512684 368226
rect 512740 368192 512774 368226
rect 512830 368192 512864 368226
rect 512920 368192 512954 368226
rect 513010 368192 513044 368226
rect 513100 368192 513134 368226
rect 512560 367392 512594 367426
rect 512650 367392 512684 367426
rect 512740 367392 512774 367426
rect 512830 367392 512864 367426
rect 512920 367392 512954 367426
rect 513010 367392 513044 367426
rect 513100 367392 513134 367426
rect 512560 367302 512594 367336
rect 512650 367302 512684 367336
rect 512740 367302 512774 367336
rect 512830 367302 512864 367336
rect 512920 367302 512954 367336
rect 513010 367302 513044 367336
rect 513100 367302 513134 367336
rect 512560 367212 512594 367246
rect 512650 367212 512684 367246
rect 512740 367212 512774 367246
rect 512830 367212 512864 367246
rect 512920 367212 512954 367246
rect 513010 367212 513044 367246
rect 513100 367212 513134 367246
rect 512560 367122 512594 367156
rect 512650 367122 512684 367156
rect 512740 367122 512774 367156
rect 512830 367122 512864 367156
rect 512920 367122 512954 367156
rect 513010 367122 513044 367156
rect 513100 367122 513134 367156
rect 512560 367032 512594 367066
rect 512650 367032 512684 367066
rect 512740 367032 512774 367066
rect 512830 367032 512864 367066
rect 512920 367032 512954 367066
rect 513010 367032 513044 367066
rect 513100 367032 513134 367066
rect 512560 366942 512594 366976
rect 512650 366942 512684 366976
rect 512740 366942 512774 366976
rect 512830 366942 512864 366976
rect 512920 366942 512954 366976
rect 513010 366942 513044 366976
rect 513100 366942 513134 366976
rect 512560 366852 512594 366886
rect 512650 366852 512684 366886
rect 512740 366852 512774 366886
rect 512830 366852 512864 366886
rect 512920 366852 512954 366886
rect 513010 366852 513044 366886
rect 513100 366852 513134 366886
rect 523439 368975 523473 369009
rect 523507 368975 523541 369009
rect 523575 368975 523609 369009
rect 523643 368975 523677 369009
rect 523711 368975 523745 369009
rect 523779 368975 523813 369009
rect 523847 368975 523881 369009
rect 523915 368975 523949 369009
rect 523983 368975 524017 369009
rect 524051 368975 524085 369009
rect 524119 368975 524153 369009
rect 524187 368975 524221 369009
rect 524255 368975 524289 369009
rect 524323 368975 524357 369009
rect 524391 368975 524425 369009
rect 524459 368975 524493 369009
rect 524527 368975 524561 369009
rect 524595 368975 524629 369009
rect 524663 368975 524697 369009
rect 523439 368517 523473 368551
rect 523507 368517 523541 368551
rect 523575 368517 523609 368551
rect 523643 368517 523677 368551
rect 523711 368517 523745 368551
rect 523779 368517 523813 368551
rect 523847 368517 523881 368551
rect 523915 368517 523949 368551
rect 523983 368517 524017 368551
rect 524051 368517 524085 368551
rect 524119 368517 524153 368551
rect 524187 368517 524221 368551
rect 524255 368517 524289 368551
rect 524323 368517 524357 368551
rect 524391 368517 524425 368551
rect 524459 368517 524493 368551
rect 524527 368517 524561 368551
rect 524595 368517 524629 368551
rect 524663 368517 524697 368551
rect 523439 368059 523473 368093
rect 523507 368059 523541 368093
rect 523575 368059 523609 368093
rect 523643 368059 523677 368093
rect 523711 368059 523745 368093
rect 523779 368059 523813 368093
rect 523847 368059 523881 368093
rect 523915 368059 523949 368093
rect 523983 368059 524017 368093
rect 524051 368059 524085 368093
rect 524119 368059 524153 368093
rect 524187 368059 524221 368093
rect 524255 368059 524289 368093
rect 524323 368059 524357 368093
rect 524391 368059 524425 368093
rect 524459 368059 524493 368093
rect 524527 368059 524561 368093
rect 524595 368059 524629 368093
rect 524663 368059 524697 368093
rect 523439 367601 523473 367635
rect 523507 367601 523541 367635
rect 523575 367601 523609 367635
rect 523643 367601 523677 367635
rect 523711 367601 523745 367635
rect 523779 367601 523813 367635
rect 523847 367601 523881 367635
rect 523915 367601 523949 367635
rect 523983 367601 524017 367635
rect 524051 367601 524085 367635
rect 524119 367601 524153 367635
rect 524187 367601 524221 367635
rect 524255 367601 524289 367635
rect 524323 367601 524357 367635
rect 524391 367601 524425 367635
rect 524459 367601 524493 367635
rect 524527 367601 524561 367635
rect 524595 367601 524629 367635
rect 524663 367601 524697 367635
rect 523439 367143 523473 367177
rect 523507 367143 523541 367177
rect 523575 367143 523609 367177
rect 523643 367143 523677 367177
rect 523711 367143 523745 367177
rect 523779 367143 523813 367177
rect 523847 367143 523881 367177
rect 523915 367143 523949 367177
rect 523983 367143 524017 367177
rect 524051 367143 524085 367177
rect 524119 367143 524153 367177
rect 524187 367143 524221 367177
rect 524255 367143 524289 367177
rect 524323 367143 524357 367177
rect 524391 367143 524425 367177
rect 524459 367143 524493 367177
rect 524527 367143 524561 367177
rect 524595 367143 524629 367177
rect 524663 367143 524697 367177
rect 523439 366685 523473 366719
rect 523507 366685 523541 366719
rect 523575 366685 523609 366719
rect 523643 366685 523677 366719
rect 523711 366685 523745 366719
rect 523779 366685 523813 366719
rect 523847 366685 523881 366719
rect 523915 366685 523949 366719
rect 523983 366685 524017 366719
rect 524051 366685 524085 366719
rect 524119 366685 524153 366719
rect 524187 366685 524221 366719
rect 524255 366685 524289 366719
rect 524323 366685 524357 366719
rect 524391 366685 524425 366719
rect 524459 366685 524493 366719
rect 524527 366685 524561 366719
rect 524595 366685 524629 366719
rect 524663 366685 524697 366719
rect 512560 366052 512594 366086
rect 512650 366052 512684 366086
rect 512740 366052 512774 366086
rect 512830 366052 512864 366086
rect 512920 366052 512954 366086
rect 513010 366052 513044 366086
rect 513100 366052 513134 366086
rect 512560 365962 512594 365996
rect 512650 365962 512684 365996
rect 512740 365962 512774 365996
rect 512830 365962 512864 365996
rect 512920 365962 512954 365996
rect 513010 365962 513044 365996
rect 513100 365962 513134 365996
rect 512560 365872 512594 365906
rect 512650 365872 512684 365906
rect 512740 365872 512774 365906
rect 512830 365872 512864 365906
rect 512920 365872 512954 365906
rect 513010 365872 513044 365906
rect 513100 365872 513134 365906
rect 512560 365782 512594 365816
rect 512650 365782 512684 365816
rect 512740 365782 512774 365816
rect 512830 365782 512864 365816
rect 512920 365782 512954 365816
rect 513010 365782 513044 365816
rect 513100 365782 513134 365816
rect 512560 365692 512594 365726
rect 512650 365692 512684 365726
rect 512740 365692 512774 365726
rect 512830 365692 512864 365726
rect 512920 365692 512954 365726
rect 513010 365692 513044 365726
rect 513100 365692 513134 365726
rect 512560 365602 512594 365636
rect 512650 365602 512684 365636
rect 512740 365602 512774 365636
rect 512830 365602 512864 365636
rect 512920 365602 512954 365636
rect 513010 365602 513044 365636
rect 513100 365602 513134 365636
rect 512560 365512 512594 365546
rect 512650 365512 512684 365546
rect 512740 365512 512774 365546
rect 512830 365512 512864 365546
rect 512920 365512 512954 365546
rect 513010 365512 513044 365546
rect 513100 365512 513134 365546
rect 512560 364712 512594 364746
rect 512650 364712 512684 364746
rect 512740 364712 512774 364746
rect 512830 364712 512864 364746
rect 512920 364712 512954 364746
rect 513010 364712 513044 364746
rect 513100 364712 513134 364746
rect 512560 364622 512594 364656
rect 512650 364622 512684 364656
rect 512740 364622 512774 364656
rect 512830 364622 512864 364656
rect 512920 364622 512954 364656
rect 513010 364622 513044 364656
rect 513100 364622 513134 364656
rect 512560 364532 512594 364566
rect 512650 364532 512684 364566
rect 512740 364532 512774 364566
rect 512830 364532 512864 364566
rect 512920 364532 512954 364566
rect 513010 364532 513044 364566
rect 513100 364532 513134 364566
rect 512560 364442 512594 364476
rect 512650 364442 512684 364476
rect 512740 364442 512774 364476
rect 512830 364442 512864 364476
rect 512920 364442 512954 364476
rect 513010 364442 513044 364476
rect 513100 364442 513134 364476
rect 512560 364352 512594 364386
rect 512650 364352 512684 364386
rect 512740 364352 512774 364386
rect 512830 364352 512864 364386
rect 512920 364352 512954 364386
rect 513010 364352 513044 364386
rect 513100 364352 513134 364386
rect 512560 364262 512594 364296
rect 512650 364262 512684 364296
rect 512740 364262 512774 364296
rect 512830 364262 512864 364296
rect 512920 364262 512954 364296
rect 513010 364262 513044 364296
rect 513100 364262 513134 364296
rect 512560 364172 512594 364206
rect 512650 364172 512684 364206
rect 512740 364172 512774 364206
rect 512830 364172 512864 364206
rect 512920 364172 512954 364206
rect 513010 364172 513044 364206
rect 513100 364172 513134 364206
rect 523439 366227 523473 366261
rect 523507 366227 523541 366261
rect 523575 366227 523609 366261
rect 523643 366227 523677 366261
rect 523711 366227 523745 366261
rect 523779 366227 523813 366261
rect 523847 366227 523881 366261
rect 523915 366227 523949 366261
rect 523983 366227 524017 366261
rect 524051 366227 524085 366261
rect 524119 366227 524153 366261
rect 524187 366227 524221 366261
rect 524255 366227 524289 366261
rect 524323 366227 524357 366261
rect 524391 366227 524425 366261
rect 524459 366227 524493 366261
rect 524527 366227 524561 366261
rect 524595 366227 524629 366261
rect 524663 366227 524697 366261
rect 523439 365769 523473 365803
rect 523507 365769 523541 365803
rect 523575 365769 523609 365803
rect 523643 365769 523677 365803
rect 523711 365769 523745 365803
rect 523779 365769 523813 365803
rect 523847 365769 523881 365803
rect 523915 365769 523949 365803
rect 523983 365769 524017 365803
rect 524051 365769 524085 365803
rect 524119 365769 524153 365803
rect 524187 365769 524221 365803
rect 524255 365769 524289 365803
rect 524323 365769 524357 365803
rect 524391 365769 524425 365803
rect 524459 365769 524493 365803
rect 524527 365769 524561 365803
rect 524595 365769 524629 365803
rect 524663 365769 524697 365803
rect 523439 365311 523473 365345
rect 523507 365311 523541 365345
rect 523575 365311 523609 365345
rect 523643 365311 523677 365345
rect 523711 365311 523745 365345
rect 523779 365311 523813 365345
rect 523847 365311 523881 365345
rect 523915 365311 523949 365345
rect 523983 365311 524017 365345
rect 524051 365311 524085 365345
rect 524119 365311 524153 365345
rect 524187 365311 524221 365345
rect 524255 365311 524289 365345
rect 524323 365311 524357 365345
rect 524391 365311 524425 365345
rect 524459 365311 524493 365345
rect 524527 365311 524561 365345
rect 524595 365311 524629 365345
rect 524663 365311 524697 365345
rect 523439 364853 523473 364887
rect 523507 364853 523541 364887
rect 523575 364853 523609 364887
rect 523643 364853 523677 364887
rect 523711 364853 523745 364887
rect 523779 364853 523813 364887
rect 523847 364853 523881 364887
rect 523915 364853 523949 364887
rect 523983 364853 524017 364887
rect 524051 364853 524085 364887
rect 524119 364853 524153 364887
rect 524187 364853 524221 364887
rect 524255 364853 524289 364887
rect 524323 364853 524357 364887
rect 524391 364853 524425 364887
rect 524459 364853 524493 364887
rect 524527 364853 524561 364887
rect 524595 364853 524629 364887
rect 524663 364853 524697 364887
rect 523439 364395 523473 364429
rect 523507 364395 523541 364429
rect 523575 364395 523609 364429
rect 523643 364395 523677 364429
rect 523711 364395 523745 364429
rect 523779 364395 523813 364429
rect 523847 364395 523881 364429
rect 523915 364395 523949 364429
rect 523983 364395 524017 364429
rect 524051 364395 524085 364429
rect 524119 364395 524153 364429
rect 524187 364395 524221 364429
rect 524255 364395 524289 364429
rect 524323 364395 524357 364429
rect 524391 364395 524425 364429
rect 524459 364395 524493 364429
rect 524527 364395 524561 364429
rect 524595 364395 524629 364429
rect 524663 364395 524697 364429
rect 523439 363937 523473 363971
rect 523507 363937 523541 363971
rect 523575 363937 523609 363971
rect 523643 363937 523677 363971
rect 523711 363937 523745 363971
rect 523779 363937 523813 363971
rect 523847 363937 523881 363971
rect 523915 363937 523949 363971
rect 523983 363937 524017 363971
rect 524051 363937 524085 363971
rect 524119 363937 524153 363971
rect 524187 363937 524221 363971
rect 524255 363937 524289 363971
rect 524323 363937 524357 363971
rect 524391 363937 524425 363971
rect 524459 363937 524493 363971
rect 524527 363937 524561 363971
rect 524595 363937 524629 363971
rect 524663 363937 524697 363971
rect 512560 363372 512594 363406
rect 512650 363372 512684 363406
rect 512740 363372 512774 363406
rect 512830 363372 512864 363406
rect 512920 363372 512954 363406
rect 513010 363372 513044 363406
rect 513100 363372 513134 363406
rect 512560 363282 512594 363316
rect 512650 363282 512684 363316
rect 512740 363282 512774 363316
rect 512830 363282 512864 363316
rect 512920 363282 512954 363316
rect 513010 363282 513044 363316
rect 513100 363282 513134 363316
rect 512560 363192 512594 363226
rect 512650 363192 512684 363226
rect 512740 363192 512774 363226
rect 512830 363192 512864 363226
rect 512920 363192 512954 363226
rect 513010 363192 513044 363226
rect 513100 363192 513134 363226
rect 512560 363102 512594 363136
rect 512650 363102 512684 363136
rect 512740 363102 512774 363136
rect 512830 363102 512864 363136
rect 512920 363102 512954 363136
rect 513010 363102 513044 363136
rect 513100 363102 513134 363136
rect 512560 363012 512594 363046
rect 512650 363012 512684 363046
rect 512740 363012 512774 363046
rect 512830 363012 512864 363046
rect 512920 363012 512954 363046
rect 513010 363012 513044 363046
rect 513100 363012 513134 363046
rect 512560 362922 512594 362956
rect 512650 362922 512684 362956
rect 512740 362922 512774 362956
rect 512830 362922 512864 362956
rect 512920 362922 512954 362956
rect 513010 362922 513044 362956
rect 513100 362922 513134 362956
rect 512560 362832 512594 362866
rect 512650 362832 512684 362866
rect 512740 362832 512774 362866
rect 512830 362832 512864 362866
rect 512920 362832 512954 362866
rect 513010 362832 513044 362866
rect 513100 362832 513134 362866
rect 523439 363479 523473 363513
rect 523507 363479 523541 363513
rect 523575 363479 523609 363513
rect 523643 363479 523677 363513
rect 523711 363479 523745 363513
rect 523779 363479 523813 363513
rect 523847 363479 523881 363513
rect 523915 363479 523949 363513
rect 523983 363479 524017 363513
rect 524051 363479 524085 363513
rect 524119 363479 524153 363513
rect 524187 363479 524221 363513
rect 524255 363479 524289 363513
rect 524323 363479 524357 363513
rect 524391 363479 524425 363513
rect 524459 363479 524493 363513
rect 524527 363479 524561 363513
rect 524595 363479 524629 363513
rect 524663 363479 524697 363513
rect 523439 363021 523473 363055
rect 523507 363021 523541 363055
rect 523575 363021 523609 363055
rect 523643 363021 523677 363055
rect 523711 363021 523745 363055
rect 523779 363021 523813 363055
rect 523847 363021 523881 363055
rect 523915 363021 523949 363055
rect 523983 363021 524017 363055
rect 524051 363021 524085 363055
rect 524119 363021 524153 363055
rect 524187 363021 524221 363055
rect 524255 363021 524289 363055
rect 524323 363021 524357 363055
rect 524391 363021 524425 363055
rect 524459 363021 524493 363055
rect 524527 363021 524561 363055
rect 524595 363021 524629 363055
rect 524663 363021 524697 363055
rect 523439 362563 523473 362597
rect 523507 362563 523541 362597
rect 523575 362563 523609 362597
rect 523643 362563 523677 362597
rect 523711 362563 523745 362597
rect 523779 362563 523813 362597
rect 523847 362563 523881 362597
rect 523915 362563 523949 362597
rect 523983 362563 524017 362597
rect 524051 362563 524085 362597
rect 524119 362563 524153 362597
rect 524187 362563 524221 362597
rect 524255 362563 524289 362597
rect 524323 362563 524357 362597
rect 524391 362563 524425 362597
rect 524459 362563 524493 362597
rect 524527 362563 524561 362597
rect 524595 362563 524629 362597
rect 524663 362563 524697 362597
rect 574691 357922 574725 358898
rect 574949 357922 574983 358898
rect 575207 357922 575241 358898
rect 575465 357922 575499 358898
rect 575723 357922 575757 358898
rect 575981 357922 576015 358898
rect 576239 357922 576273 358898
rect 576497 357922 576531 358898
rect 576755 357922 576789 358898
rect 577013 357922 577047 358898
rect 577271 357922 577305 358898
rect 577529 357922 577563 358898
rect 577787 357922 577821 358898
rect 578045 357922 578079 358898
rect 578303 357922 578337 358898
rect 578561 357922 578595 358898
rect 578819 357922 578853 358898
rect 579077 357922 579111 358898
rect 579335 357922 579369 358898
rect 579593 357922 579627 358898
rect 579851 357922 579885 358898
rect 575139 311754 575173 312730
rect 575397 311754 575431 312730
rect 575655 311754 575689 312730
rect 575913 311754 575947 312730
rect 576171 311754 576205 312730
rect 576429 311754 576463 312730
rect 576687 311754 576721 312730
rect 576945 311754 576979 312730
rect 577203 311754 577237 312730
rect 577461 311754 577495 312730
rect 577719 311754 577753 312730
rect 577977 311754 578011 312730
rect 578235 311754 578269 312730
rect 578493 311754 578527 312730
rect 578751 311754 578785 312730
rect 579009 311754 579043 312730
rect 579267 311754 579301 312730
rect 579525 311754 579559 312730
rect 579783 311754 579817 312730
rect 580041 311754 580075 312730
rect 580299 311754 580333 312730
<< psubdiff >>
rect 565886 492100 565926 492140
rect 562148 492068 562268 492070
rect 562148 492032 562184 492068
rect 562228 492032 562268 492068
rect 562148 492020 562268 492032
rect 563448 492068 563568 492070
rect 563448 492032 563484 492068
rect 563528 492032 563568 492068
rect 563448 492020 563568 492032
rect 564748 492068 564868 492070
rect 564748 492032 564784 492068
rect 564828 492032 564868 492068
rect 564748 492020 564868 492032
rect 565886 492020 565926 492060
rect 560630 402958 560670 402998
rect 504684 402902 505972 402936
rect 504684 402868 504742 402902
rect 504776 402868 504832 402902
rect 504866 402868 504922 402902
rect 504956 402868 505012 402902
rect 505046 402868 505102 402902
rect 505136 402868 505192 402902
rect 505226 402868 505282 402902
rect 505316 402868 505372 402902
rect 505406 402868 505462 402902
rect 505496 402868 505552 402902
rect 505586 402868 505642 402902
rect 505676 402868 505732 402902
rect 505766 402868 505822 402902
rect 505856 402868 505972 402902
rect 560630 402878 560670 402918
rect 561688 402926 561808 402928
rect 561688 402890 561728 402926
rect 561772 402890 561808 402926
rect 561688 402878 561808 402890
rect 562988 402926 563108 402928
rect 562988 402890 563028 402926
rect 563072 402890 563108 402926
rect 562988 402878 563108 402890
rect 564288 402926 564408 402928
rect 564288 402890 564328 402926
rect 564372 402890 564408 402926
rect 564288 402878 564408 402890
rect 504684 402835 505972 402868
rect 504684 402806 504785 402835
rect 504684 402772 504719 402806
rect 504753 402772 504785 402806
rect 505871 402806 505972 402835
rect 504684 402716 504785 402772
rect 504684 402682 504719 402716
rect 504753 402682 504785 402716
rect 504684 402626 504785 402682
rect 504684 402592 504719 402626
rect 504753 402592 504785 402626
rect 504684 402536 504785 402592
rect 504684 402502 504719 402536
rect 504753 402502 504785 402536
rect 504684 402446 504785 402502
rect 504684 402412 504719 402446
rect 504753 402412 504785 402446
rect 504684 402356 504785 402412
rect 504684 402322 504719 402356
rect 504753 402322 504785 402356
rect 504684 402266 504785 402322
rect 504684 402232 504719 402266
rect 504753 402232 504785 402266
rect 504684 402176 504785 402232
rect 504684 402142 504719 402176
rect 504753 402142 504785 402176
rect 504684 402086 504785 402142
rect 504684 402052 504719 402086
rect 504753 402052 504785 402086
rect 504684 401996 504785 402052
rect 504684 401962 504719 401996
rect 504753 401962 504785 401996
rect 504684 401906 504785 401962
rect 504684 401872 504719 401906
rect 504753 401872 504785 401906
rect 504684 401816 504785 401872
rect 504684 401782 504719 401816
rect 504753 401782 504785 401816
rect 505871 402772 505906 402806
rect 505940 402772 505972 402806
rect 505871 402716 505972 402772
rect 505871 402682 505906 402716
rect 505940 402682 505972 402716
rect 505871 402626 505972 402682
rect 505871 402592 505906 402626
rect 505940 402592 505972 402626
rect 505871 402536 505972 402592
rect 505871 402502 505906 402536
rect 505940 402502 505972 402536
rect 505871 402446 505972 402502
rect 505871 402412 505906 402446
rect 505940 402412 505972 402446
rect 505871 402356 505972 402412
rect 505871 402322 505906 402356
rect 505940 402322 505972 402356
rect 505871 402266 505972 402322
rect 505871 402232 505906 402266
rect 505940 402232 505972 402266
rect 505871 402176 505972 402232
rect 505871 402142 505906 402176
rect 505940 402142 505972 402176
rect 505871 402086 505972 402142
rect 505871 402052 505906 402086
rect 505940 402052 505972 402086
rect 505871 401996 505972 402052
rect 505871 401962 505906 401996
rect 505940 401962 505972 401996
rect 505871 401906 505972 401962
rect 505871 401872 505906 401906
rect 505940 401872 505972 401906
rect 505871 401816 505972 401872
rect 504684 401749 504785 401782
rect 505871 401782 505906 401816
rect 505940 401782 505972 401816
rect 505871 401749 505972 401782
rect 504684 401715 505972 401749
rect 504684 401681 504742 401715
rect 504776 401681 504832 401715
rect 504866 401681 504922 401715
rect 504956 401681 505012 401715
rect 505046 401681 505102 401715
rect 505136 401681 505192 401715
rect 505226 401681 505282 401715
rect 505316 401681 505372 401715
rect 505406 401681 505462 401715
rect 505496 401681 505552 401715
rect 505586 401681 505642 401715
rect 505676 401681 505732 401715
rect 505766 401681 505822 401715
rect 505856 401681 505972 401715
rect 504684 401648 505972 401681
rect 498548 400893 498668 400896
rect 498548 400859 498591 400893
rect 498625 400859 498668 400893
rect 498548 400856 498668 400859
rect 505298 400277 505478 400364
rect 505298 399835 505337 400277
rect 505439 399835 505478 400277
rect 505298 399748 505478 399835
rect 505298 397533 505478 397620
rect 505298 397091 505337 397533
rect 505439 397091 505478 397533
rect 505298 397004 505478 397091
rect 512818 397435 512998 397522
rect 512818 396993 512857 397435
rect 512959 396993 512998 397435
rect 512818 396906 512998 396993
rect 494018 393123 494198 393210
rect 494018 392681 494057 393123
rect 494159 392681 494198 393123
rect 494018 392594 494198 392681
rect 505298 394501 505478 394588
rect 505298 394059 505337 394501
rect 505439 394059 505478 394501
rect 505298 393972 505478 394059
rect 509058 394691 509238 394778
rect 509058 394249 509097 394691
rect 509199 394249 509238 394691
rect 509058 394162 509238 394249
rect 512818 394691 512998 394778
rect 512818 394249 512857 394691
rect 512959 394249 512998 394691
rect 512818 394162 512998 394249
rect 494788 391093 494908 391096
rect 494788 391059 494831 391093
rect 494865 391059 494908 391093
rect 494788 391056 494908 391059
rect 505298 391457 505478 391544
rect 505298 391015 505337 391457
rect 505439 391015 505478 391457
rect 505298 390928 505478 391015
rect 509058 391659 509238 391746
rect 509058 391217 509097 391659
rect 509199 391217 509238 391659
rect 509058 391130 509238 391217
rect 512818 391947 512998 392034
rect 512818 391505 512857 391947
rect 512959 391505 512998 391947
rect 512818 391418 512998 391505
rect 516578 391555 516758 391642
rect 516578 391113 516617 391555
rect 516719 391113 516758 391555
rect 516578 391026 516758 391113
rect 506068 389593 506188 389596
rect 506068 389559 506111 389593
rect 506145 389559 506188 389593
rect 506068 389556 506188 389559
rect 517348 389593 517468 389596
rect 517348 389559 517391 389593
rect 517425 389559 517468 389593
rect 517348 389556 517468 389559
rect 506138 388491 506188 388536
rect 506138 388457 506141 388491
rect 506175 388457 506188 388491
rect 506138 388416 506188 388457
rect 520338 390085 520518 390172
rect 520338 389643 520377 390085
rect 520479 389643 520518 390085
rect 520338 389556 520518 389643
rect 517418 388491 517468 388536
rect 517418 388457 517421 388491
rect 517455 388457 517468 388491
rect 517418 388416 517468 388457
rect 506138 387191 506188 387236
rect 506138 387157 506141 387191
rect 506175 387157 506188 387191
rect 506138 387116 506188 387157
rect 512818 386753 512998 386840
rect 512818 386311 512857 386753
rect 512959 386311 512998 386753
rect 512818 386224 512998 386311
rect 517418 387191 517468 387236
rect 517418 387157 517421 387191
rect 517455 387157 517468 387191
rect 517418 387116 517468 387157
rect 520338 386753 520518 386840
rect 520338 386311 520377 386753
rect 520479 386311 520518 386753
rect 520338 386224 520518 386311
rect 520338 384009 520518 384096
rect 520338 383567 520377 384009
rect 520479 383567 520518 384009
rect 520338 383480 520518 383567
rect 520338 380775 520518 380862
rect 520338 380333 520377 380775
rect 520479 380333 520518 380775
rect 520338 380246 520518 380333
rect 502308 377735 502428 377738
rect 502308 377701 502351 377735
rect 502385 377701 502428 377735
rect 502308 377698 502428 377701
rect 502378 376633 502428 376678
rect 502378 376599 502381 376633
rect 502415 376599 502428 376633
rect 502378 376558 502428 376599
rect 502378 375333 502428 375378
rect 502378 375299 502381 375333
rect 502415 375299 502428 375333
rect 502378 375258 502428 375299
rect 516578 376561 516758 376648
rect 516578 376119 516617 376561
rect 516719 376119 516758 376561
rect 516578 376032 516758 376119
rect 520338 376561 520518 376648
rect 520338 376119 520377 376561
rect 520479 376119 520518 376561
rect 520338 376032 520518 376119
rect 500924 373110 502212 373144
rect 500924 373076 500982 373110
rect 501016 373076 501072 373110
rect 501106 373076 501162 373110
rect 501196 373076 501252 373110
rect 501286 373076 501342 373110
rect 501376 373076 501432 373110
rect 501466 373076 501522 373110
rect 501556 373076 501612 373110
rect 501646 373076 501702 373110
rect 501736 373076 501792 373110
rect 501826 373076 501882 373110
rect 501916 373076 501972 373110
rect 502006 373076 502062 373110
rect 502096 373076 502212 373110
rect 500924 373043 502212 373076
rect 500924 373014 501025 373043
rect 500924 372980 500959 373014
rect 500993 372980 501025 373014
rect 502111 373014 502212 373043
rect 500924 372924 501025 372980
rect 500924 372890 500959 372924
rect 500993 372890 501025 372924
rect 500924 372834 501025 372890
rect 500924 372800 500959 372834
rect 500993 372800 501025 372834
rect 500924 372744 501025 372800
rect 500924 372710 500959 372744
rect 500993 372710 501025 372744
rect 500924 372654 501025 372710
rect 500924 372620 500959 372654
rect 500993 372620 501025 372654
rect 500924 372564 501025 372620
rect 500924 372530 500959 372564
rect 500993 372530 501025 372564
rect 500924 372474 501025 372530
rect 500924 372440 500959 372474
rect 500993 372440 501025 372474
rect 500924 372384 501025 372440
rect 500924 372350 500959 372384
rect 500993 372350 501025 372384
rect 500924 372294 501025 372350
rect 500924 372260 500959 372294
rect 500993 372260 501025 372294
rect 500924 372204 501025 372260
rect 500924 372170 500959 372204
rect 500993 372170 501025 372204
rect 500924 372114 501025 372170
rect 500924 372080 500959 372114
rect 500993 372080 501025 372114
rect 500924 372024 501025 372080
rect 500924 371990 500959 372024
rect 500993 371990 501025 372024
rect 502111 372980 502146 373014
rect 502180 372980 502212 373014
rect 502111 372924 502212 372980
rect 502111 372890 502146 372924
rect 502180 372890 502212 372924
rect 502111 372834 502212 372890
rect 502111 372800 502146 372834
rect 502180 372800 502212 372834
rect 502111 372744 502212 372800
rect 502111 372710 502146 372744
rect 502180 372710 502212 372744
rect 502111 372654 502212 372710
rect 502111 372620 502146 372654
rect 502180 372620 502212 372654
rect 502111 372564 502212 372620
rect 502111 372530 502146 372564
rect 502180 372530 502212 372564
rect 502111 372474 502212 372530
rect 502111 372440 502146 372474
rect 502180 372440 502212 372474
rect 502111 372384 502212 372440
rect 502111 372350 502146 372384
rect 502180 372350 502212 372384
rect 502111 372294 502212 372350
rect 502111 372260 502146 372294
rect 502180 372260 502212 372294
rect 502111 372204 502212 372260
rect 502111 372170 502146 372204
rect 502180 372170 502212 372204
rect 502111 372114 502212 372170
rect 502111 372080 502146 372114
rect 502180 372080 502212 372114
rect 502111 372024 502212 372080
rect 497164 371934 498452 371968
rect 497164 371900 497222 371934
rect 497256 371900 497312 371934
rect 497346 371900 497402 371934
rect 497436 371900 497492 371934
rect 497526 371900 497582 371934
rect 497616 371900 497672 371934
rect 497706 371900 497762 371934
rect 497796 371900 497852 371934
rect 497886 371900 497942 371934
rect 497976 371900 498032 371934
rect 498066 371900 498122 371934
rect 498156 371900 498212 371934
rect 498246 371900 498302 371934
rect 498336 371900 498452 371934
rect 497164 371867 498452 371900
rect 497164 371838 497265 371867
rect 497164 371804 497199 371838
rect 497233 371804 497265 371838
rect 498351 371838 498452 371867
rect 497164 371748 497265 371804
rect 497164 371714 497199 371748
rect 497233 371714 497265 371748
rect 497164 371658 497265 371714
rect 497164 371624 497199 371658
rect 497233 371624 497265 371658
rect 497164 371568 497265 371624
rect 497164 371534 497199 371568
rect 497233 371534 497265 371568
rect 497164 371478 497265 371534
rect 497164 371444 497199 371478
rect 497233 371444 497265 371478
rect 497164 371388 497265 371444
rect 497164 371354 497199 371388
rect 497233 371354 497265 371388
rect 497164 371298 497265 371354
rect 497164 371264 497199 371298
rect 497233 371264 497265 371298
rect 497164 371208 497265 371264
rect 497164 371174 497199 371208
rect 497233 371174 497265 371208
rect 497164 371118 497265 371174
rect 497164 371084 497199 371118
rect 497233 371084 497265 371118
rect 497164 371028 497265 371084
rect 497164 370994 497199 371028
rect 497233 370994 497265 371028
rect 497164 370938 497265 370994
rect 497164 370904 497199 370938
rect 497233 370904 497265 370938
rect 497164 370848 497265 370904
rect 497164 370814 497199 370848
rect 497233 370814 497265 370848
rect 498351 371804 498386 371838
rect 498420 371804 498452 371838
rect 498351 371748 498452 371804
rect 498351 371714 498386 371748
rect 498420 371714 498452 371748
rect 498351 371658 498452 371714
rect 498351 371624 498386 371658
rect 498420 371624 498452 371658
rect 498351 371568 498452 371624
rect 498351 371534 498386 371568
rect 498420 371534 498452 371568
rect 498351 371478 498452 371534
rect 498351 371444 498386 371478
rect 498420 371444 498452 371478
rect 498351 371388 498452 371444
rect 498351 371354 498386 371388
rect 498420 371354 498452 371388
rect 498351 371298 498452 371354
rect 498351 371264 498386 371298
rect 498420 371264 498452 371298
rect 498351 371208 498452 371264
rect 498351 371174 498386 371208
rect 498420 371174 498452 371208
rect 498351 371118 498452 371174
rect 498351 371084 498386 371118
rect 498420 371084 498452 371118
rect 498351 371028 498452 371084
rect 498351 370994 498386 371028
rect 498420 370994 498452 371028
rect 498351 370938 498452 370994
rect 498351 370904 498386 370938
rect 498420 370904 498452 370938
rect 498351 370848 498452 370904
rect 497164 370781 497265 370814
rect 498351 370814 498386 370848
rect 498420 370814 498452 370848
rect 498351 370781 498452 370814
rect 497164 370747 498452 370781
rect 497164 370713 497222 370747
rect 497256 370713 497312 370747
rect 497346 370713 497402 370747
rect 497436 370713 497492 370747
rect 497526 370713 497582 370747
rect 497616 370713 497672 370747
rect 497706 370713 497762 370747
rect 497796 370713 497852 370747
rect 497886 370713 497942 370747
rect 497976 370713 498032 370747
rect 498066 370713 498122 370747
rect 498156 370713 498212 370747
rect 498246 370713 498302 370747
rect 498336 370713 498452 370747
rect 497164 370594 498452 370713
rect 497164 370560 497222 370594
rect 497256 370560 497312 370594
rect 497346 370560 497402 370594
rect 497436 370560 497492 370594
rect 497526 370560 497582 370594
rect 497616 370560 497672 370594
rect 497706 370560 497762 370594
rect 497796 370560 497852 370594
rect 497886 370560 497942 370594
rect 497976 370560 498032 370594
rect 498066 370560 498122 370594
rect 498156 370560 498212 370594
rect 498246 370560 498302 370594
rect 498336 370560 498452 370594
rect 497164 370527 498452 370560
rect 497164 370498 497265 370527
rect 497164 370464 497199 370498
rect 497233 370464 497265 370498
rect 498351 370498 498452 370527
rect 497164 370408 497265 370464
rect 497164 370374 497199 370408
rect 497233 370374 497265 370408
rect 497164 370318 497265 370374
rect 497164 370284 497199 370318
rect 497233 370284 497265 370318
rect 497164 370228 497265 370284
rect 497164 370194 497199 370228
rect 497233 370194 497265 370228
rect 497164 370138 497265 370194
rect 497164 370104 497199 370138
rect 497233 370104 497265 370138
rect 497164 370048 497265 370104
rect 497164 370014 497199 370048
rect 497233 370014 497265 370048
rect 497164 369958 497265 370014
rect 497164 369924 497199 369958
rect 497233 369924 497265 369958
rect 497164 369868 497265 369924
rect 497164 369834 497199 369868
rect 497233 369834 497265 369868
rect 497164 369778 497265 369834
rect 497164 369744 497199 369778
rect 497233 369744 497265 369778
rect 497164 369688 497265 369744
rect 497164 369654 497199 369688
rect 497233 369654 497265 369688
rect 497164 369598 497265 369654
rect 497164 369564 497199 369598
rect 497233 369564 497265 369598
rect 497164 369508 497265 369564
rect 497164 369474 497199 369508
rect 497233 369474 497265 369508
rect 498351 370464 498386 370498
rect 498420 370464 498452 370498
rect 498351 370408 498452 370464
rect 498351 370374 498386 370408
rect 498420 370374 498452 370408
rect 498351 370318 498452 370374
rect 498351 370284 498386 370318
rect 498420 370284 498452 370318
rect 498351 370228 498452 370284
rect 498351 370194 498386 370228
rect 498420 370194 498452 370228
rect 498351 370138 498452 370194
rect 498351 370104 498386 370138
rect 498420 370104 498452 370138
rect 498351 370048 498452 370104
rect 498351 370014 498386 370048
rect 498420 370014 498452 370048
rect 498351 369958 498452 370014
rect 498351 369924 498386 369958
rect 498420 369924 498452 369958
rect 498351 369868 498452 369924
rect 498351 369834 498386 369868
rect 498420 369834 498452 369868
rect 498351 369778 498452 369834
rect 498351 369744 498386 369778
rect 498420 369744 498452 369778
rect 498351 369688 498452 369744
rect 498351 369654 498386 369688
rect 498420 369654 498452 369688
rect 498351 369598 498452 369654
rect 498351 369564 498386 369598
rect 498420 369564 498452 369598
rect 498351 369508 498452 369564
rect 497164 369441 497265 369474
rect 498351 369474 498386 369508
rect 498420 369474 498452 369508
rect 498351 369441 498452 369474
rect 497164 369407 498452 369441
rect 497164 369373 497222 369407
rect 497256 369373 497312 369407
rect 497346 369373 497402 369407
rect 497436 369373 497492 369407
rect 497526 369373 497582 369407
rect 497616 369373 497672 369407
rect 497706 369373 497762 369407
rect 497796 369373 497852 369407
rect 497886 369373 497942 369407
rect 497976 369373 498032 369407
rect 498066 369373 498122 369407
rect 498156 369373 498212 369407
rect 498246 369373 498302 369407
rect 498336 369373 498452 369407
rect 497164 369254 498452 369373
rect 497164 369220 497222 369254
rect 497256 369220 497312 369254
rect 497346 369220 497402 369254
rect 497436 369220 497492 369254
rect 497526 369220 497582 369254
rect 497616 369220 497672 369254
rect 497706 369220 497762 369254
rect 497796 369220 497852 369254
rect 497886 369220 497942 369254
rect 497976 369220 498032 369254
rect 498066 369220 498122 369254
rect 498156 369220 498212 369254
rect 498246 369220 498302 369254
rect 498336 369220 498452 369254
rect 497164 369187 498452 369220
rect 497164 369158 497265 369187
rect 497164 369124 497199 369158
rect 497233 369124 497265 369158
rect 498351 369158 498452 369187
rect 497164 369068 497265 369124
rect 497164 369034 497199 369068
rect 497233 369034 497265 369068
rect 497164 368978 497265 369034
rect 497164 368944 497199 368978
rect 497233 368944 497265 368978
rect 497164 368888 497265 368944
rect 497164 368854 497199 368888
rect 497233 368854 497265 368888
rect 497164 368798 497265 368854
rect 497164 368764 497199 368798
rect 497233 368764 497265 368798
rect 497164 368708 497265 368764
rect 497164 368674 497199 368708
rect 497233 368674 497265 368708
rect 497164 368618 497265 368674
rect 497164 368584 497199 368618
rect 497233 368584 497265 368618
rect 497164 368528 497265 368584
rect 497164 368494 497199 368528
rect 497233 368494 497265 368528
rect 497164 368438 497265 368494
rect 497164 368404 497199 368438
rect 497233 368404 497265 368438
rect 497164 368348 497265 368404
rect 497164 368314 497199 368348
rect 497233 368314 497265 368348
rect 497164 368258 497265 368314
rect 497164 368224 497199 368258
rect 497233 368224 497265 368258
rect 497164 368168 497265 368224
rect 497164 368134 497199 368168
rect 497233 368134 497265 368168
rect 498351 369124 498386 369158
rect 498420 369124 498452 369158
rect 498351 369068 498452 369124
rect 498351 369034 498386 369068
rect 498420 369034 498452 369068
rect 498351 368978 498452 369034
rect 498351 368944 498386 368978
rect 498420 368944 498452 368978
rect 498351 368888 498452 368944
rect 498351 368854 498386 368888
rect 498420 368854 498452 368888
rect 498351 368798 498452 368854
rect 498351 368764 498386 368798
rect 498420 368764 498452 368798
rect 498351 368708 498452 368764
rect 498351 368674 498386 368708
rect 498420 368674 498452 368708
rect 498351 368618 498452 368674
rect 498351 368584 498386 368618
rect 498420 368584 498452 368618
rect 498351 368528 498452 368584
rect 498351 368494 498386 368528
rect 498420 368494 498452 368528
rect 498351 368438 498452 368494
rect 498351 368404 498386 368438
rect 498420 368404 498452 368438
rect 498351 368348 498452 368404
rect 498351 368314 498386 368348
rect 498420 368314 498452 368348
rect 498351 368258 498452 368314
rect 498351 368224 498386 368258
rect 498420 368224 498452 368258
rect 498351 368168 498452 368224
rect 497164 368101 497265 368134
rect 498351 368134 498386 368168
rect 498420 368134 498452 368168
rect 498351 368101 498452 368134
rect 497164 368067 498452 368101
rect 497164 368033 497222 368067
rect 497256 368033 497312 368067
rect 497346 368033 497402 368067
rect 497436 368033 497492 368067
rect 497526 368033 497582 368067
rect 497616 368033 497672 368067
rect 497706 368033 497762 368067
rect 497796 368033 497852 368067
rect 497886 368033 497942 368067
rect 497976 368033 498032 368067
rect 498066 368033 498122 368067
rect 498156 368033 498212 368067
rect 498246 368033 498302 368067
rect 498336 368033 498452 368067
rect 497164 367914 498452 368033
rect 497164 367880 497222 367914
rect 497256 367880 497312 367914
rect 497346 367880 497402 367914
rect 497436 367880 497492 367914
rect 497526 367880 497582 367914
rect 497616 367880 497672 367914
rect 497706 367880 497762 367914
rect 497796 367880 497852 367914
rect 497886 367880 497942 367914
rect 497976 367880 498032 367914
rect 498066 367880 498122 367914
rect 498156 367880 498212 367914
rect 498246 367880 498302 367914
rect 498336 367880 498452 367914
rect 497164 367847 498452 367880
rect 497164 367818 497265 367847
rect 497164 367784 497199 367818
rect 497233 367784 497265 367818
rect 498351 367818 498452 367847
rect 497164 367728 497265 367784
rect 497164 367694 497199 367728
rect 497233 367694 497265 367728
rect 497164 367638 497265 367694
rect 497164 367604 497199 367638
rect 497233 367604 497265 367638
rect 497164 367548 497265 367604
rect 497164 367514 497199 367548
rect 497233 367514 497265 367548
rect 497164 367458 497265 367514
rect 497164 367424 497199 367458
rect 497233 367424 497265 367458
rect 497164 367368 497265 367424
rect 497164 367334 497199 367368
rect 497233 367334 497265 367368
rect 497164 367278 497265 367334
rect 497164 367244 497199 367278
rect 497233 367244 497265 367278
rect 497164 367188 497265 367244
rect 497164 367154 497199 367188
rect 497233 367154 497265 367188
rect 497164 367098 497265 367154
rect 497164 367064 497199 367098
rect 497233 367064 497265 367098
rect 497164 367008 497265 367064
rect 497164 366974 497199 367008
rect 497233 366974 497265 367008
rect 497164 366918 497265 366974
rect 497164 366884 497199 366918
rect 497233 366884 497265 366918
rect 497164 366828 497265 366884
rect 497164 366794 497199 366828
rect 497233 366794 497265 366828
rect 498351 367784 498386 367818
rect 498420 367784 498452 367818
rect 498351 367728 498452 367784
rect 498351 367694 498386 367728
rect 498420 367694 498452 367728
rect 498351 367638 498452 367694
rect 498351 367604 498386 367638
rect 498420 367604 498452 367638
rect 498351 367548 498452 367604
rect 498351 367514 498386 367548
rect 498420 367514 498452 367548
rect 498351 367458 498452 367514
rect 498351 367424 498386 367458
rect 498420 367424 498452 367458
rect 498351 367368 498452 367424
rect 498351 367334 498386 367368
rect 498420 367334 498452 367368
rect 498351 367278 498452 367334
rect 498351 367244 498386 367278
rect 498420 367244 498452 367278
rect 498351 367188 498452 367244
rect 498351 367154 498386 367188
rect 498420 367154 498452 367188
rect 498351 367098 498452 367154
rect 498351 367064 498386 367098
rect 498420 367064 498452 367098
rect 498351 367008 498452 367064
rect 498351 366974 498386 367008
rect 498420 366974 498452 367008
rect 498351 366918 498452 366974
rect 498351 366884 498386 366918
rect 498420 366884 498452 366918
rect 498351 366828 498452 366884
rect 497164 366761 497265 366794
rect 498351 366794 498386 366828
rect 498420 366794 498452 366828
rect 498351 366761 498452 366794
rect 497164 366727 498452 366761
rect 497164 366693 497222 366727
rect 497256 366693 497312 366727
rect 497346 366693 497402 366727
rect 497436 366693 497492 366727
rect 497526 366693 497582 366727
rect 497616 366693 497672 366727
rect 497706 366693 497762 366727
rect 497796 366693 497852 366727
rect 497886 366693 497942 366727
rect 497976 366693 498032 366727
rect 498066 366693 498122 366727
rect 498156 366693 498212 366727
rect 498246 366693 498302 366727
rect 498336 366693 498452 366727
rect 497164 366574 498452 366693
rect 497164 366540 497222 366574
rect 497256 366540 497312 366574
rect 497346 366540 497402 366574
rect 497436 366540 497492 366574
rect 497526 366540 497582 366574
rect 497616 366540 497672 366574
rect 497706 366540 497762 366574
rect 497796 366540 497852 366574
rect 497886 366540 497942 366574
rect 497976 366540 498032 366574
rect 498066 366540 498122 366574
rect 498156 366540 498212 366574
rect 498246 366540 498302 366574
rect 498336 366540 498452 366574
rect 497164 366507 498452 366540
rect 497164 366478 497265 366507
rect 497164 366444 497199 366478
rect 497233 366444 497265 366478
rect 498351 366478 498452 366507
rect 497164 366388 497265 366444
rect 497164 366354 497199 366388
rect 497233 366354 497265 366388
rect 497164 366298 497265 366354
rect 497164 366264 497199 366298
rect 497233 366264 497265 366298
rect 497164 366208 497265 366264
rect 497164 366174 497199 366208
rect 497233 366174 497265 366208
rect 497164 366118 497265 366174
rect 497164 366084 497199 366118
rect 497233 366084 497265 366118
rect 497164 366028 497265 366084
rect 497164 365994 497199 366028
rect 497233 365994 497265 366028
rect 497164 365938 497265 365994
rect 497164 365904 497199 365938
rect 497233 365904 497265 365938
rect 497164 365848 497265 365904
rect 497164 365814 497199 365848
rect 497233 365814 497265 365848
rect 497164 365758 497265 365814
rect 497164 365724 497199 365758
rect 497233 365724 497265 365758
rect 497164 365668 497265 365724
rect 497164 365634 497199 365668
rect 497233 365634 497265 365668
rect 497164 365578 497265 365634
rect 497164 365544 497199 365578
rect 497233 365544 497265 365578
rect 497164 365488 497265 365544
rect 497164 365454 497199 365488
rect 497233 365454 497265 365488
rect 498351 366444 498386 366478
rect 498420 366444 498452 366478
rect 498351 366388 498452 366444
rect 498351 366354 498386 366388
rect 498420 366354 498452 366388
rect 498351 366298 498452 366354
rect 498351 366264 498386 366298
rect 498420 366264 498452 366298
rect 498351 366208 498452 366264
rect 498351 366174 498386 366208
rect 498420 366174 498452 366208
rect 498351 366118 498452 366174
rect 498351 366084 498386 366118
rect 498420 366084 498452 366118
rect 498351 366028 498452 366084
rect 498351 365994 498386 366028
rect 498420 365994 498452 366028
rect 498351 365938 498452 365994
rect 498351 365904 498386 365938
rect 498420 365904 498452 365938
rect 498351 365848 498452 365904
rect 498351 365814 498386 365848
rect 498420 365814 498452 365848
rect 498351 365758 498452 365814
rect 498351 365724 498386 365758
rect 498420 365724 498452 365758
rect 498351 365668 498452 365724
rect 498351 365634 498386 365668
rect 498420 365634 498452 365668
rect 498351 365578 498452 365634
rect 498351 365544 498386 365578
rect 498420 365544 498452 365578
rect 498351 365488 498452 365544
rect 497164 365421 497265 365454
rect 498351 365454 498386 365488
rect 498420 365454 498452 365488
rect 498351 365421 498452 365454
rect 497164 365387 498452 365421
rect 497164 365353 497222 365387
rect 497256 365353 497312 365387
rect 497346 365353 497402 365387
rect 497436 365353 497492 365387
rect 497526 365353 497582 365387
rect 497616 365353 497672 365387
rect 497706 365353 497762 365387
rect 497796 365353 497852 365387
rect 497886 365353 497942 365387
rect 497976 365353 498032 365387
rect 498066 365353 498122 365387
rect 498156 365353 498212 365387
rect 498246 365353 498302 365387
rect 498336 365353 498452 365387
rect 497164 365234 498452 365353
rect 497164 365200 497222 365234
rect 497256 365200 497312 365234
rect 497346 365200 497402 365234
rect 497436 365200 497492 365234
rect 497526 365200 497582 365234
rect 497616 365200 497672 365234
rect 497706 365200 497762 365234
rect 497796 365200 497852 365234
rect 497886 365200 497942 365234
rect 497976 365200 498032 365234
rect 498066 365200 498122 365234
rect 498156 365200 498212 365234
rect 498246 365200 498302 365234
rect 498336 365200 498452 365234
rect 497164 365167 498452 365200
rect 497164 365138 497265 365167
rect 497164 365104 497199 365138
rect 497233 365104 497265 365138
rect 498351 365138 498452 365167
rect 497164 365048 497265 365104
rect 497164 365014 497199 365048
rect 497233 365014 497265 365048
rect 497164 364958 497265 365014
rect 497164 364924 497199 364958
rect 497233 364924 497265 364958
rect 497164 364868 497265 364924
rect 497164 364834 497199 364868
rect 497233 364834 497265 364868
rect 497164 364778 497265 364834
rect 497164 364744 497199 364778
rect 497233 364744 497265 364778
rect 497164 364688 497265 364744
rect 497164 364654 497199 364688
rect 497233 364654 497265 364688
rect 497164 364598 497265 364654
rect 497164 364564 497199 364598
rect 497233 364564 497265 364598
rect 497164 364508 497265 364564
rect 497164 364474 497199 364508
rect 497233 364474 497265 364508
rect 497164 364418 497265 364474
rect 497164 364384 497199 364418
rect 497233 364384 497265 364418
rect 497164 364328 497265 364384
rect 497164 364294 497199 364328
rect 497233 364294 497265 364328
rect 497164 364238 497265 364294
rect 497164 364204 497199 364238
rect 497233 364204 497265 364238
rect 497164 364148 497265 364204
rect 497164 364114 497199 364148
rect 497233 364114 497265 364148
rect 498351 365104 498386 365138
rect 498420 365104 498452 365138
rect 498351 365048 498452 365104
rect 498351 365014 498386 365048
rect 498420 365014 498452 365048
rect 498351 364958 498452 365014
rect 498351 364924 498386 364958
rect 498420 364924 498452 364958
rect 498351 364868 498452 364924
rect 498351 364834 498386 364868
rect 498420 364834 498452 364868
rect 498351 364778 498452 364834
rect 498351 364744 498386 364778
rect 498420 364744 498452 364778
rect 498351 364688 498452 364744
rect 498351 364654 498386 364688
rect 498420 364654 498452 364688
rect 498351 364598 498452 364654
rect 498351 364564 498386 364598
rect 498420 364564 498452 364598
rect 498351 364508 498452 364564
rect 498351 364474 498386 364508
rect 498420 364474 498452 364508
rect 498351 364418 498452 364474
rect 498351 364384 498386 364418
rect 498420 364384 498452 364418
rect 498351 364328 498452 364384
rect 498351 364294 498386 364328
rect 498420 364294 498452 364328
rect 498351 364238 498452 364294
rect 498351 364204 498386 364238
rect 498420 364204 498452 364238
rect 498351 364148 498452 364204
rect 497164 364081 497265 364114
rect 498351 364114 498386 364148
rect 498420 364114 498452 364148
rect 498351 364081 498452 364114
rect 497164 364047 498452 364081
rect 497164 364013 497222 364047
rect 497256 364013 497312 364047
rect 497346 364013 497402 364047
rect 497436 364013 497492 364047
rect 497526 364013 497582 364047
rect 497616 364013 497672 364047
rect 497706 364013 497762 364047
rect 497796 364013 497852 364047
rect 497886 364013 497942 364047
rect 497976 364013 498032 364047
rect 498066 364013 498122 364047
rect 498156 364013 498212 364047
rect 498246 364013 498302 364047
rect 498336 364013 498452 364047
rect 497164 363894 498452 364013
rect 497164 363860 497222 363894
rect 497256 363860 497312 363894
rect 497346 363860 497402 363894
rect 497436 363860 497492 363894
rect 497526 363860 497582 363894
rect 497616 363860 497672 363894
rect 497706 363860 497762 363894
rect 497796 363860 497852 363894
rect 497886 363860 497942 363894
rect 497976 363860 498032 363894
rect 498066 363860 498122 363894
rect 498156 363860 498212 363894
rect 498246 363860 498302 363894
rect 498336 363860 498452 363894
rect 497164 363827 498452 363860
rect 497164 363798 497265 363827
rect 497164 363764 497199 363798
rect 497233 363764 497265 363798
rect 498351 363798 498452 363827
rect 497164 363708 497265 363764
rect 497164 363674 497199 363708
rect 497233 363674 497265 363708
rect 497164 363618 497265 363674
rect 497164 363584 497199 363618
rect 497233 363584 497265 363618
rect 497164 363528 497265 363584
rect 497164 363494 497199 363528
rect 497233 363494 497265 363528
rect 497164 363438 497265 363494
rect 497164 363404 497199 363438
rect 497233 363404 497265 363438
rect 497164 363348 497265 363404
rect 497164 363314 497199 363348
rect 497233 363314 497265 363348
rect 497164 363258 497265 363314
rect 497164 363224 497199 363258
rect 497233 363224 497265 363258
rect 497164 363168 497265 363224
rect 497164 363134 497199 363168
rect 497233 363134 497265 363168
rect 497164 363078 497265 363134
rect 497164 363044 497199 363078
rect 497233 363044 497265 363078
rect 497164 362988 497265 363044
rect 497164 362954 497199 362988
rect 497233 362954 497265 362988
rect 497164 362898 497265 362954
rect 497164 362864 497199 362898
rect 497233 362864 497265 362898
rect 497164 362808 497265 362864
rect 497164 362774 497199 362808
rect 497233 362774 497265 362808
rect 498351 363764 498386 363798
rect 498420 363764 498452 363798
rect 498351 363708 498452 363764
rect 498351 363674 498386 363708
rect 498420 363674 498452 363708
rect 498351 363618 498452 363674
rect 498351 363584 498386 363618
rect 498420 363584 498452 363618
rect 498351 363528 498452 363584
rect 498351 363494 498386 363528
rect 498420 363494 498452 363528
rect 498351 363438 498452 363494
rect 498351 363404 498386 363438
rect 498420 363404 498452 363438
rect 498351 363348 498452 363404
rect 498351 363314 498386 363348
rect 498420 363314 498452 363348
rect 498351 363258 498452 363314
rect 498351 363224 498386 363258
rect 498420 363224 498452 363258
rect 498351 363168 498452 363224
rect 498351 363134 498386 363168
rect 498420 363134 498452 363168
rect 498351 363078 498452 363134
rect 498351 363044 498386 363078
rect 498420 363044 498452 363078
rect 498351 362988 498452 363044
rect 498351 362954 498386 362988
rect 498420 362954 498452 362988
rect 498351 362898 498452 362954
rect 498351 362864 498386 362898
rect 498420 362864 498452 362898
rect 498351 362808 498452 362864
rect 497164 362741 497265 362774
rect 498351 362774 498386 362808
rect 498420 362774 498452 362808
rect 498351 362741 498452 362774
rect 497164 362707 498452 362741
rect 497164 362673 497222 362707
rect 497256 362673 497312 362707
rect 497346 362673 497402 362707
rect 497436 362673 497492 362707
rect 497526 362673 497582 362707
rect 497616 362673 497672 362707
rect 497706 362673 497762 362707
rect 497796 362673 497852 362707
rect 497886 362673 497942 362707
rect 497976 362673 498032 362707
rect 498066 362673 498122 362707
rect 498156 362673 498212 362707
rect 498246 362673 498302 362707
rect 498336 362673 498452 362707
rect 497164 362640 498452 362673
rect 500924 371957 501025 371990
rect 502111 371990 502146 372024
rect 502180 371990 502212 372024
rect 502111 371957 502212 371990
rect 500924 371923 502212 371957
rect 500924 371889 500982 371923
rect 501016 371889 501072 371923
rect 501106 371889 501162 371923
rect 501196 371889 501252 371923
rect 501286 371889 501342 371923
rect 501376 371889 501432 371923
rect 501466 371889 501522 371923
rect 501556 371889 501612 371923
rect 501646 371889 501702 371923
rect 501736 371889 501792 371923
rect 501826 371889 501882 371923
rect 501916 371889 501972 371923
rect 502006 371889 502062 371923
rect 502096 371889 502212 371923
rect 500924 371770 502212 371889
rect 500924 371736 500982 371770
rect 501016 371736 501072 371770
rect 501106 371736 501162 371770
rect 501196 371736 501252 371770
rect 501286 371736 501342 371770
rect 501376 371736 501432 371770
rect 501466 371736 501522 371770
rect 501556 371736 501612 371770
rect 501646 371736 501702 371770
rect 501736 371736 501792 371770
rect 501826 371736 501882 371770
rect 501916 371736 501972 371770
rect 502006 371736 502062 371770
rect 502096 371736 502212 371770
rect 500924 371703 502212 371736
rect 500924 371674 501025 371703
rect 500924 371640 500959 371674
rect 500993 371640 501025 371674
rect 502111 371674 502212 371703
rect 500924 371584 501025 371640
rect 500924 371550 500959 371584
rect 500993 371550 501025 371584
rect 500924 371494 501025 371550
rect 500924 371460 500959 371494
rect 500993 371460 501025 371494
rect 500924 371404 501025 371460
rect 500924 371370 500959 371404
rect 500993 371370 501025 371404
rect 500924 371314 501025 371370
rect 500924 371280 500959 371314
rect 500993 371280 501025 371314
rect 500924 371224 501025 371280
rect 500924 371190 500959 371224
rect 500993 371190 501025 371224
rect 500924 371134 501025 371190
rect 500924 371100 500959 371134
rect 500993 371100 501025 371134
rect 500924 371044 501025 371100
rect 500924 371010 500959 371044
rect 500993 371010 501025 371044
rect 500924 370954 501025 371010
rect 500924 370920 500959 370954
rect 500993 370920 501025 370954
rect 500924 370864 501025 370920
rect 500924 370830 500959 370864
rect 500993 370830 501025 370864
rect 500924 370774 501025 370830
rect 500924 370740 500959 370774
rect 500993 370740 501025 370774
rect 500924 370684 501025 370740
rect 500924 370650 500959 370684
rect 500993 370650 501025 370684
rect 502111 371640 502146 371674
rect 502180 371640 502212 371674
rect 502111 371584 502212 371640
rect 502111 371550 502146 371584
rect 502180 371550 502212 371584
rect 502111 371494 502212 371550
rect 502111 371460 502146 371494
rect 502180 371460 502212 371494
rect 502111 371404 502212 371460
rect 502111 371370 502146 371404
rect 502180 371370 502212 371404
rect 502111 371314 502212 371370
rect 502111 371280 502146 371314
rect 502180 371280 502212 371314
rect 502111 371224 502212 371280
rect 502111 371190 502146 371224
rect 502180 371190 502212 371224
rect 502111 371134 502212 371190
rect 502111 371100 502146 371134
rect 502180 371100 502212 371134
rect 502111 371044 502212 371100
rect 502111 371010 502146 371044
rect 502180 371010 502212 371044
rect 502111 370954 502212 371010
rect 502111 370920 502146 370954
rect 502180 370920 502212 370954
rect 502111 370864 502212 370920
rect 502111 370830 502146 370864
rect 502180 370830 502212 370864
rect 502111 370774 502212 370830
rect 502111 370740 502146 370774
rect 502180 370740 502212 370774
rect 502111 370684 502212 370740
rect 500924 370617 501025 370650
rect 502111 370650 502146 370684
rect 502180 370650 502212 370684
rect 502111 370617 502212 370650
rect 500924 370583 502212 370617
rect 500924 370549 500982 370583
rect 501016 370549 501072 370583
rect 501106 370549 501162 370583
rect 501196 370549 501252 370583
rect 501286 370549 501342 370583
rect 501376 370549 501432 370583
rect 501466 370549 501522 370583
rect 501556 370549 501612 370583
rect 501646 370549 501702 370583
rect 501736 370549 501792 370583
rect 501826 370549 501882 370583
rect 501916 370549 501972 370583
rect 502006 370549 502062 370583
rect 502096 370549 502212 370583
rect 500924 370430 502212 370549
rect 500924 370396 500982 370430
rect 501016 370396 501072 370430
rect 501106 370396 501162 370430
rect 501196 370396 501252 370430
rect 501286 370396 501342 370430
rect 501376 370396 501432 370430
rect 501466 370396 501522 370430
rect 501556 370396 501612 370430
rect 501646 370396 501702 370430
rect 501736 370396 501792 370430
rect 501826 370396 501882 370430
rect 501916 370396 501972 370430
rect 502006 370396 502062 370430
rect 502096 370396 502212 370430
rect 500924 370363 502212 370396
rect 500924 370334 501025 370363
rect 500924 370300 500959 370334
rect 500993 370300 501025 370334
rect 502111 370334 502212 370363
rect 500924 370244 501025 370300
rect 500924 370210 500959 370244
rect 500993 370210 501025 370244
rect 500924 370154 501025 370210
rect 500924 370120 500959 370154
rect 500993 370120 501025 370154
rect 500924 370064 501025 370120
rect 500924 370030 500959 370064
rect 500993 370030 501025 370064
rect 500924 369974 501025 370030
rect 500924 369940 500959 369974
rect 500993 369940 501025 369974
rect 500924 369884 501025 369940
rect 500924 369850 500959 369884
rect 500993 369850 501025 369884
rect 500924 369794 501025 369850
rect 500924 369760 500959 369794
rect 500993 369760 501025 369794
rect 500924 369704 501025 369760
rect 500924 369670 500959 369704
rect 500993 369670 501025 369704
rect 500924 369614 501025 369670
rect 500924 369580 500959 369614
rect 500993 369580 501025 369614
rect 500924 369524 501025 369580
rect 500924 369490 500959 369524
rect 500993 369490 501025 369524
rect 500924 369434 501025 369490
rect 500924 369400 500959 369434
rect 500993 369400 501025 369434
rect 500924 369344 501025 369400
rect 500924 369310 500959 369344
rect 500993 369310 501025 369344
rect 502111 370300 502146 370334
rect 502180 370300 502212 370334
rect 502111 370244 502212 370300
rect 502111 370210 502146 370244
rect 502180 370210 502212 370244
rect 502111 370154 502212 370210
rect 502111 370120 502146 370154
rect 502180 370120 502212 370154
rect 502111 370064 502212 370120
rect 502111 370030 502146 370064
rect 502180 370030 502212 370064
rect 502111 369974 502212 370030
rect 502111 369940 502146 369974
rect 502180 369940 502212 369974
rect 502111 369884 502212 369940
rect 502111 369850 502146 369884
rect 502180 369850 502212 369884
rect 502111 369794 502212 369850
rect 502111 369760 502146 369794
rect 502180 369760 502212 369794
rect 502111 369704 502212 369760
rect 502111 369670 502146 369704
rect 502180 369670 502212 369704
rect 502111 369614 502212 369670
rect 502111 369580 502146 369614
rect 502180 369580 502212 369614
rect 502111 369524 502212 369580
rect 502111 369490 502146 369524
rect 502180 369490 502212 369524
rect 502111 369434 502212 369490
rect 502111 369400 502146 369434
rect 502180 369400 502212 369434
rect 502111 369344 502212 369400
rect 500924 369277 501025 369310
rect 502111 369310 502146 369344
rect 502180 369310 502212 369344
rect 502111 369277 502212 369310
rect 500924 369243 502212 369277
rect 500924 369209 500982 369243
rect 501016 369209 501072 369243
rect 501106 369209 501162 369243
rect 501196 369209 501252 369243
rect 501286 369209 501342 369243
rect 501376 369209 501432 369243
rect 501466 369209 501522 369243
rect 501556 369209 501612 369243
rect 501646 369209 501702 369243
rect 501736 369209 501792 369243
rect 501826 369209 501882 369243
rect 501916 369209 501972 369243
rect 502006 369209 502062 369243
rect 502096 369209 502212 369243
rect 500924 369090 502212 369209
rect 500924 369056 500982 369090
rect 501016 369056 501072 369090
rect 501106 369056 501162 369090
rect 501196 369056 501252 369090
rect 501286 369056 501342 369090
rect 501376 369056 501432 369090
rect 501466 369056 501522 369090
rect 501556 369056 501612 369090
rect 501646 369056 501702 369090
rect 501736 369056 501792 369090
rect 501826 369056 501882 369090
rect 501916 369056 501972 369090
rect 502006 369056 502062 369090
rect 502096 369056 502212 369090
rect 500924 369023 502212 369056
rect 500924 368994 501025 369023
rect 500924 368960 500959 368994
rect 500993 368960 501025 368994
rect 502111 368994 502212 369023
rect 500924 368904 501025 368960
rect 500924 368870 500959 368904
rect 500993 368870 501025 368904
rect 500924 368814 501025 368870
rect 500924 368780 500959 368814
rect 500993 368780 501025 368814
rect 500924 368724 501025 368780
rect 500924 368690 500959 368724
rect 500993 368690 501025 368724
rect 500924 368634 501025 368690
rect 500924 368600 500959 368634
rect 500993 368600 501025 368634
rect 500924 368544 501025 368600
rect 500924 368510 500959 368544
rect 500993 368510 501025 368544
rect 500924 368454 501025 368510
rect 500924 368420 500959 368454
rect 500993 368420 501025 368454
rect 500924 368364 501025 368420
rect 500924 368330 500959 368364
rect 500993 368330 501025 368364
rect 500924 368274 501025 368330
rect 500924 368240 500959 368274
rect 500993 368240 501025 368274
rect 500924 368184 501025 368240
rect 500924 368150 500959 368184
rect 500993 368150 501025 368184
rect 500924 368094 501025 368150
rect 500924 368060 500959 368094
rect 500993 368060 501025 368094
rect 500924 368004 501025 368060
rect 500924 367970 500959 368004
rect 500993 367970 501025 368004
rect 502111 368960 502146 368994
rect 502180 368960 502212 368994
rect 502111 368904 502212 368960
rect 502111 368870 502146 368904
rect 502180 368870 502212 368904
rect 502111 368814 502212 368870
rect 502111 368780 502146 368814
rect 502180 368780 502212 368814
rect 502111 368724 502212 368780
rect 502111 368690 502146 368724
rect 502180 368690 502212 368724
rect 502111 368634 502212 368690
rect 502111 368600 502146 368634
rect 502180 368600 502212 368634
rect 502111 368544 502212 368600
rect 502111 368510 502146 368544
rect 502180 368510 502212 368544
rect 502111 368454 502212 368510
rect 502111 368420 502146 368454
rect 502180 368420 502212 368454
rect 502111 368364 502212 368420
rect 502111 368330 502146 368364
rect 502180 368330 502212 368364
rect 502111 368274 502212 368330
rect 502111 368240 502146 368274
rect 502180 368240 502212 368274
rect 502111 368184 502212 368240
rect 502111 368150 502146 368184
rect 502180 368150 502212 368184
rect 502111 368094 502212 368150
rect 502111 368060 502146 368094
rect 502180 368060 502212 368094
rect 502111 368004 502212 368060
rect 500924 367937 501025 367970
rect 502111 367970 502146 368004
rect 502180 367970 502212 368004
rect 502111 367937 502212 367970
rect 500924 367903 502212 367937
rect 500924 367869 500982 367903
rect 501016 367869 501072 367903
rect 501106 367869 501162 367903
rect 501196 367869 501252 367903
rect 501286 367869 501342 367903
rect 501376 367869 501432 367903
rect 501466 367869 501522 367903
rect 501556 367869 501612 367903
rect 501646 367869 501702 367903
rect 501736 367869 501792 367903
rect 501826 367869 501882 367903
rect 501916 367869 501972 367903
rect 502006 367869 502062 367903
rect 502096 367869 502212 367903
rect 500924 367750 502212 367869
rect 500924 367716 500982 367750
rect 501016 367716 501072 367750
rect 501106 367716 501162 367750
rect 501196 367716 501252 367750
rect 501286 367716 501342 367750
rect 501376 367716 501432 367750
rect 501466 367716 501522 367750
rect 501556 367716 501612 367750
rect 501646 367716 501702 367750
rect 501736 367716 501792 367750
rect 501826 367716 501882 367750
rect 501916 367716 501972 367750
rect 502006 367716 502062 367750
rect 502096 367716 502212 367750
rect 500924 367683 502212 367716
rect 500924 367654 501025 367683
rect 500924 367620 500959 367654
rect 500993 367620 501025 367654
rect 502111 367654 502212 367683
rect 500924 367564 501025 367620
rect 500924 367530 500959 367564
rect 500993 367530 501025 367564
rect 500924 367474 501025 367530
rect 500924 367440 500959 367474
rect 500993 367440 501025 367474
rect 500924 367384 501025 367440
rect 500924 367350 500959 367384
rect 500993 367350 501025 367384
rect 500924 367294 501025 367350
rect 500924 367260 500959 367294
rect 500993 367260 501025 367294
rect 500924 367204 501025 367260
rect 500924 367170 500959 367204
rect 500993 367170 501025 367204
rect 500924 367114 501025 367170
rect 500924 367080 500959 367114
rect 500993 367080 501025 367114
rect 500924 367024 501025 367080
rect 500924 366990 500959 367024
rect 500993 366990 501025 367024
rect 500924 366934 501025 366990
rect 500924 366900 500959 366934
rect 500993 366900 501025 366934
rect 500924 366844 501025 366900
rect 500924 366810 500959 366844
rect 500993 366810 501025 366844
rect 500924 366754 501025 366810
rect 500924 366720 500959 366754
rect 500993 366720 501025 366754
rect 500924 366664 501025 366720
rect 500924 366630 500959 366664
rect 500993 366630 501025 366664
rect 502111 367620 502146 367654
rect 502180 367620 502212 367654
rect 502111 367564 502212 367620
rect 502111 367530 502146 367564
rect 502180 367530 502212 367564
rect 502111 367474 502212 367530
rect 502111 367440 502146 367474
rect 502180 367440 502212 367474
rect 502111 367384 502212 367440
rect 502111 367350 502146 367384
rect 502180 367350 502212 367384
rect 502111 367294 502212 367350
rect 502111 367260 502146 367294
rect 502180 367260 502212 367294
rect 502111 367204 502212 367260
rect 502111 367170 502146 367204
rect 502180 367170 502212 367204
rect 502111 367114 502212 367170
rect 502111 367080 502146 367114
rect 502180 367080 502212 367114
rect 502111 367024 502212 367080
rect 502111 366990 502146 367024
rect 502180 366990 502212 367024
rect 502111 366934 502212 366990
rect 502111 366900 502146 366934
rect 502180 366900 502212 366934
rect 502111 366844 502212 366900
rect 502111 366810 502146 366844
rect 502180 366810 502212 366844
rect 502111 366754 502212 366810
rect 502111 366720 502146 366754
rect 502180 366720 502212 366754
rect 502111 366664 502212 366720
rect 500924 366597 501025 366630
rect 502111 366630 502146 366664
rect 502180 366630 502212 366664
rect 502111 366597 502212 366630
rect 500924 366563 502212 366597
rect 500924 366529 500982 366563
rect 501016 366529 501072 366563
rect 501106 366529 501162 366563
rect 501196 366529 501252 366563
rect 501286 366529 501342 366563
rect 501376 366529 501432 366563
rect 501466 366529 501522 366563
rect 501556 366529 501612 366563
rect 501646 366529 501702 366563
rect 501736 366529 501792 366563
rect 501826 366529 501882 366563
rect 501916 366529 501972 366563
rect 502006 366529 502062 366563
rect 502096 366529 502212 366563
rect 500924 366410 502212 366529
rect 500924 366376 500982 366410
rect 501016 366376 501072 366410
rect 501106 366376 501162 366410
rect 501196 366376 501252 366410
rect 501286 366376 501342 366410
rect 501376 366376 501432 366410
rect 501466 366376 501522 366410
rect 501556 366376 501612 366410
rect 501646 366376 501702 366410
rect 501736 366376 501792 366410
rect 501826 366376 501882 366410
rect 501916 366376 501972 366410
rect 502006 366376 502062 366410
rect 502096 366376 502212 366410
rect 500924 366343 502212 366376
rect 500924 366314 501025 366343
rect 500924 366280 500959 366314
rect 500993 366280 501025 366314
rect 502111 366314 502212 366343
rect 500924 366224 501025 366280
rect 500924 366190 500959 366224
rect 500993 366190 501025 366224
rect 500924 366134 501025 366190
rect 500924 366100 500959 366134
rect 500993 366100 501025 366134
rect 500924 366044 501025 366100
rect 500924 366010 500959 366044
rect 500993 366010 501025 366044
rect 500924 365954 501025 366010
rect 500924 365920 500959 365954
rect 500993 365920 501025 365954
rect 500924 365864 501025 365920
rect 500924 365830 500959 365864
rect 500993 365830 501025 365864
rect 500924 365774 501025 365830
rect 500924 365740 500959 365774
rect 500993 365740 501025 365774
rect 500924 365684 501025 365740
rect 500924 365650 500959 365684
rect 500993 365650 501025 365684
rect 500924 365594 501025 365650
rect 500924 365560 500959 365594
rect 500993 365560 501025 365594
rect 500924 365504 501025 365560
rect 500924 365470 500959 365504
rect 500993 365470 501025 365504
rect 500924 365414 501025 365470
rect 500924 365380 500959 365414
rect 500993 365380 501025 365414
rect 500924 365324 501025 365380
rect 500924 365290 500959 365324
rect 500993 365290 501025 365324
rect 502111 366280 502146 366314
rect 502180 366280 502212 366314
rect 502111 366224 502212 366280
rect 502111 366190 502146 366224
rect 502180 366190 502212 366224
rect 502111 366134 502212 366190
rect 502111 366100 502146 366134
rect 502180 366100 502212 366134
rect 502111 366044 502212 366100
rect 502111 366010 502146 366044
rect 502180 366010 502212 366044
rect 502111 365954 502212 366010
rect 502111 365920 502146 365954
rect 502180 365920 502212 365954
rect 502111 365864 502212 365920
rect 502111 365830 502146 365864
rect 502180 365830 502212 365864
rect 502111 365774 502212 365830
rect 502111 365740 502146 365774
rect 502180 365740 502212 365774
rect 502111 365684 502212 365740
rect 502111 365650 502146 365684
rect 502180 365650 502212 365684
rect 502111 365594 502212 365650
rect 502111 365560 502146 365594
rect 502180 365560 502212 365594
rect 502111 365504 502212 365560
rect 502111 365470 502146 365504
rect 502180 365470 502212 365504
rect 502111 365414 502212 365470
rect 502111 365380 502146 365414
rect 502180 365380 502212 365414
rect 502111 365324 502212 365380
rect 500924 365257 501025 365290
rect 502111 365290 502146 365324
rect 502180 365290 502212 365324
rect 502111 365257 502212 365290
rect 500924 365223 502212 365257
rect 500924 365189 500982 365223
rect 501016 365189 501072 365223
rect 501106 365189 501162 365223
rect 501196 365189 501252 365223
rect 501286 365189 501342 365223
rect 501376 365189 501432 365223
rect 501466 365189 501522 365223
rect 501556 365189 501612 365223
rect 501646 365189 501702 365223
rect 501736 365189 501792 365223
rect 501826 365189 501882 365223
rect 501916 365189 501972 365223
rect 502006 365189 502062 365223
rect 502096 365189 502212 365223
rect 500924 365070 502212 365189
rect 500924 365036 500982 365070
rect 501016 365036 501072 365070
rect 501106 365036 501162 365070
rect 501196 365036 501252 365070
rect 501286 365036 501342 365070
rect 501376 365036 501432 365070
rect 501466 365036 501522 365070
rect 501556 365036 501612 365070
rect 501646 365036 501702 365070
rect 501736 365036 501792 365070
rect 501826 365036 501882 365070
rect 501916 365036 501972 365070
rect 502006 365036 502062 365070
rect 502096 365036 502212 365070
rect 500924 365003 502212 365036
rect 500924 364974 501025 365003
rect 500924 364940 500959 364974
rect 500993 364940 501025 364974
rect 502111 364974 502212 365003
rect 500924 364884 501025 364940
rect 500924 364850 500959 364884
rect 500993 364850 501025 364884
rect 500924 364794 501025 364850
rect 500924 364760 500959 364794
rect 500993 364760 501025 364794
rect 500924 364704 501025 364760
rect 500924 364670 500959 364704
rect 500993 364670 501025 364704
rect 500924 364614 501025 364670
rect 500924 364580 500959 364614
rect 500993 364580 501025 364614
rect 500924 364524 501025 364580
rect 500924 364490 500959 364524
rect 500993 364490 501025 364524
rect 500924 364434 501025 364490
rect 500924 364400 500959 364434
rect 500993 364400 501025 364434
rect 500924 364344 501025 364400
rect 500924 364310 500959 364344
rect 500993 364310 501025 364344
rect 500924 364254 501025 364310
rect 500924 364220 500959 364254
rect 500993 364220 501025 364254
rect 500924 364164 501025 364220
rect 500924 364130 500959 364164
rect 500993 364130 501025 364164
rect 500924 364074 501025 364130
rect 500924 364040 500959 364074
rect 500993 364040 501025 364074
rect 500924 363984 501025 364040
rect 500924 363950 500959 363984
rect 500993 363950 501025 363984
rect 502111 364940 502146 364974
rect 502180 364940 502212 364974
rect 502111 364884 502212 364940
rect 502111 364850 502146 364884
rect 502180 364850 502212 364884
rect 502111 364794 502212 364850
rect 502111 364760 502146 364794
rect 502180 364760 502212 364794
rect 502111 364704 502212 364760
rect 502111 364670 502146 364704
rect 502180 364670 502212 364704
rect 502111 364614 502212 364670
rect 502111 364580 502146 364614
rect 502180 364580 502212 364614
rect 502111 364524 502212 364580
rect 502111 364490 502146 364524
rect 502180 364490 502212 364524
rect 502111 364434 502212 364490
rect 502111 364400 502146 364434
rect 502180 364400 502212 364434
rect 502111 364344 502212 364400
rect 502111 364310 502146 364344
rect 502180 364310 502212 364344
rect 502111 364254 502212 364310
rect 502111 364220 502146 364254
rect 502180 364220 502212 364254
rect 502111 364164 502212 364220
rect 502111 364130 502146 364164
rect 502180 364130 502212 364164
rect 502111 364074 502212 364130
rect 502111 364040 502146 364074
rect 502180 364040 502212 364074
rect 502111 363984 502212 364040
rect 500924 363917 501025 363950
rect 502111 363950 502146 363984
rect 502180 363950 502212 363984
rect 502111 363917 502212 363950
rect 500924 363883 502212 363917
rect 500924 363849 500982 363883
rect 501016 363849 501072 363883
rect 501106 363849 501162 363883
rect 501196 363849 501252 363883
rect 501286 363849 501342 363883
rect 501376 363849 501432 363883
rect 501466 363849 501522 363883
rect 501556 363849 501612 363883
rect 501646 363849 501702 363883
rect 501736 363849 501792 363883
rect 501826 363849 501882 363883
rect 501916 363849 501972 363883
rect 502006 363849 502062 363883
rect 502096 363849 502212 363883
rect 500924 363730 502212 363849
rect 500924 363696 500982 363730
rect 501016 363696 501072 363730
rect 501106 363696 501162 363730
rect 501196 363696 501252 363730
rect 501286 363696 501342 363730
rect 501376 363696 501432 363730
rect 501466 363696 501522 363730
rect 501556 363696 501612 363730
rect 501646 363696 501702 363730
rect 501736 363696 501792 363730
rect 501826 363696 501882 363730
rect 501916 363696 501972 363730
rect 502006 363696 502062 363730
rect 502096 363696 502212 363730
rect 500924 363663 502212 363696
rect 500924 363634 501025 363663
rect 500924 363600 500959 363634
rect 500993 363600 501025 363634
rect 502111 363634 502212 363663
rect 500924 363544 501025 363600
rect 500924 363510 500959 363544
rect 500993 363510 501025 363544
rect 500924 363454 501025 363510
rect 500924 363420 500959 363454
rect 500993 363420 501025 363454
rect 500924 363364 501025 363420
rect 500924 363330 500959 363364
rect 500993 363330 501025 363364
rect 500924 363274 501025 363330
rect 500924 363240 500959 363274
rect 500993 363240 501025 363274
rect 500924 363184 501025 363240
rect 500924 363150 500959 363184
rect 500993 363150 501025 363184
rect 500924 363094 501025 363150
rect 500924 363060 500959 363094
rect 500993 363060 501025 363094
rect 500924 363004 501025 363060
rect 500924 362970 500959 363004
rect 500993 362970 501025 363004
rect 500924 362914 501025 362970
rect 500924 362880 500959 362914
rect 500993 362880 501025 362914
rect 500924 362824 501025 362880
rect 500924 362790 500959 362824
rect 500993 362790 501025 362824
rect 500924 362734 501025 362790
rect 500924 362700 500959 362734
rect 500993 362700 501025 362734
rect 500924 362644 501025 362700
rect 500924 362610 500959 362644
rect 500993 362610 501025 362644
rect 502111 363600 502146 363634
rect 502180 363600 502212 363634
rect 502111 363544 502212 363600
rect 502111 363510 502146 363544
rect 502180 363510 502212 363544
rect 502111 363454 502212 363510
rect 502111 363420 502146 363454
rect 502180 363420 502212 363454
rect 502111 363364 502212 363420
rect 502111 363330 502146 363364
rect 502180 363330 502212 363364
rect 502111 363274 502212 363330
rect 502111 363240 502146 363274
rect 502180 363240 502212 363274
rect 502111 363184 502212 363240
rect 502111 363150 502146 363184
rect 502180 363150 502212 363184
rect 502111 363094 502212 363150
rect 502111 363060 502146 363094
rect 502180 363060 502212 363094
rect 502111 363004 502212 363060
rect 502111 362970 502146 363004
rect 502180 362970 502212 363004
rect 502111 362914 502212 362970
rect 502111 362880 502146 362914
rect 502180 362880 502212 362914
rect 502111 362824 502212 362880
rect 502111 362790 502146 362824
rect 502180 362790 502212 362824
rect 502111 362734 502212 362790
rect 502111 362700 502146 362734
rect 502180 362700 502212 362734
rect 502111 362644 502212 362700
rect 500924 362577 501025 362610
rect 502111 362610 502146 362644
rect 502180 362610 502212 362644
rect 502111 362577 502212 362610
rect 500924 362543 502212 362577
rect 500924 362509 500982 362543
rect 501016 362509 501072 362543
rect 501106 362509 501162 362543
rect 501196 362509 501252 362543
rect 501286 362509 501342 362543
rect 501376 362509 501432 362543
rect 501466 362509 501522 362543
rect 501556 362509 501612 362543
rect 501646 362509 501702 362543
rect 501736 362509 501792 362543
rect 501826 362509 501882 362543
rect 501916 362509 501972 362543
rect 502006 362509 502062 362543
rect 502096 362509 502212 362543
rect 500924 362476 502212 362509
rect 504684 373110 505972 373144
rect 504684 373076 504742 373110
rect 504776 373076 504832 373110
rect 504866 373076 504922 373110
rect 504956 373076 505012 373110
rect 505046 373076 505102 373110
rect 505136 373076 505192 373110
rect 505226 373076 505282 373110
rect 505316 373076 505372 373110
rect 505406 373076 505462 373110
rect 505496 373076 505552 373110
rect 505586 373076 505642 373110
rect 505676 373076 505732 373110
rect 505766 373076 505822 373110
rect 505856 373076 505972 373110
rect 504684 373043 505972 373076
rect 504684 373014 504785 373043
rect 504684 372980 504719 373014
rect 504753 372980 504785 373014
rect 505871 373014 505972 373043
rect 504684 372924 504785 372980
rect 504684 372890 504719 372924
rect 504753 372890 504785 372924
rect 504684 372834 504785 372890
rect 504684 372800 504719 372834
rect 504753 372800 504785 372834
rect 504684 372744 504785 372800
rect 504684 372710 504719 372744
rect 504753 372710 504785 372744
rect 504684 372654 504785 372710
rect 504684 372620 504719 372654
rect 504753 372620 504785 372654
rect 504684 372564 504785 372620
rect 504684 372530 504719 372564
rect 504753 372530 504785 372564
rect 504684 372474 504785 372530
rect 504684 372440 504719 372474
rect 504753 372440 504785 372474
rect 504684 372384 504785 372440
rect 504684 372350 504719 372384
rect 504753 372350 504785 372384
rect 504684 372294 504785 372350
rect 504684 372260 504719 372294
rect 504753 372260 504785 372294
rect 504684 372204 504785 372260
rect 504684 372170 504719 372204
rect 504753 372170 504785 372204
rect 504684 372114 504785 372170
rect 504684 372080 504719 372114
rect 504753 372080 504785 372114
rect 504684 372024 504785 372080
rect 504684 371990 504719 372024
rect 504753 371990 504785 372024
rect 505871 372980 505906 373014
rect 505940 372980 505972 373014
rect 505871 372924 505972 372980
rect 505871 372890 505906 372924
rect 505940 372890 505972 372924
rect 505871 372834 505972 372890
rect 505871 372800 505906 372834
rect 505940 372800 505972 372834
rect 505871 372744 505972 372800
rect 505871 372710 505906 372744
rect 505940 372710 505972 372744
rect 505871 372654 505972 372710
rect 505871 372620 505906 372654
rect 505940 372620 505972 372654
rect 505871 372564 505972 372620
rect 505871 372530 505906 372564
rect 505940 372530 505972 372564
rect 505871 372474 505972 372530
rect 505871 372440 505906 372474
rect 505940 372440 505972 372474
rect 505871 372384 505972 372440
rect 505871 372350 505906 372384
rect 505940 372350 505972 372384
rect 505871 372294 505972 372350
rect 505871 372260 505906 372294
rect 505940 372260 505972 372294
rect 505871 372204 505972 372260
rect 505871 372170 505906 372204
rect 505940 372170 505972 372204
rect 505871 372114 505972 372170
rect 505871 372080 505906 372114
rect 505940 372080 505972 372114
rect 505871 372024 505972 372080
rect 504684 371957 504785 371990
rect 505871 371990 505906 372024
rect 505940 371990 505972 372024
rect 505871 371957 505972 371990
rect 504684 371923 505972 371957
rect 504684 371889 504742 371923
rect 504776 371889 504832 371923
rect 504866 371889 504922 371923
rect 504956 371889 505012 371923
rect 505046 371889 505102 371923
rect 505136 371889 505192 371923
rect 505226 371889 505282 371923
rect 505316 371889 505372 371923
rect 505406 371889 505462 371923
rect 505496 371889 505552 371923
rect 505586 371889 505642 371923
rect 505676 371889 505732 371923
rect 505766 371889 505822 371923
rect 505856 371889 505972 371923
rect 504684 371770 505972 371889
rect 504684 371736 504742 371770
rect 504776 371736 504832 371770
rect 504866 371736 504922 371770
rect 504956 371736 505012 371770
rect 505046 371736 505102 371770
rect 505136 371736 505192 371770
rect 505226 371736 505282 371770
rect 505316 371736 505372 371770
rect 505406 371736 505462 371770
rect 505496 371736 505552 371770
rect 505586 371736 505642 371770
rect 505676 371736 505732 371770
rect 505766 371736 505822 371770
rect 505856 371736 505972 371770
rect 504684 371703 505972 371736
rect 504684 371674 504785 371703
rect 504684 371640 504719 371674
rect 504753 371640 504785 371674
rect 505871 371674 505972 371703
rect 504684 371584 504785 371640
rect 504684 371550 504719 371584
rect 504753 371550 504785 371584
rect 504684 371494 504785 371550
rect 504684 371460 504719 371494
rect 504753 371460 504785 371494
rect 504684 371404 504785 371460
rect 504684 371370 504719 371404
rect 504753 371370 504785 371404
rect 504684 371314 504785 371370
rect 504684 371280 504719 371314
rect 504753 371280 504785 371314
rect 504684 371224 504785 371280
rect 504684 371190 504719 371224
rect 504753 371190 504785 371224
rect 504684 371134 504785 371190
rect 504684 371100 504719 371134
rect 504753 371100 504785 371134
rect 504684 371044 504785 371100
rect 504684 371010 504719 371044
rect 504753 371010 504785 371044
rect 504684 370954 504785 371010
rect 504684 370920 504719 370954
rect 504753 370920 504785 370954
rect 504684 370864 504785 370920
rect 504684 370830 504719 370864
rect 504753 370830 504785 370864
rect 504684 370774 504785 370830
rect 504684 370740 504719 370774
rect 504753 370740 504785 370774
rect 504684 370684 504785 370740
rect 504684 370650 504719 370684
rect 504753 370650 504785 370684
rect 505871 371640 505906 371674
rect 505940 371640 505972 371674
rect 505871 371584 505972 371640
rect 505871 371550 505906 371584
rect 505940 371550 505972 371584
rect 505871 371494 505972 371550
rect 505871 371460 505906 371494
rect 505940 371460 505972 371494
rect 505871 371404 505972 371460
rect 505871 371370 505906 371404
rect 505940 371370 505972 371404
rect 505871 371314 505972 371370
rect 505871 371280 505906 371314
rect 505940 371280 505972 371314
rect 505871 371224 505972 371280
rect 505871 371190 505906 371224
rect 505940 371190 505972 371224
rect 505871 371134 505972 371190
rect 505871 371100 505906 371134
rect 505940 371100 505972 371134
rect 505871 371044 505972 371100
rect 505871 371010 505906 371044
rect 505940 371010 505972 371044
rect 505871 370954 505972 371010
rect 505871 370920 505906 370954
rect 505940 370920 505972 370954
rect 505871 370864 505972 370920
rect 505871 370830 505906 370864
rect 505940 370830 505972 370864
rect 505871 370774 505972 370830
rect 505871 370740 505906 370774
rect 505940 370740 505972 370774
rect 505871 370684 505972 370740
rect 504684 370617 504785 370650
rect 505871 370650 505906 370684
rect 505940 370650 505972 370684
rect 505871 370617 505972 370650
rect 504684 370583 505972 370617
rect 504684 370549 504742 370583
rect 504776 370549 504832 370583
rect 504866 370549 504922 370583
rect 504956 370549 505012 370583
rect 505046 370549 505102 370583
rect 505136 370549 505192 370583
rect 505226 370549 505282 370583
rect 505316 370549 505372 370583
rect 505406 370549 505462 370583
rect 505496 370549 505552 370583
rect 505586 370549 505642 370583
rect 505676 370549 505732 370583
rect 505766 370549 505822 370583
rect 505856 370549 505972 370583
rect 504684 370430 505972 370549
rect 504684 370396 504742 370430
rect 504776 370396 504832 370430
rect 504866 370396 504922 370430
rect 504956 370396 505012 370430
rect 505046 370396 505102 370430
rect 505136 370396 505192 370430
rect 505226 370396 505282 370430
rect 505316 370396 505372 370430
rect 505406 370396 505462 370430
rect 505496 370396 505552 370430
rect 505586 370396 505642 370430
rect 505676 370396 505732 370430
rect 505766 370396 505822 370430
rect 505856 370396 505972 370430
rect 504684 370363 505972 370396
rect 504684 370334 504785 370363
rect 504684 370300 504719 370334
rect 504753 370300 504785 370334
rect 505871 370334 505972 370363
rect 504684 370244 504785 370300
rect 504684 370210 504719 370244
rect 504753 370210 504785 370244
rect 504684 370154 504785 370210
rect 504684 370120 504719 370154
rect 504753 370120 504785 370154
rect 504684 370064 504785 370120
rect 504684 370030 504719 370064
rect 504753 370030 504785 370064
rect 504684 369974 504785 370030
rect 504684 369940 504719 369974
rect 504753 369940 504785 369974
rect 504684 369884 504785 369940
rect 504684 369850 504719 369884
rect 504753 369850 504785 369884
rect 504684 369794 504785 369850
rect 504684 369760 504719 369794
rect 504753 369760 504785 369794
rect 504684 369704 504785 369760
rect 504684 369670 504719 369704
rect 504753 369670 504785 369704
rect 504684 369614 504785 369670
rect 504684 369580 504719 369614
rect 504753 369580 504785 369614
rect 504684 369524 504785 369580
rect 504684 369490 504719 369524
rect 504753 369490 504785 369524
rect 504684 369434 504785 369490
rect 504684 369400 504719 369434
rect 504753 369400 504785 369434
rect 504684 369344 504785 369400
rect 504684 369310 504719 369344
rect 504753 369310 504785 369344
rect 505871 370300 505906 370334
rect 505940 370300 505972 370334
rect 505871 370244 505972 370300
rect 505871 370210 505906 370244
rect 505940 370210 505972 370244
rect 505871 370154 505972 370210
rect 505871 370120 505906 370154
rect 505940 370120 505972 370154
rect 505871 370064 505972 370120
rect 505871 370030 505906 370064
rect 505940 370030 505972 370064
rect 505871 369974 505972 370030
rect 505871 369940 505906 369974
rect 505940 369940 505972 369974
rect 505871 369884 505972 369940
rect 505871 369850 505906 369884
rect 505940 369850 505972 369884
rect 505871 369794 505972 369850
rect 505871 369760 505906 369794
rect 505940 369760 505972 369794
rect 505871 369704 505972 369760
rect 505871 369670 505906 369704
rect 505940 369670 505972 369704
rect 505871 369614 505972 369670
rect 505871 369580 505906 369614
rect 505940 369580 505972 369614
rect 505871 369524 505972 369580
rect 505871 369490 505906 369524
rect 505940 369490 505972 369524
rect 505871 369434 505972 369490
rect 505871 369400 505906 369434
rect 505940 369400 505972 369434
rect 505871 369344 505972 369400
rect 504684 369277 504785 369310
rect 505871 369310 505906 369344
rect 505940 369310 505972 369344
rect 505871 369277 505972 369310
rect 504684 369243 505972 369277
rect 504684 369209 504742 369243
rect 504776 369209 504832 369243
rect 504866 369209 504922 369243
rect 504956 369209 505012 369243
rect 505046 369209 505102 369243
rect 505136 369209 505192 369243
rect 505226 369209 505282 369243
rect 505316 369209 505372 369243
rect 505406 369209 505462 369243
rect 505496 369209 505552 369243
rect 505586 369209 505642 369243
rect 505676 369209 505732 369243
rect 505766 369209 505822 369243
rect 505856 369209 505972 369243
rect 504684 369090 505972 369209
rect 504684 369056 504742 369090
rect 504776 369056 504832 369090
rect 504866 369056 504922 369090
rect 504956 369056 505012 369090
rect 505046 369056 505102 369090
rect 505136 369056 505192 369090
rect 505226 369056 505282 369090
rect 505316 369056 505372 369090
rect 505406 369056 505462 369090
rect 505496 369056 505552 369090
rect 505586 369056 505642 369090
rect 505676 369056 505732 369090
rect 505766 369056 505822 369090
rect 505856 369056 505972 369090
rect 504684 369023 505972 369056
rect 504684 368994 504785 369023
rect 504684 368960 504719 368994
rect 504753 368960 504785 368994
rect 505871 368994 505972 369023
rect 504684 368904 504785 368960
rect 504684 368870 504719 368904
rect 504753 368870 504785 368904
rect 504684 368814 504785 368870
rect 504684 368780 504719 368814
rect 504753 368780 504785 368814
rect 504684 368724 504785 368780
rect 504684 368690 504719 368724
rect 504753 368690 504785 368724
rect 504684 368634 504785 368690
rect 504684 368600 504719 368634
rect 504753 368600 504785 368634
rect 504684 368544 504785 368600
rect 504684 368510 504719 368544
rect 504753 368510 504785 368544
rect 504684 368454 504785 368510
rect 504684 368420 504719 368454
rect 504753 368420 504785 368454
rect 504684 368364 504785 368420
rect 504684 368330 504719 368364
rect 504753 368330 504785 368364
rect 504684 368274 504785 368330
rect 504684 368240 504719 368274
rect 504753 368240 504785 368274
rect 504684 368184 504785 368240
rect 504684 368150 504719 368184
rect 504753 368150 504785 368184
rect 504684 368094 504785 368150
rect 504684 368060 504719 368094
rect 504753 368060 504785 368094
rect 504684 368004 504785 368060
rect 504684 367970 504719 368004
rect 504753 367970 504785 368004
rect 505871 368960 505906 368994
rect 505940 368960 505972 368994
rect 505871 368904 505972 368960
rect 505871 368870 505906 368904
rect 505940 368870 505972 368904
rect 505871 368814 505972 368870
rect 505871 368780 505906 368814
rect 505940 368780 505972 368814
rect 505871 368724 505972 368780
rect 505871 368690 505906 368724
rect 505940 368690 505972 368724
rect 505871 368634 505972 368690
rect 505871 368600 505906 368634
rect 505940 368600 505972 368634
rect 505871 368544 505972 368600
rect 505871 368510 505906 368544
rect 505940 368510 505972 368544
rect 505871 368454 505972 368510
rect 505871 368420 505906 368454
rect 505940 368420 505972 368454
rect 505871 368364 505972 368420
rect 505871 368330 505906 368364
rect 505940 368330 505972 368364
rect 505871 368274 505972 368330
rect 505871 368240 505906 368274
rect 505940 368240 505972 368274
rect 505871 368184 505972 368240
rect 505871 368150 505906 368184
rect 505940 368150 505972 368184
rect 505871 368094 505972 368150
rect 505871 368060 505906 368094
rect 505940 368060 505972 368094
rect 505871 368004 505972 368060
rect 504684 367937 504785 367970
rect 505871 367970 505906 368004
rect 505940 367970 505972 368004
rect 505871 367937 505972 367970
rect 504684 367903 505972 367937
rect 504684 367869 504742 367903
rect 504776 367869 504832 367903
rect 504866 367869 504922 367903
rect 504956 367869 505012 367903
rect 505046 367869 505102 367903
rect 505136 367869 505192 367903
rect 505226 367869 505282 367903
rect 505316 367869 505372 367903
rect 505406 367869 505462 367903
rect 505496 367869 505552 367903
rect 505586 367869 505642 367903
rect 505676 367869 505732 367903
rect 505766 367869 505822 367903
rect 505856 367869 505972 367903
rect 504684 367750 505972 367869
rect 504684 367716 504742 367750
rect 504776 367716 504832 367750
rect 504866 367716 504922 367750
rect 504956 367716 505012 367750
rect 505046 367716 505102 367750
rect 505136 367716 505192 367750
rect 505226 367716 505282 367750
rect 505316 367716 505372 367750
rect 505406 367716 505462 367750
rect 505496 367716 505552 367750
rect 505586 367716 505642 367750
rect 505676 367716 505732 367750
rect 505766 367716 505822 367750
rect 505856 367716 505972 367750
rect 504684 367683 505972 367716
rect 504684 367654 504785 367683
rect 504684 367620 504719 367654
rect 504753 367620 504785 367654
rect 505871 367654 505972 367683
rect 504684 367564 504785 367620
rect 504684 367530 504719 367564
rect 504753 367530 504785 367564
rect 504684 367474 504785 367530
rect 504684 367440 504719 367474
rect 504753 367440 504785 367474
rect 504684 367384 504785 367440
rect 504684 367350 504719 367384
rect 504753 367350 504785 367384
rect 504684 367294 504785 367350
rect 504684 367260 504719 367294
rect 504753 367260 504785 367294
rect 504684 367204 504785 367260
rect 504684 367170 504719 367204
rect 504753 367170 504785 367204
rect 504684 367114 504785 367170
rect 504684 367080 504719 367114
rect 504753 367080 504785 367114
rect 504684 367024 504785 367080
rect 504684 366990 504719 367024
rect 504753 366990 504785 367024
rect 504684 366934 504785 366990
rect 504684 366900 504719 366934
rect 504753 366900 504785 366934
rect 504684 366844 504785 366900
rect 504684 366810 504719 366844
rect 504753 366810 504785 366844
rect 504684 366754 504785 366810
rect 504684 366720 504719 366754
rect 504753 366720 504785 366754
rect 504684 366664 504785 366720
rect 504684 366630 504719 366664
rect 504753 366630 504785 366664
rect 505871 367620 505906 367654
rect 505940 367620 505972 367654
rect 505871 367564 505972 367620
rect 505871 367530 505906 367564
rect 505940 367530 505972 367564
rect 505871 367474 505972 367530
rect 505871 367440 505906 367474
rect 505940 367440 505972 367474
rect 505871 367384 505972 367440
rect 505871 367350 505906 367384
rect 505940 367350 505972 367384
rect 505871 367294 505972 367350
rect 505871 367260 505906 367294
rect 505940 367260 505972 367294
rect 505871 367204 505972 367260
rect 505871 367170 505906 367204
rect 505940 367170 505972 367204
rect 505871 367114 505972 367170
rect 505871 367080 505906 367114
rect 505940 367080 505972 367114
rect 505871 367024 505972 367080
rect 505871 366990 505906 367024
rect 505940 366990 505972 367024
rect 505871 366934 505972 366990
rect 505871 366900 505906 366934
rect 505940 366900 505972 366934
rect 505871 366844 505972 366900
rect 505871 366810 505906 366844
rect 505940 366810 505972 366844
rect 505871 366754 505972 366810
rect 505871 366720 505906 366754
rect 505940 366720 505972 366754
rect 505871 366664 505972 366720
rect 504684 366597 504785 366630
rect 505871 366630 505906 366664
rect 505940 366630 505972 366664
rect 505871 366597 505972 366630
rect 504684 366563 505972 366597
rect 504684 366529 504742 366563
rect 504776 366529 504832 366563
rect 504866 366529 504922 366563
rect 504956 366529 505012 366563
rect 505046 366529 505102 366563
rect 505136 366529 505192 366563
rect 505226 366529 505282 366563
rect 505316 366529 505372 366563
rect 505406 366529 505462 366563
rect 505496 366529 505552 366563
rect 505586 366529 505642 366563
rect 505676 366529 505732 366563
rect 505766 366529 505822 366563
rect 505856 366529 505972 366563
rect 504684 366410 505972 366529
rect 504684 366376 504742 366410
rect 504776 366376 504832 366410
rect 504866 366376 504922 366410
rect 504956 366376 505012 366410
rect 505046 366376 505102 366410
rect 505136 366376 505192 366410
rect 505226 366376 505282 366410
rect 505316 366376 505372 366410
rect 505406 366376 505462 366410
rect 505496 366376 505552 366410
rect 505586 366376 505642 366410
rect 505676 366376 505732 366410
rect 505766 366376 505822 366410
rect 505856 366376 505972 366410
rect 504684 366343 505972 366376
rect 504684 366314 504785 366343
rect 504684 366280 504719 366314
rect 504753 366280 504785 366314
rect 505871 366314 505972 366343
rect 504684 366224 504785 366280
rect 504684 366190 504719 366224
rect 504753 366190 504785 366224
rect 504684 366134 504785 366190
rect 504684 366100 504719 366134
rect 504753 366100 504785 366134
rect 504684 366044 504785 366100
rect 504684 366010 504719 366044
rect 504753 366010 504785 366044
rect 504684 365954 504785 366010
rect 504684 365920 504719 365954
rect 504753 365920 504785 365954
rect 504684 365864 504785 365920
rect 504684 365830 504719 365864
rect 504753 365830 504785 365864
rect 504684 365774 504785 365830
rect 504684 365740 504719 365774
rect 504753 365740 504785 365774
rect 504684 365684 504785 365740
rect 504684 365650 504719 365684
rect 504753 365650 504785 365684
rect 504684 365594 504785 365650
rect 504684 365560 504719 365594
rect 504753 365560 504785 365594
rect 504684 365504 504785 365560
rect 504684 365470 504719 365504
rect 504753 365470 504785 365504
rect 504684 365414 504785 365470
rect 504684 365380 504719 365414
rect 504753 365380 504785 365414
rect 504684 365324 504785 365380
rect 504684 365290 504719 365324
rect 504753 365290 504785 365324
rect 505871 366280 505906 366314
rect 505940 366280 505972 366314
rect 505871 366224 505972 366280
rect 505871 366190 505906 366224
rect 505940 366190 505972 366224
rect 505871 366134 505972 366190
rect 505871 366100 505906 366134
rect 505940 366100 505972 366134
rect 505871 366044 505972 366100
rect 505871 366010 505906 366044
rect 505940 366010 505972 366044
rect 505871 365954 505972 366010
rect 505871 365920 505906 365954
rect 505940 365920 505972 365954
rect 505871 365864 505972 365920
rect 505871 365830 505906 365864
rect 505940 365830 505972 365864
rect 505871 365774 505972 365830
rect 505871 365740 505906 365774
rect 505940 365740 505972 365774
rect 505871 365684 505972 365740
rect 505871 365650 505906 365684
rect 505940 365650 505972 365684
rect 505871 365594 505972 365650
rect 505871 365560 505906 365594
rect 505940 365560 505972 365594
rect 505871 365504 505972 365560
rect 505871 365470 505906 365504
rect 505940 365470 505972 365504
rect 505871 365414 505972 365470
rect 505871 365380 505906 365414
rect 505940 365380 505972 365414
rect 505871 365324 505972 365380
rect 504684 365257 504785 365290
rect 505871 365290 505906 365324
rect 505940 365290 505972 365324
rect 505871 365257 505972 365290
rect 504684 365223 505972 365257
rect 504684 365189 504742 365223
rect 504776 365189 504832 365223
rect 504866 365189 504922 365223
rect 504956 365189 505012 365223
rect 505046 365189 505102 365223
rect 505136 365189 505192 365223
rect 505226 365189 505282 365223
rect 505316 365189 505372 365223
rect 505406 365189 505462 365223
rect 505496 365189 505552 365223
rect 505586 365189 505642 365223
rect 505676 365189 505732 365223
rect 505766 365189 505822 365223
rect 505856 365189 505972 365223
rect 504684 365070 505972 365189
rect 504684 365036 504742 365070
rect 504776 365036 504832 365070
rect 504866 365036 504922 365070
rect 504956 365036 505012 365070
rect 505046 365036 505102 365070
rect 505136 365036 505192 365070
rect 505226 365036 505282 365070
rect 505316 365036 505372 365070
rect 505406 365036 505462 365070
rect 505496 365036 505552 365070
rect 505586 365036 505642 365070
rect 505676 365036 505732 365070
rect 505766 365036 505822 365070
rect 505856 365036 505972 365070
rect 504684 365003 505972 365036
rect 504684 364974 504785 365003
rect 504684 364940 504719 364974
rect 504753 364940 504785 364974
rect 505871 364974 505972 365003
rect 504684 364884 504785 364940
rect 504684 364850 504719 364884
rect 504753 364850 504785 364884
rect 504684 364794 504785 364850
rect 504684 364760 504719 364794
rect 504753 364760 504785 364794
rect 504684 364704 504785 364760
rect 504684 364670 504719 364704
rect 504753 364670 504785 364704
rect 504684 364614 504785 364670
rect 504684 364580 504719 364614
rect 504753 364580 504785 364614
rect 504684 364524 504785 364580
rect 504684 364490 504719 364524
rect 504753 364490 504785 364524
rect 504684 364434 504785 364490
rect 504684 364400 504719 364434
rect 504753 364400 504785 364434
rect 504684 364344 504785 364400
rect 504684 364310 504719 364344
rect 504753 364310 504785 364344
rect 504684 364254 504785 364310
rect 504684 364220 504719 364254
rect 504753 364220 504785 364254
rect 504684 364164 504785 364220
rect 504684 364130 504719 364164
rect 504753 364130 504785 364164
rect 504684 364074 504785 364130
rect 504684 364040 504719 364074
rect 504753 364040 504785 364074
rect 504684 363984 504785 364040
rect 504684 363950 504719 363984
rect 504753 363950 504785 363984
rect 505871 364940 505906 364974
rect 505940 364940 505972 364974
rect 505871 364884 505972 364940
rect 505871 364850 505906 364884
rect 505940 364850 505972 364884
rect 505871 364794 505972 364850
rect 505871 364760 505906 364794
rect 505940 364760 505972 364794
rect 505871 364704 505972 364760
rect 505871 364670 505906 364704
rect 505940 364670 505972 364704
rect 505871 364614 505972 364670
rect 505871 364580 505906 364614
rect 505940 364580 505972 364614
rect 505871 364524 505972 364580
rect 505871 364490 505906 364524
rect 505940 364490 505972 364524
rect 505871 364434 505972 364490
rect 505871 364400 505906 364434
rect 505940 364400 505972 364434
rect 505871 364344 505972 364400
rect 505871 364310 505906 364344
rect 505940 364310 505972 364344
rect 505871 364254 505972 364310
rect 505871 364220 505906 364254
rect 505940 364220 505972 364254
rect 505871 364164 505972 364220
rect 505871 364130 505906 364164
rect 505940 364130 505972 364164
rect 505871 364074 505972 364130
rect 505871 364040 505906 364074
rect 505940 364040 505972 364074
rect 505871 363984 505972 364040
rect 504684 363917 504785 363950
rect 505871 363950 505906 363984
rect 505940 363950 505972 363984
rect 505871 363917 505972 363950
rect 504684 363883 505972 363917
rect 504684 363849 504742 363883
rect 504776 363849 504832 363883
rect 504866 363849 504922 363883
rect 504956 363849 505012 363883
rect 505046 363849 505102 363883
rect 505136 363849 505192 363883
rect 505226 363849 505282 363883
rect 505316 363849 505372 363883
rect 505406 363849 505462 363883
rect 505496 363849 505552 363883
rect 505586 363849 505642 363883
rect 505676 363849 505732 363883
rect 505766 363849 505822 363883
rect 505856 363849 505972 363883
rect 504684 363730 505972 363849
rect 504684 363696 504742 363730
rect 504776 363696 504832 363730
rect 504866 363696 504922 363730
rect 504956 363696 505012 363730
rect 505046 363696 505102 363730
rect 505136 363696 505192 363730
rect 505226 363696 505282 363730
rect 505316 363696 505372 363730
rect 505406 363696 505462 363730
rect 505496 363696 505552 363730
rect 505586 363696 505642 363730
rect 505676 363696 505732 363730
rect 505766 363696 505822 363730
rect 505856 363696 505972 363730
rect 504684 363663 505972 363696
rect 504684 363634 504785 363663
rect 504684 363600 504719 363634
rect 504753 363600 504785 363634
rect 505871 363634 505972 363663
rect 504684 363544 504785 363600
rect 504684 363510 504719 363544
rect 504753 363510 504785 363544
rect 504684 363454 504785 363510
rect 504684 363420 504719 363454
rect 504753 363420 504785 363454
rect 504684 363364 504785 363420
rect 504684 363330 504719 363364
rect 504753 363330 504785 363364
rect 504684 363274 504785 363330
rect 504684 363240 504719 363274
rect 504753 363240 504785 363274
rect 504684 363184 504785 363240
rect 504684 363150 504719 363184
rect 504753 363150 504785 363184
rect 504684 363094 504785 363150
rect 504684 363060 504719 363094
rect 504753 363060 504785 363094
rect 504684 363004 504785 363060
rect 504684 362970 504719 363004
rect 504753 362970 504785 363004
rect 504684 362914 504785 362970
rect 504684 362880 504719 362914
rect 504753 362880 504785 362914
rect 504684 362824 504785 362880
rect 504684 362790 504719 362824
rect 504753 362790 504785 362824
rect 504684 362734 504785 362790
rect 504684 362700 504719 362734
rect 504753 362700 504785 362734
rect 504684 362644 504785 362700
rect 504684 362610 504719 362644
rect 504753 362610 504785 362644
rect 505871 363600 505906 363634
rect 505940 363600 505972 363634
rect 505871 363544 505972 363600
rect 505871 363510 505906 363544
rect 505940 363510 505972 363544
rect 505871 363454 505972 363510
rect 505871 363420 505906 363454
rect 505940 363420 505972 363454
rect 505871 363364 505972 363420
rect 505871 363330 505906 363364
rect 505940 363330 505972 363364
rect 505871 363274 505972 363330
rect 505871 363240 505906 363274
rect 505940 363240 505972 363274
rect 505871 363184 505972 363240
rect 505871 363150 505906 363184
rect 505940 363150 505972 363184
rect 505871 363094 505972 363150
rect 505871 363060 505906 363094
rect 505940 363060 505972 363094
rect 505871 363004 505972 363060
rect 505871 362970 505906 363004
rect 505940 362970 505972 363004
rect 505871 362914 505972 362970
rect 505871 362880 505906 362914
rect 505940 362880 505972 362914
rect 505871 362824 505972 362880
rect 505871 362790 505906 362824
rect 505940 362790 505972 362824
rect 505871 362734 505972 362790
rect 505871 362700 505906 362734
rect 505940 362700 505972 362734
rect 505871 362644 505972 362700
rect 504684 362577 504785 362610
rect 505871 362610 505906 362644
rect 505940 362610 505972 362644
rect 505871 362577 505972 362610
rect 504684 362543 505972 362577
rect 504684 362509 504742 362543
rect 504776 362509 504832 362543
rect 504866 362509 504922 362543
rect 504956 362509 505012 362543
rect 505046 362509 505102 362543
rect 505136 362509 505192 362543
rect 505226 362509 505282 362543
rect 505316 362509 505372 362543
rect 505406 362509 505462 362543
rect 505496 362509 505552 362543
rect 505586 362509 505642 362543
rect 505676 362509 505732 362543
rect 505766 362509 505822 362543
rect 505856 362509 505972 362543
rect 504684 362476 505972 362509
rect 508444 373110 509732 373144
rect 508444 373076 508502 373110
rect 508536 373076 508592 373110
rect 508626 373076 508682 373110
rect 508716 373076 508772 373110
rect 508806 373076 508862 373110
rect 508896 373076 508952 373110
rect 508986 373076 509042 373110
rect 509076 373076 509132 373110
rect 509166 373076 509222 373110
rect 509256 373076 509312 373110
rect 509346 373076 509402 373110
rect 509436 373076 509492 373110
rect 509526 373076 509582 373110
rect 509616 373076 509732 373110
rect 508444 373043 509732 373076
rect 508444 373014 508545 373043
rect 508444 372980 508479 373014
rect 508513 372980 508545 373014
rect 509631 373014 509732 373043
rect 508444 372924 508545 372980
rect 508444 372890 508479 372924
rect 508513 372890 508545 372924
rect 508444 372834 508545 372890
rect 508444 372800 508479 372834
rect 508513 372800 508545 372834
rect 508444 372744 508545 372800
rect 508444 372710 508479 372744
rect 508513 372710 508545 372744
rect 508444 372654 508545 372710
rect 508444 372620 508479 372654
rect 508513 372620 508545 372654
rect 508444 372564 508545 372620
rect 508444 372530 508479 372564
rect 508513 372530 508545 372564
rect 508444 372474 508545 372530
rect 508444 372440 508479 372474
rect 508513 372440 508545 372474
rect 508444 372384 508545 372440
rect 508444 372350 508479 372384
rect 508513 372350 508545 372384
rect 508444 372294 508545 372350
rect 508444 372260 508479 372294
rect 508513 372260 508545 372294
rect 508444 372204 508545 372260
rect 508444 372170 508479 372204
rect 508513 372170 508545 372204
rect 508444 372114 508545 372170
rect 508444 372080 508479 372114
rect 508513 372080 508545 372114
rect 508444 372024 508545 372080
rect 508444 371990 508479 372024
rect 508513 371990 508545 372024
rect 509631 372980 509666 373014
rect 509700 372980 509732 373014
rect 509631 372924 509732 372980
rect 509631 372890 509666 372924
rect 509700 372890 509732 372924
rect 509631 372834 509732 372890
rect 509631 372800 509666 372834
rect 509700 372800 509732 372834
rect 509631 372744 509732 372800
rect 509631 372710 509666 372744
rect 509700 372710 509732 372744
rect 509631 372654 509732 372710
rect 509631 372620 509666 372654
rect 509700 372620 509732 372654
rect 509631 372564 509732 372620
rect 509631 372530 509666 372564
rect 509700 372530 509732 372564
rect 509631 372474 509732 372530
rect 509631 372440 509666 372474
rect 509700 372440 509732 372474
rect 509631 372384 509732 372440
rect 509631 372350 509666 372384
rect 509700 372350 509732 372384
rect 509631 372294 509732 372350
rect 509631 372260 509666 372294
rect 509700 372260 509732 372294
rect 509631 372204 509732 372260
rect 509631 372170 509666 372204
rect 509700 372170 509732 372204
rect 509631 372114 509732 372170
rect 509631 372080 509666 372114
rect 509700 372080 509732 372114
rect 509631 372024 509732 372080
rect 508444 371957 508545 371990
rect 509631 371990 509666 372024
rect 509700 371990 509732 372024
rect 509631 371957 509732 371990
rect 508444 371923 509732 371957
rect 508444 371889 508502 371923
rect 508536 371889 508592 371923
rect 508626 371889 508682 371923
rect 508716 371889 508772 371923
rect 508806 371889 508862 371923
rect 508896 371889 508952 371923
rect 508986 371889 509042 371923
rect 509076 371889 509132 371923
rect 509166 371889 509222 371923
rect 509256 371889 509312 371923
rect 509346 371889 509402 371923
rect 509436 371889 509492 371923
rect 509526 371889 509582 371923
rect 509616 371889 509732 371923
rect 508444 371770 509732 371889
rect 508444 371736 508502 371770
rect 508536 371736 508592 371770
rect 508626 371736 508682 371770
rect 508716 371736 508772 371770
rect 508806 371736 508862 371770
rect 508896 371736 508952 371770
rect 508986 371736 509042 371770
rect 509076 371736 509132 371770
rect 509166 371736 509222 371770
rect 509256 371736 509312 371770
rect 509346 371736 509402 371770
rect 509436 371736 509492 371770
rect 509526 371736 509582 371770
rect 509616 371736 509732 371770
rect 508444 371703 509732 371736
rect 508444 371674 508545 371703
rect 508444 371640 508479 371674
rect 508513 371640 508545 371674
rect 509631 371674 509732 371703
rect 508444 371584 508545 371640
rect 508444 371550 508479 371584
rect 508513 371550 508545 371584
rect 508444 371494 508545 371550
rect 508444 371460 508479 371494
rect 508513 371460 508545 371494
rect 508444 371404 508545 371460
rect 508444 371370 508479 371404
rect 508513 371370 508545 371404
rect 508444 371314 508545 371370
rect 508444 371280 508479 371314
rect 508513 371280 508545 371314
rect 508444 371224 508545 371280
rect 508444 371190 508479 371224
rect 508513 371190 508545 371224
rect 508444 371134 508545 371190
rect 508444 371100 508479 371134
rect 508513 371100 508545 371134
rect 508444 371044 508545 371100
rect 508444 371010 508479 371044
rect 508513 371010 508545 371044
rect 508444 370954 508545 371010
rect 508444 370920 508479 370954
rect 508513 370920 508545 370954
rect 508444 370864 508545 370920
rect 508444 370830 508479 370864
rect 508513 370830 508545 370864
rect 508444 370774 508545 370830
rect 508444 370740 508479 370774
rect 508513 370740 508545 370774
rect 508444 370684 508545 370740
rect 508444 370650 508479 370684
rect 508513 370650 508545 370684
rect 509631 371640 509666 371674
rect 509700 371640 509732 371674
rect 509631 371584 509732 371640
rect 509631 371550 509666 371584
rect 509700 371550 509732 371584
rect 509631 371494 509732 371550
rect 509631 371460 509666 371494
rect 509700 371460 509732 371494
rect 509631 371404 509732 371460
rect 509631 371370 509666 371404
rect 509700 371370 509732 371404
rect 509631 371314 509732 371370
rect 509631 371280 509666 371314
rect 509700 371280 509732 371314
rect 509631 371224 509732 371280
rect 509631 371190 509666 371224
rect 509700 371190 509732 371224
rect 509631 371134 509732 371190
rect 509631 371100 509666 371134
rect 509700 371100 509732 371134
rect 509631 371044 509732 371100
rect 509631 371010 509666 371044
rect 509700 371010 509732 371044
rect 509631 370954 509732 371010
rect 509631 370920 509666 370954
rect 509700 370920 509732 370954
rect 509631 370864 509732 370920
rect 509631 370830 509666 370864
rect 509700 370830 509732 370864
rect 509631 370774 509732 370830
rect 509631 370740 509666 370774
rect 509700 370740 509732 370774
rect 509631 370684 509732 370740
rect 508444 370617 508545 370650
rect 509631 370650 509666 370684
rect 509700 370650 509732 370684
rect 509631 370617 509732 370650
rect 508444 370583 509732 370617
rect 508444 370549 508502 370583
rect 508536 370549 508592 370583
rect 508626 370549 508682 370583
rect 508716 370549 508772 370583
rect 508806 370549 508862 370583
rect 508896 370549 508952 370583
rect 508986 370549 509042 370583
rect 509076 370549 509132 370583
rect 509166 370549 509222 370583
rect 509256 370549 509312 370583
rect 509346 370549 509402 370583
rect 509436 370549 509492 370583
rect 509526 370549 509582 370583
rect 509616 370549 509732 370583
rect 508444 370430 509732 370549
rect 508444 370396 508502 370430
rect 508536 370396 508592 370430
rect 508626 370396 508682 370430
rect 508716 370396 508772 370430
rect 508806 370396 508862 370430
rect 508896 370396 508952 370430
rect 508986 370396 509042 370430
rect 509076 370396 509132 370430
rect 509166 370396 509222 370430
rect 509256 370396 509312 370430
rect 509346 370396 509402 370430
rect 509436 370396 509492 370430
rect 509526 370396 509582 370430
rect 509616 370396 509732 370430
rect 508444 370363 509732 370396
rect 508444 370334 508545 370363
rect 508444 370300 508479 370334
rect 508513 370300 508545 370334
rect 509631 370334 509732 370363
rect 508444 370244 508545 370300
rect 508444 370210 508479 370244
rect 508513 370210 508545 370244
rect 508444 370154 508545 370210
rect 508444 370120 508479 370154
rect 508513 370120 508545 370154
rect 508444 370064 508545 370120
rect 508444 370030 508479 370064
rect 508513 370030 508545 370064
rect 508444 369974 508545 370030
rect 508444 369940 508479 369974
rect 508513 369940 508545 369974
rect 508444 369884 508545 369940
rect 508444 369850 508479 369884
rect 508513 369850 508545 369884
rect 508444 369794 508545 369850
rect 508444 369760 508479 369794
rect 508513 369760 508545 369794
rect 508444 369704 508545 369760
rect 508444 369670 508479 369704
rect 508513 369670 508545 369704
rect 508444 369614 508545 369670
rect 508444 369580 508479 369614
rect 508513 369580 508545 369614
rect 508444 369524 508545 369580
rect 508444 369490 508479 369524
rect 508513 369490 508545 369524
rect 508444 369434 508545 369490
rect 508444 369400 508479 369434
rect 508513 369400 508545 369434
rect 508444 369344 508545 369400
rect 508444 369310 508479 369344
rect 508513 369310 508545 369344
rect 509631 370300 509666 370334
rect 509700 370300 509732 370334
rect 509631 370244 509732 370300
rect 509631 370210 509666 370244
rect 509700 370210 509732 370244
rect 509631 370154 509732 370210
rect 509631 370120 509666 370154
rect 509700 370120 509732 370154
rect 509631 370064 509732 370120
rect 509631 370030 509666 370064
rect 509700 370030 509732 370064
rect 509631 369974 509732 370030
rect 509631 369940 509666 369974
rect 509700 369940 509732 369974
rect 509631 369884 509732 369940
rect 509631 369850 509666 369884
rect 509700 369850 509732 369884
rect 509631 369794 509732 369850
rect 509631 369760 509666 369794
rect 509700 369760 509732 369794
rect 509631 369704 509732 369760
rect 509631 369670 509666 369704
rect 509700 369670 509732 369704
rect 509631 369614 509732 369670
rect 509631 369580 509666 369614
rect 509700 369580 509732 369614
rect 509631 369524 509732 369580
rect 509631 369490 509666 369524
rect 509700 369490 509732 369524
rect 509631 369434 509732 369490
rect 509631 369400 509666 369434
rect 509700 369400 509732 369434
rect 509631 369344 509732 369400
rect 508444 369277 508545 369310
rect 509631 369310 509666 369344
rect 509700 369310 509732 369344
rect 509631 369277 509732 369310
rect 508444 369243 509732 369277
rect 508444 369209 508502 369243
rect 508536 369209 508592 369243
rect 508626 369209 508682 369243
rect 508716 369209 508772 369243
rect 508806 369209 508862 369243
rect 508896 369209 508952 369243
rect 508986 369209 509042 369243
rect 509076 369209 509132 369243
rect 509166 369209 509222 369243
rect 509256 369209 509312 369243
rect 509346 369209 509402 369243
rect 509436 369209 509492 369243
rect 509526 369209 509582 369243
rect 509616 369209 509732 369243
rect 508444 369090 509732 369209
rect 508444 369056 508502 369090
rect 508536 369056 508592 369090
rect 508626 369056 508682 369090
rect 508716 369056 508772 369090
rect 508806 369056 508862 369090
rect 508896 369056 508952 369090
rect 508986 369056 509042 369090
rect 509076 369056 509132 369090
rect 509166 369056 509222 369090
rect 509256 369056 509312 369090
rect 509346 369056 509402 369090
rect 509436 369056 509492 369090
rect 509526 369056 509582 369090
rect 509616 369056 509732 369090
rect 508444 369023 509732 369056
rect 508444 368994 508545 369023
rect 508444 368960 508479 368994
rect 508513 368960 508545 368994
rect 509631 368994 509732 369023
rect 508444 368904 508545 368960
rect 508444 368870 508479 368904
rect 508513 368870 508545 368904
rect 508444 368814 508545 368870
rect 508444 368780 508479 368814
rect 508513 368780 508545 368814
rect 508444 368724 508545 368780
rect 508444 368690 508479 368724
rect 508513 368690 508545 368724
rect 508444 368634 508545 368690
rect 508444 368600 508479 368634
rect 508513 368600 508545 368634
rect 508444 368544 508545 368600
rect 508444 368510 508479 368544
rect 508513 368510 508545 368544
rect 508444 368454 508545 368510
rect 508444 368420 508479 368454
rect 508513 368420 508545 368454
rect 508444 368364 508545 368420
rect 508444 368330 508479 368364
rect 508513 368330 508545 368364
rect 508444 368274 508545 368330
rect 508444 368240 508479 368274
rect 508513 368240 508545 368274
rect 508444 368184 508545 368240
rect 508444 368150 508479 368184
rect 508513 368150 508545 368184
rect 508444 368094 508545 368150
rect 508444 368060 508479 368094
rect 508513 368060 508545 368094
rect 508444 368004 508545 368060
rect 508444 367970 508479 368004
rect 508513 367970 508545 368004
rect 509631 368960 509666 368994
rect 509700 368960 509732 368994
rect 509631 368904 509732 368960
rect 509631 368870 509666 368904
rect 509700 368870 509732 368904
rect 509631 368814 509732 368870
rect 509631 368780 509666 368814
rect 509700 368780 509732 368814
rect 509631 368724 509732 368780
rect 509631 368690 509666 368724
rect 509700 368690 509732 368724
rect 509631 368634 509732 368690
rect 509631 368600 509666 368634
rect 509700 368600 509732 368634
rect 509631 368544 509732 368600
rect 509631 368510 509666 368544
rect 509700 368510 509732 368544
rect 509631 368454 509732 368510
rect 509631 368420 509666 368454
rect 509700 368420 509732 368454
rect 509631 368364 509732 368420
rect 509631 368330 509666 368364
rect 509700 368330 509732 368364
rect 509631 368274 509732 368330
rect 509631 368240 509666 368274
rect 509700 368240 509732 368274
rect 509631 368184 509732 368240
rect 509631 368150 509666 368184
rect 509700 368150 509732 368184
rect 509631 368094 509732 368150
rect 509631 368060 509666 368094
rect 509700 368060 509732 368094
rect 509631 368004 509732 368060
rect 508444 367937 508545 367970
rect 509631 367970 509666 368004
rect 509700 367970 509732 368004
rect 509631 367937 509732 367970
rect 508444 367903 509732 367937
rect 508444 367869 508502 367903
rect 508536 367869 508592 367903
rect 508626 367869 508682 367903
rect 508716 367869 508772 367903
rect 508806 367869 508862 367903
rect 508896 367869 508952 367903
rect 508986 367869 509042 367903
rect 509076 367869 509132 367903
rect 509166 367869 509222 367903
rect 509256 367869 509312 367903
rect 509346 367869 509402 367903
rect 509436 367869 509492 367903
rect 509526 367869 509582 367903
rect 509616 367869 509732 367903
rect 508444 367750 509732 367869
rect 508444 367716 508502 367750
rect 508536 367716 508592 367750
rect 508626 367716 508682 367750
rect 508716 367716 508772 367750
rect 508806 367716 508862 367750
rect 508896 367716 508952 367750
rect 508986 367716 509042 367750
rect 509076 367716 509132 367750
rect 509166 367716 509222 367750
rect 509256 367716 509312 367750
rect 509346 367716 509402 367750
rect 509436 367716 509492 367750
rect 509526 367716 509582 367750
rect 509616 367716 509732 367750
rect 508444 367683 509732 367716
rect 508444 367654 508545 367683
rect 508444 367620 508479 367654
rect 508513 367620 508545 367654
rect 509631 367654 509732 367683
rect 508444 367564 508545 367620
rect 508444 367530 508479 367564
rect 508513 367530 508545 367564
rect 508444 367474 508545 367530
rect 508444 367440 508479 367474
rect 508513 367440 508545 367474
rect 508444 367384 508545 367440
rect 508444 367350 508479 367384
rect 508513 367350 508545 367384
rect 508444 367294 508545 367350
rect 508444 367260 508479 367294
rect 508513 367260 508545 367294
rect 508444 367204 508545 367260
rect 508444 367170 508479 367204
rect 508513 367170 508545 367204
rect 508444 367114 508545 367170
rect 508444 367080 508479 367114
rect 508513 367080 508545 367114
rect 508444 367024 508545 367080
rect 508444 366990 508479 367024
rect 508513 366990 508545 367024
rect 508444 366934 508545 366990
rect 508444 366900 508479 366934
rect 508513 366900 508545 366934
rect 508444 366844 508545 366900
rect 508444 366810 508479 366844
rect 508513 366810 508545 366844
rect 508444 366754 508545 366810
rect 508444 366720 508479 366754
rect 508513 366720 508545 366754
rect 508444 366664 508545 366720
rect 508444 366630 508479 366664
rect 508513 366630 508545 366664
rect 509631 367620 509666 367654
rect 509700 367620 509732 367654
rect 509631 367564 509732 367620
rect 509631 367530 509666 367564
rect 509700 367530 509732 367564
rect 509631 367474 509732 367530
rect 509631 367440 509666 367474
rect 509700 367440 509732 367474
rect 509631 367384 509732 367440
rect 509631 367350 509666 367384
rect 509700 367350 509732 367384
rect 509631 367294 509732 367350
rect 509631 367260 509666 367294
rect 509700 367260 509732 367294
rect 509631 367204 509732 367260
rect 509631 367170 509666 367204
rect 509700 367170 509732 367204
rect 509631 367114 509732 367170
rect 509631 367080 509666 367114
rect 509700 367080 509732 367114
rect 509631 367024 509732 367080
rect 509631 366990 509666 367024
rect 509700 366990 509732 367024
rect 509631 366934 509732 366990
rect 509631 366900 509666 366934
rect 509700 366900 509732 366934
rect 509631 366844 509732 366900
rect 509631 366810 509666 366844
rect 509700 366810 509732 366844
rect 509631 366754 509732 366810
rect 509631 366720 509666 366754
rect 509700 366720 509732 366754
rect 509631 366664 509732 366720
rect 508444 366597 508545 366630
rect 509631 366630 509666 366664
rect 509700 366630 509732 366664
rect 509631 366597 509732 366630
rect 508444 366563 509732 366597
rect 508444 366529 508502 366563
rect 508536 366529 508592 366563
rect 508626 366529 508682 366563
rect 508716 366529 508772 366563
rect 508806 366529 508862 366563
rect 508896 366529 508952 366563
rect 508986 366529 509042 366563
rect 509076 366529 509132 366563
rect 509166 366529 509222 366563
rect 509256 366529 509312 366563
rect 509346 366529 509402 366563
rect 509436 366529 509492 366563
rect 509526 366529 509582 366563
rect 509616 366529 509732 366563
rect 508444 366410 509732 366529
rect 508444 366376 508502 366410
rect 508536 366376 508592 366410
rect 508626 366376 508682 366410
rect 508716 366376 508772 366410
rect 508806 366376 508862 366410
rect 508896 366376 508952 366410
rect 508986 366376 509042 366410
rect 509076 366376 509132 366410
rect 509166 366376 509222 366410
rect 509256 366376 509312 366410
rect 509346 366376 509402 366410
rect 509436 366376 509492 366410
rect 509526 366376 509582 366410
rect 509616 366376 509732 366410
rect 508444 366343 509732 366376
rect 508444 366314 508545 366343
rect 508444 366280 508479 366314
rect 508513 366280 508545 366314
rect 509631 366314 509732 366343
rect 508444 366224 508545 366280
rect 508444 366190 508479 366224
rect 508513 366190 508545 366224
rect 508444 366134 508545 366190
rect 508444 366100 508479 366134
rect 508513 366100 508545 366134
rect 508444 366044 508545 366100
rect 508444 366010 508479 366044
rect 508513 366010 508545 366044
rect 508444 365954 508545 366010
rect 508444 365920 508479 365954
rect 508513 365920 508545 365954
rect 508444 365864 508545 365920
rect 508444 365830 508479 365864
rect 508513 365830 508545 365864
rect 508444 365774 508545 365830
rect 508444 365740 508479 365774
rect 508513 365740 508545 365774
rect 508444 365684 508545 365740
rect 508444 365650 508479 365684
rect 508513 365650 508545 365684
rect 508444 365594 508545 365650
rect 508444 365560 508479 365594
rect 508513 365560 508545 365594
rect 508444 365504 508545 365560
rect 508444 365470 508479 365504
rect 508513 365470 508545 365504
rect 508444 365414 508545 365470
rect 508444 365380 508479 365414
rect 508513 365380 508545 365414
rect 508444 365324 508545 365380
rect 508444 365290 508479 365324
rect 508513 365290 508545 365324
rect 509631 366280 509666 366314
rect 509700 366280 509732 366314
rect 509631 366224 509732 366280
rect 509631 366190 509666 366224
rect 509700 366190 509732 366224
rect 509631 366134 509732 366190
rect 509631 366100 509666 366134
rect 509700 366100 509732 366134
rect 509631 366044 509732 366100
rect 509631 366010 509666 366044
rect 509700 366010 509732 366044
rect 509631 365954 509732 366010
rect 509631 365920 509666 365954
rect 509700 365920 509732 365954
rect 509631 365864 509732 365920
rect 509631 365830 509666 365864
rect 509700 365830 509732 365864
rect 509631 365774 509732 365830
rect 509631 365740 509666 365774
rect 509700 365740 509732 365774
rect 509631 365684 509732 365740
rect 509631 365650 509666 365684
rect 509700 365650 509732 365684
rect 509631 365594 509732 365650
rect 509631 365560 509666 365594
rect 509700 365560 509732 365594
rect 509631 365504 509732 365560
rect 509631 365470 509666 365504
rect 509700 365470 509732 365504
rect 509631 365414 509732 365470
rect 509631 365380 509666 365414
rect 509700 365380 509732 365414
rect 509631 365324 509732 365380
rect 508444 365257 508545 365290
rect 509631 365290 509666 365324
rect 509700 365290 509732 365324
rect 509631 365257 509732 365290
rect 508444 365223 509732 365257
rect 508444 365189 508502 365223
rect 508536 365189 508592 365223
rect 508626 365189 508682 365223
rect 508716 365189 508772 365223
rect 508806 365189 508862 365223
rect 508896 365189 508952 365223
rect 508986 365189 509042 365223
rect 509076 365189 509132 365223
rect 509166 365189 509222 365223
rect 509256 365189 509312 365223
rect 509346 365189 509402 365223
rect 509436 365189 509492 365223
rect 509526 365189 509582 365223
rect 509616 365189 509732 365223
rect 508444 365070 509732 365189
rect 508444 365036 508502 365070
rect 508536 365036 508592 365070
rect 508626 365036 508682 365070
rect 508716 365036 508772 365070
rect 508806 365036 508862 365070
rect 508896 365036 508952 365070
rect 508986 365036 509042 365070
rect 509076 365036 509132 365070
rect 509166 365036 509222 365070
rect 509256 365036 509312 365070
rect 509346 365036 509402 365070
rect 509436 365036 509492 365070
rect 509526 365036 509582 365070
rect 509616 365036 509732 365070
rect 508444 365003 509732 365036
rect 508444 364974 508545 365003
rect 508444 364940 508479 364974
rect 508513 364940 508545 364974
rect 509631 364974 509732 365003
rect 508444 364884 508545 364940
rect 508444 364850 508479 364884
rect 508513 364850 508545 364884
rect 508444 364794 508545 364850
rect 508444 364760 508479 364794
rect 508513 364760 508545 364794
rect 508444 364704 508545 364760
rect 508444 364670 508479 364704
rect 508513 364670 508545 364704
rect 508444 364614 508545 364670
rect 508444 364580 508479 364614
rect 508513 364580 508545 364614
rect 508444 364524 508545 364580
rect 508444 364490 508479 364524
rect 508513 364490 508545 364524
rect 508444 364434 508545 364490
rect 508444 364400 508479 364434
rect 508513 364400 508545 364434
rect 508444 364344 508545 364400
rect 508444 364310 508479 364344
rect 508513 364310 508545 364344
rect 508444 364254 508545 364310
rect 508444 364220 508479 364254
rect 508513 364220 508545 364254
rect 508444 364164 508545 364220
rect 508444 364130 508479 364164
rect 508513 364130 508545 364164
rect 508444 364074 508545 364130
rect 508444 364040 508479 364074
rect 508513 364040 508545 364074
rect 508444 363984 508545 364040
rect 508444 363950 508479 363984
rect 508513 363950 508545 363984
rect 509631 364940 509666 364974
rect 509700 364940 509732 364974
rect 509631 364884 509732 364940
rect 509631 364850 509666 364884
rect 509700 364850 509732 364884
rect 509631 364794 509732 364850
rect 509631 364760 509666 364794
rect 509700 364760 509732 364794
rect 509631 364704 509732 364760
rect 509631 364670 509666 364704
rect 509700 364670 509732 364704
rect 509631 364614 509732 364670
rect 509631 364580 509666 364614
rect 509700 364580 509732 364614
rect 509631 364524 509732 364580
rect 509631 364490 509666 364524
rect 509700 364490 509732 364524
rect 509631 364434 509732 364490
rect 509631 364400 509666 364434
rect 509700 364400 509732 364434
rect 509631 364344 509732 364400
rect 509631 364310 509666 364344
rect 509700 364310 509732 364344
rect 509631 364254 509732 364310
rect 509631 364220 509666 364254
rect 509700 364220 509732 364254
rect 509631 364164 509732 364220
rect 509631 364130 509666 364164
rect 509700 364130 509732 364164
rect 509631 364074 509732 364130
rect 509631 364040 509666 364074
rect 509700 364040 509732 364074
rect 509631 363984 509732 364040
rect 508444 363917 508545 363950
rect 509631 363950 509666 363984
rect 509700 363950 509732 363984
rect 509631 363917 509732 363950
rect 508444 363883 509732 363917
rect 508444 363849 508502 363883
rect 508536 363849 508592 363883
rect 508626 363849 508682 363883
rect 508716 363849 508772 363883
rect 508806 363849 508862 363883
rect 508896 363849 508952 363883
rect 508986 363849 509042 363883
rect 509076 363849 509132 363883
rect 509166 363849 509222 363883
rect 509256 363849 509312 363883
rect 509346 363849 509402 363883
rect 509436 363849 509492 363883
rect 509526 363849 509582 363883
rect 509616 363849 509732 363883
rect 508444 363730 509732 363849
rect 508444 363696 508502 363730
rect 508536 363696 508592 363730
rect 508626 363696 508682 363730
rect 508716 363696 508772 363730
rect 508806 363696 508862 363730
rect 508896 363696 508952 363730
rect 508986 363696 509042 363730
rect 509076 363696 509132 363730
rect 509166 363696 509222 363730
rect 509256 363696 509312 363730
rect 509346 363696 509402 363730
rect 509436 363696 509492 363730
rect 509526 363696 509582 363730
rect 509616 363696 509732 363730
rect 508444 363663 509732 363696
rect 508444 363634 508545 363663
rect 508444 363600 508479 363634
rect 508513 363600 508545 363634
rect 509631 363634 509732 363663
rect 508444 363544 508545 363600
rect 508444 363510 508479 363544
rect 508513 363510 508545 363544
rect 508444 363454 508545 363510
rect 508444 363420 508479 363454
rect 508513 363420 508545 363454
rect 508444 363364 508545 363420
rect 508444 363330 508479 363364
rect 508513 363330 508545 363364
rect 508444 363274 508545 363330
rect 508444 363240 508479 363274
rect 508513 363240 508545 363274
rect 508444 363184 508545 363240
rect 508444 363150 508479 363184
rect 508513 363150 508545 363184
rect 508444 363094 508545 363150
rect 508444 363060 508479 363094
rect 508513 363060 508545 363094
rect 508444 363004 508545 363060
rect 508444 362970 508479 363004
rect 508513 362970 508545 363004
rect 508444 362914 508545 362970
rect 508444 362880 508479 362914
rect 508513 362880 508545 362914
rect 508444 362824 508545 362880
rect 508444 362790 508479 362824
rect 508513 362790 508545 362824
rect 508444 362734 508545 362790
rect 508444 362700 508479 362734
rect 508513 362700 508545 362734
rect 508444 362644 508545 362700
rect 508444 362610 508479 362644
rect 508513 362610 508545 362644
rect 509631 363600 509666 363634
rect 509700 363600 509732 363634
rect 509631 363544 509732 363600
rect 509631 363510 509666 363544
rect 509700 363510 509732 363544
rect 509631 363454 509732 363510
rect 509631 363420 509666 363454
rect 509700 363420 509732 363454
rect 509631 363364 509732 363420
rect 509631 363330 509666 363364
rect 509700 363330 509732 363364
rect 509631 363274 509732 363330
rect 509631 363240 509666 363274
rect 509700 363240 509732 363274
rect 509631 363184 509732 363240
rect 509631 363150 509666 363184
rect 509700 363150 509732 363184
rect 509631 363094 509732 363150
rect 509631 363060 509666 363094
rect 509700 363060 509732 363094
rect 509631 363004 509732 363060
rect 509631 362970 509666 363004
rect 509700 362970 509732 363004
rect 509631 362914 509732 362970
rect 509631 362880 509666 362914
rect 509700 362880 509732 362914
rect 509631 362824 509732 362880
rect 509631 362790 509666 362824
rect 509700 362790 509732 362824
rect 509631 362734 509732 362790
rect 509631 362700 509666 362734
rect 509700 362700 509732 362734
rect 509631 362644 509732 362700
rect 508444 362577 508545 362610
rect 509631 362610 509666 362644
rect 509700 362610 509732 362644
rect 509631 362577 509732 362610
rect 508444 362543 509732 362577
rect 508444 362509 508502 362543
rect 508536 362509 508592 362543
rect 508626 362509 508682 362543
rect 508716 362509 508772 362543
rect 508806 362509 508862 362543
rect 508896 362509 508952 362543
rect 508986 362509 509042 362543
rect 509076 362509 509132 362543
rect 509166 362509 509222 362543
rect 509256 362509 509312 362543
rect 509346 362509 509402 362543
rect 509436 362509 509492 362543
rect 509526 362509 509582 362543
rect 509616 362509 509732 362543
rect 508444 362476 509732 362509
rect 512204 373110 513492 373144
rect 512204 373076 512262 373110
rect 512296 373076 512352 373110
rect 512386 373076 512442 373110
rect 512476 373076 512532 373110
rect 512566 373076 512622 373110
rect 512656 373076 512712 373110
rect 512746 373076 512802 373110
rect 512836 373076 512892 373110
rect 512926 373076 512982 373110
rect 513016 373076 513072 373110
rect 513106 373076 513162 373110
rect 513196 373076 513252 373110
rect 513286 373076 513342 373110
rect 513376 373076 513492 373110
rect 512204 373043 513492 373076
rect 512204 373014 512305 373043
rect 512204 372980 512239 373014
rect 512273 372980 512305 373014
rect 513391 373014 513492 373043
rect 512204 372924 512305 372980
rect 512204 372890 512239 372924
rect 512273 372890 512305 372924
rect 512204 372834 512305 372890
rect 512204 372800 512239 372834
rect 512273 372800 512305 372834
rect 512204 372744 512305 372800
rect 512204 372710 512239 372744
rect 512273 372710 512305 372744
rect 512204 372654 512305 372710
rect 512204 372620 512239 372654
rect 512273 372620 512305 372654
rect 512204 372564 512305 372620
rect 512204 372530 512239 372564
rect 512273 372530 512305 372564
rect 512204 372474 512305 372530
rect 512204 372440 512239 372474
rect 512273 372440 512305 372474
rect 512204 372384 512305 372440
rect 512204 372350 512239 372384
rect 512273 372350 512305 372384
rect 512204 372294 512305 372350
rect 512204 372260 512239 372294
rect 512273 372260 512305 372294
rect 512204 372204 512305 372260
rect 512204 372170 512239 372204
rect 512273 372170 512305 372204
rect 512204 372114 512305 372170
rect 512204 372080 512239 372114
rect 512273 372080 512305 372114
rect 512204 372024 512305 372080
rect 512204 371990 512239 372024
rect 512273 371990 512305 372024
rect 513391 372980 513426 373014
rect 513460 372980 513492 373014
rect 513391 372924 513492 372980
rect 513391 372890 513426 372924
rect 513460 372890 513492 372924
rect 513391 372834 513492 372890
rect 513391 372800 513426 372834
rect 513460 372800 513492 372834
rect 513391 372744 513492 372800
rect 513391 372710 513426 372744
rect 513460 372710 513492 372744
rect 513391 372654 513492 372710
rect 513391 372620 513426 372654
rect 513460 372620 513492 372654
rect 513391 372564 513492 372620
rect 513391 372530 513426 372564
rect 513460 372530 513492 372564
rect 513391 372474 513492 372530
rect 513391 372440 513426 372474
rect 513460 372440 513492 372474
rect 513391 372384 513492 372440
rect 513391 372350 513426 372384
rect 513460 372350 513492 372384
rect 516578 373817 516758 373904
rect 516578 373375 516617 373817
rect 516719 373375 516758 373817
rect 516578 373288 516758 373375
rect 520338 373817 520518 373904
rect 520338 373375 520377 373817
rect 520479 373375 520518 373817
rect 520338 373288 520518 373375
rect 513391 372294 513492 372350
rect 513391 372260 513426 372294
rect 513460 372260 513492 372294
rect 513391 372204 513492 372260
rect 513391 372170 513426 372204
rect 513460 372170 513492 372204
rect 513391 372114 513492 372170
rect 513391 372080 513426 372114
rect 513460 372080 513492 372114
rect 513391 372024 513492 372080
rect 512204 371957 512305 371990
rect 513391 371990 513426 372024
rect 513460 371990 513492 372024
rect 513391 371957 513492 371990
rect 512204 371923 513492 371957
rect 512204 371889 512262 371923
rect 512296 371889 512352 371923
rect 512386 371889 512442 371923
rect 512476 371889 512532 371923
rect 512566 371889 512622 371923
rect 512656 371889 512712 371923
rect 512746 371889 512802 371923
rect 512836 371889 512892 371923
rect 512926 371889 512982 371923
rect 513016 371889 513072 371923
rect 513106 371889 513162 371923
rect 513196 371889 513252 371923
rect 513286 371889 513342 371923
rect 513376 371889 513492 371923
rect 512204 371770 513492 371889
rect 512204 371736 512262 371770
rect 512296 371736 512352 371770
rect 512386 371736 512442 371770
rect 512476 371736 512532 371770
rect 512566 371736 512622 371770
rect 512656 371736 512712 371770
rect 512746 371736 512802 371770
rect 512836 371736 512892 371770
rect 512926 371736 512982 371770
rect 513016 371736 513072 371770
rect 513106 371736 513162 371770
rect 513196 371736 513252 371770
rect 513286 371736 513342 371770
rect 513376 371736 513492 371770
rect 512204 371703 513492 371736
rect 512204 371674 512305 371703
rect 512204 371640 512239 371674
rect 512273 371640 512305 371674
rect 513391 371674 513492 371703
rect 512204 371584 512305 371640
rect 512204 371550 512239 371584
rect 512273 371550 512305 371584
rect 512204 371494 512305 371550
rect 512204 371460 512239 371494
rect 512273 371460 512305 371494
rect 512204 371404 512305 371460
rect 512204 371370 512239 371404
rect 512273 371370 512305 371404
rect 512204 371314 512305 371370
rect 512204 371280 512239 371314
rect 512273 371280 512305 371314
rect 512204 371224 512305 371280
rect 512204 371190 512239 371224
rect 512273 371190 512305 371224
rect 512204 371134 512305 371190
rect 512204 371100 512239 371134
rect 512273 371100 512305 371134
rect 512204 371044 512305 371100
rect 512204 371010 512239 371044
rect 512273 371010 512305 371044
rect 512204 370954 512305 371010
rect 512204 370920 512239 370954
rect 512273 370920 512305 370954
rect 512204 370864 512305 370920
rect 512204 370830 512239 370864
rect 512273 370830 512305 370864
rect 512204 370774 512305 370830
rect 512204 370740 512239 370774
rect 512273 370740 512305 370774
rect 512204 370684 512305 370740
rect 512204 370650 512239 370684
rect 512273 370650 512305 370684
rect 513391 371640 513426 371674
rect 513460 371640 513492 371674
rect 513391 371584 513492 371640
rect 513391 371550 513426 371584
rect 513460 371550 513492 371584
rect 513391 371494 513492 371550
rect 513391 371460 513426 371494
rect 513460 371460 513492 371494
rect 513391 371404 513492 371460
rect 513391 371370 513426 371404
rect 513460 371370 513492 371404
rect 513391 371314 513492 371370
rect 513391 371280 513426 371314
rect 513460 371280 513492 371314
rect 513391 371224 513492 371280
rect 513391 371190 513426 371224
rect 513460 371190 513492 371224
rect 513391 371134 513492 371190
rect 513391 371100 513426 371134
rect 513460 371100 513492 371134
rect 513391 371044 513492 371100
rect 513391 371010 513426 371044
rect 513460 371010 513492 371044
rect 513391 370954 513492 371010
rect 513391 370920 513426 370954
rect 513460 370920 513492 370954
rect 513391 370864 513492 370920
rect 513391 370830 513426 370864
rect 513460 370830 513492 370864
rect 513391 370774 513492 370830
rect 513391 370740 513426 370774
rect 513460 370740 513492 370774
rect 513391 370684 513492 370740
rect 512204 370617 512305 370650
rect 513391 370650 513426 370684
rect 513460 370650 513492 370684
rect 513391 370617 513492 370650
rect 512204 370583 513492 370617
rect 512204 370549 512262 370583
rect 512296 370549 512352 370583
rect 512386 370549 512442 370583
rect 512476 370549 512532 370583
rect 512566 370549 512622 370583
rect 512656 370549 512712 370583
rect 512746 370549 512802 370583
rect 512836 370549 512892 370583
rect 512926 370549 512982 370583
rect 513016 370549 513072 370583
rect 513106 370549 513162 370583
rect 513196 370549 513252 370583
rect 513286 370549 513342 370583
rect 513376 370549 513492 370583
rect 512204 370430 513492 370549
rect 512204 370396 512262 370430
rect 512296 370396 512352 370430
rect 512386 370396 512442 370430
rect 512476 370396 512532 370430
rect 512566 370396 512622 370430
rect 512656 370396 512712 370430
rect 512746 370396 512802 370430
rect 512836 370396 512892 370430
rect 512926 370396 512982 370430
rect 513016 370396 513072 370430
rect 513106 370396 513162 370430
rect 513196 370396 513252 370430
rect 513286 370396 513342 370430
rect 513376 370396 513492 370430
rect 512204 370363 513492 370396
rect 512204 370334 512305 370363
rect 512204 370300 512239 370334
rect 512273 370300 512305 370334
rect 513391 370334 513492 370363
rect 512204 370244 512305 370300
rect 512204 370210 512239 370244
rect 512273 370210 512305 370244
rect 512204 370154 512305 370210
rect 512204 370120 512239 370154
rect 512273 370120 512305 370154
rect 512204 370064 512305 370120
rect 512204 370030 512239 370064
rect 512273 370030 512305 370064
rect 512204 369974 512305 370030
rect 512204 369940 512239 369974
rect 512273 369940 512305 369974
rect 512204 369884 512305 369940
rect 512204 369850 512239 369884
rect 512273 369850 512305 369884
rect 512204 369794 512305 369850
rect 512204 369760 512239 369794
rect 512273 369760 512305 369794
rect 512204 369704 512305 369760
rect 512204 369670 512239 369704
rect 512273 369670 512305 369704
rect 512204 369614 512305 369670
rect 512204 369580 512239 369614
rect 512273 369580 512305 369614
rect 512204 369524 512305 369580
rect 512204 369490 512239 369524
rect 512273 369490 512305 369524
rect 512204 369434 512305 369490
rect 512204 369400 512239 369434
rect 512273 369400 512305 369434
rect 512204 369344 512305 369400
rect 512204 369310 512239 369344
rect 512273 369310 512305 369344
rect 513391 370300 513426 370334
rect 513460 370300 513492 370334
rect 513391 370244 513492 370300
rect 513391 370210 513426 370244
rect 513460 370210 513492 370244
rect 513391 370154 513492 370210
rect 513391 370120 513426 370154
rect 513460 370120 513492 370154
rect 513391 370064 513492 370120
rect 513391 370030 513426 370064
rect 513460 370030 513492 370064
rect 513391 369974 513492 370030
rect 513391 369940 513426 369974
rect 513460 369940 513492 369974
rect 513391 369884 513492 369940
rect 513391 369850 513426 369884
rect 513460 369850 513492 369884
rect 513391 369794 513492 369850
rect 513391 369760 513426 369794
rect 513460 369760 513492 369794
rect 513391 369704 513492 369760
rect 513391 369670 513426 369704
rect 513460 369670 513492 369704
rect 513391 369614 513492 369670
rect 516578 371073 516758 371160
rect 516578 370631 516617 371073
rect 516719 370631 516758 371073
rect 516578 370544 516758 370631
rect 513391 369580 513426 369614
rect 513460 369580 513492 369614
rect 513391 369524 513492 369580
rect 513391 369490 513426 369524
rect 513460 369490 513492 369524
rect 513391 369434 513492 369490
rect 513391 369400 513426 369434
rect 513460 369400 513492 369434
rect 513391 369344 513492 369400
rect 512204 369277 512305 369310
rect 513391 369310 513426 369344
rect 513460 369310 513492 369344
rect 513391 369277 513492 369310
rect 512204 369243 513492 369277
rect 512204 369209 512262 369243
rect 512296 369209 512352 369243
rect 512386 369209 512442 369243
rect 512476 369209 512532 369243
rect 512566 369209 512622 369243
rect 512656 369209 512712 369243
rect 512746 369209 512802 369243
rect 512836 369209 512892 369243
rect 512926 369209 512982 369243
rect 513016 369209 513072 369243
rect 513106 369209 513162 369243
rect 513196 369209 513252 369243
rect 513286 369209 513342 369243
rect 513376 369209 513492 369243
rect 512204 369090 513492 369209
rect 512204 369056 512262 369090
rect 512296 369056 512352 369090
rect 512386 369056 512442 369090
rect 512476 369056 512532 369090
rect 512566 369056 512622 369090
rect 512656 369056 512712 369090
rect 512746 369056 512802 369090
rect 512836 369056 512892 369090
rect 512926 369056 512982 369090
rect 513016 369056 513072 369090
rect 513106 369056 513162 369090
rect 513196 369056 513252 369090
rect 513286 369056 513342 369090
rect 513376 369056 513492 369090
rect 512204 369023 513492 369056
rect 512204 368994 512305 369023
rect 512204 368960 512239 368994
rect 512273 368960 512305 368994
rect 513391 368994 513492 369023
rect 512204 368904 512305 368960
rect 512204 368870 512239 368904
rect 512273 368870 512305 368904
rect 512204 368814 512305 368870
rect 512204 368780 512239 368814
rect 512273 368780 512305 368814
rect 512204 368724 512305 368780
rect 512204 368690 512239 368724
rect 512273 368690 512305 368724
rect 512204 368634 512305 368690
rect 512204 368600 512239 368634
rect 512273 368600 512305 368634
rect 512204 368544 512305 368600
rect 512204 368510 512239 368544
rect 512273 368510 512305 368544
rect 512204 368454 512305 368510
rect 512204 368420 512239 368454
rect 512273 368420 512305 368454
rect 512204 368364 512305 368420
rect 512204 368330 512239 368364
rect 512273 368330 512305 368364
rect 512204 368274 512305 368330
rect 512204 368240 512239 368274
rect 512273 368240 512305 368274
rect 512204 368184 512305 368240
rect 512204 368150 512239 368184
rect 512273 368150 512305 368184
rect 512204 368094 512305 368150
rect 512204 368060 512239 368094
rect 512273 368060 512305 368094
rect 512204 368004 512305 368060
rect 512204 367970 512239 368004
rect 512273 367970 512305 368004
rect 513391 368960 513426 368994
rect 513460 368960 513492 368994
rect 513391 368904 513492 368960
rect 513391 368870 513426 368904
rect 513460 368870 513492 368904
rect 513391 368814 513492 368870
rect 513391 368780 513426 368814
rect 513460 368780 513492 368814
rect 513391 368724 513492 368780
rect 513391 368690 513426 368724
rect 513460 368690 513492 368724
rect 513391 368634 513492 368690
rect 513391 368600 513426 368634
rect 513460 368600 513492 368634
rect 513391 368544 513492 368600
rect 513391 368510 513426 368544
rect 513460 368510 513492 368544
rect 513391 368454 513492 368510
rect 513391 368420 513426 368454
rect 513460 368420 513492 368454
rect 513391 368364 513492 368420
rect 513391 368330 513426 368364
rect 513460 368330 513492 368364
rect 513391 368274 513492 368330
rect 513391 368240 513426 368274
rect 513460 368240 513492 368274
rect 513391 368184 513492 368240
rect 513391 368150 513426 368184
rect 513460 368150 513492 368184
rect 513391 368094 513492 368150
rect 513391 368060 513426 368094
rect 513460 368060 513492 368094
rect 513391 368004 513492 368060
rect 512204 367937 512305 367970
rect 513391 367970 513426 368004
rect 513460 367970 513492 368004
rect 513391 367937 513492 367970
rect 512204 367903 513492 367937
rect 512204 367869 512262 367903
rect 512296 367869 512352 367903
rect 512386 367869 512442 367903
rect 512476 367869 512532 367903
rect 512566 367869 512622 367903
rect 512656 367869 512712 367903
rect 512746 367869 512802 367903
rect 512836 367869 512892 367903
rect 512926 367869 512982 367903
rect 513016 367869 513072 367903
rect 513106 367869 513162 367903
rect 513196 367869 513252 367903
rect 513286 367869 513342 367903
rect 513376 367869 513492 367903
rect 512204 367750 513492 367869
rect 512204 367716 512262 367750
rect 512296 367716 512352 367750
rect 512386 367716 512442 367750
rect 512476 367716 512532 367750
rect 512566 367716 512622 367750
rect 512656 367716 512712 367750
rect 512746 367716 512802 367750
rect 512836 367716 512892 367750
rect 512926 367716 512982 367750
rect 513016 367716 513072 367750
rect 513106 367716 513162 367750
rect 513196 367716 513252 367750
rect 513286 367716 513342 367750
rect 513376 367716 513492 367750
rect 512204 367683 513492 367716
rect 512204 367654 512305 367683
rect 512204 367620 512239 367654
rect 512273 367620 512305 367654
rect 513391 367654 513492 367683
rect 512204 367564 512305 367620
rect 512204 367530 512239 367564
rect 512273 367530 512305 367564
rect 512204 367474 512305 367530
rect 512204 367440 512239 367474
rect 512273 367440 512305 367474
rect 512204 367384 512305 367440
rect 512204 367350 512239 367384
rect 512273 367350 512305 367384
rect 512204 367294 512305 367350
rect 512204 367260 512239 367294
rect 512273 367260 512305 367294
rect 512204 367204 512305 367260
rect 512204 367170 512239 367204
rect 512273 367170 512305 367204
rect 512204 367114 512305 367170
rect 512204 367080 512239 367114
rect 512273 367080 512305 367114
rect 512204 367024 512305 367080
rect 512204 366990 512239 367024
rect 512273 366990 512305 367024
rect 512204 366934 512305 366990
rect 512204 366900 512239 366934
rect 512273 366900 512305 366934
rect 512204 366844 512305 366900
rect 512204 366810 512239 366844
rect 512273 366810 512305 366844
rect 512204 366754 512305 366810
rect 512204 366720 512239 366754
rect 512273 366720 512305 366754
rect 512204 366664 512305 366720
rect 512204 366630 512239 366664
rect 512273 366630 512305 366664
rect 513391 367620 513426 367654
rect 513460 367620 513492 367654
rect 513391 367564 513492 367620
rect 513391 367530 513426 367564
rect 513460 367530 513492 367564
rect 513391 367474 513492 367530
rect 513391 367440 513426 367474
rect 513460 367440 513492 367474
rect 513391 367384 513492 367440
rect 513391 367350 513426 367384
rect 513460 367350 513492 367384
rect 513391 367294 513492 367350
rect 513391 367260 513426 367294
rect 513460 367260 513492 367294
rect 513391 367204 513492 367260
rect 513391 367170 513426 367204
rect 513460 367170 513492 367204
rect 513391 367114 513492 367170
rect 513391 367080 513426 367114
rect 513460 367080 513492 367114
rect 513391 367024 513492 367080
rect 513391 366990 513426 367024
rect 513460 366990 513492 367024
rect 513391 366934 513492 366990
rect 513391 366900 513426 366934
rect 513460 366900 513492 366934
rect 513391 366844 513492 366900
rect 516578 368329 516758 368416
rect 516578 367887 516617 368329
rect 516719 367887 516758 368329
rect 516578 367800 516758 367887
rect 527858 370093 528038 370180
rect 527858 369651 527897 370093
rect 527999 369651 528038 370093
rect 527858 369564 528038 369651
rect 531618 370191 531798 370278
rect 531618 369749 531657 370191
rect 531759 369749 531798 370191
rect 531618 369662 531798 369749
rect 513391 366810 513426 366844
rect 513460 366810 513492 366844
rect 513391 366754 513492 366810
rect 513391 366720 513426 366754
rect 513460 366720 513492 366754
rect 513391 366664 513492 366720
rect 512204 366597 512305 366630
rect 513391 366630 513426 366664
rect 513460 366630 513492 366664
rect 513391 366597 513492 366630
rect 512204 366563 513492 366597
rect 512204 366529 512262 366563
rect 512296 366529 512352 366563
rect 512386 366529 512442 366563
rect 512476 366529 512532 366563
rect 512566 366529 512622 366563
rect 512656 366529 512712 366563
rect 512746 366529 512802 366563
rect 512836 366529 512892 366563
rect 512926 366529 512982 366563
rect 513016 366529 513072 366563
rect 513106 366529 513162 366563
rect 513196 366529 513252 366563
rect 513286 366529 513342 366563
rect 513376 366529 513492 366563
rect 512204 366410 513492 366529
rect 512204 366376 512262 366410
rect 512296 366376 512352 366410
rect 512386 366376 512442 366410
rect 512476 366376 512532 366410
rect 512566 366376 512622 366410
rect 512656 366376 512712 366410
rect 512746 366376 512802 366410
rect 512836 366376 512892 366410
rect 512926 366376 512982 366410
rect 513016 366376 513072 366410
rect 513106 366376 513162 366410
rect 513196 366376 513252 366410
rect 513286 366376 513342 366410
rect 513376 366376 513492 366410
rect 512204 366343 513492 366376
rect 512204 366314 512305 366343
rect 512204 366280 512239 366314
rect 512273 366280 512305 366314
rect 513391 366314 513492 366343
rect 512204 366224 512305 366280
rect 512204 366190 512239 366224
rect 512273 366190 512305 366224
rect 512204 366134 512305 366190
rect 512204 366100 512239 366134
rect 512273 366100 512305 366134
rect 512204 366044 512305 366100
rect 512204 366010 512239 366044
rect 512273 366010 512305 366044
rect 512204 365954 512305 366010
rect 512204 365920 512239 365954
rect 512273 365920 512305 365954
rect 512204 365864 512305 365920
rect 512204 365830 512239 365864
rect 512273 365830 512305 365864
rect 512204 365774 512305 365830
rect 512204 365740 512239 365774
rect 512273 365740 512305 365774
rect 512204 365684 512305 365740
rect 512204 365650 512239 365684
rect 512273 365650 512305 365684
rect 512204 365594 512305 365650
rect 512204 365560 512239 365594
rect 512273 365560 512305 365594
rect 512204 365504 512305 365560
rect 512204 365470 512239 365504
rect 512273 365470 512305 365504
rect 512204 365414 512305 365470
rect 512204 365380 512239 365414
rect 512273 365380 512305 365414
rect 512204 365324 512305 365380
rect 512204 365290 512239 365324
rect 512273 365290 512305 365324
rect 513391 366280 513426 366314
rect 513460 366280 513492 366314
rect 513391 366224 513492 366280
rect 513391 366190 513426 366224
rect 513460 366190 513492 366224
rect 513391 366134 513492 366190
rect 513391 366100 513426 366134
rect 513460 366100 513492 366134
rect 513391 366044 513492 366100
rect 513391 366010 513426 366044
rect 513460 366010 513492 366044
rect 513391 365954 513492 366010
rect 513391 365920 513426 365954
rect 513460 365920 513492 365954
rect 513391 365864 513492 365920
rect 513391 365830 513426 365864
rect 513460 365830 513492 365864
rect 513391 365774 513492 365830
rect 513391 365740 513426 365774
rect 513460 365740 513492 365774
rect 513391 365684 513492 365740
rect 513391 365650 513426 365684
rect 513460 365650 513492 365684
rect 513391 365594 513492 365650
rect 513391 365560 513426 365594
rect 513460 365560 513492 365594
rect 513391 365504 513492 365560
rect 513391 365470 513426 365504
rect 513460 365470 513492 365504
rect 513391 365414 513492 365470
rect 513391 365380 513426 365414
rect 513460 365380 513492 365414
rect 513391 365324 513492 365380
rect 512204 365257 512305 365290
rect 513391 365290 513426 365324
rect 513460 365290 513492 365324
rect 513391 365257 513492 365290
rect 512204 365223 513492 365257
rect 512204 365189 512262 365223
rect 512296 365189 512352 365223
rect 512386 365189 512442 365223
rect 512476 365189 512532 365223
rect 512566 365189 512622 365223
rect 512656 365189 512712 365223
rect 512746 365189 512802 365223
rect 512836 365189 512892 365223
rect 512926 365189 512982 365223
rect 513016 365189 513072 365223
rect 513106 365189 513162 365223
rect 513196 365189 513252 365223
rect 513286 365189 513342 365223
rect 513376 365189 513492 365223
rect 512204 365070 513492 365189
rect 512204 365036 512262 365070
rect 512296 365036 512352 365070
rect 512386 365036 512442 365070
rect 512476 365036 512532 365070
rect 512566 365036 512622 365070
rect 512656 365036 512712 365070
rect 512746 365036 512802 365070
rect 512836 365036 512892 365070
rect 512926 365036 512982 365070
rect 513016 365036 513072 365070
rect 513106 365036 513162 365070
rect 513196 365036 513252 365070
rect 513286 365036 513342 365070
rect 513376 365036 513492 365070
rect 512204 365003 513492 365036
rect 512204 364974 512305 365003
rect 512204 364940 512239 364974
rect 512273 364940 512305 364974
rect 513391 364974 513492 365003
rect 512204 364884 512305 364940
rect 512204 364850 512239 364884
rect 512273 364850 512305 364884
rect 512204 364794 512305 364850
rect 512204 364760 512239 364794
rect 512273 364760 512305 364794
rect 512204 364704 512305 364760
rect 512204 364670 512239 364704
rect 512273 364670 512305 364704
rect 512204 364614 512305 364670
rect 512204 364580 512239 364614
rect 512273 364580 512305 364614
rect 512204 364524 512305 364580
rect 512204 364490 512239 364524
rect 512273 364490 512305 364524
rect 512204 364434 512305 364490
rect 512204 364400 512239 364434
rect 512273 364400 512305 364434
rect 512204 364344 512305 364400
rect 512204 364310 512239 364344
rect 512273 364310 512305 364344
rect 512204 364254 512305 364310
rect 512204 364220 512239 364254
rect 512273 364220 512305 364254
rect 512204 364164 512305 364220
rect 512204 364130 512239 364164
rect 512273 364130 512305 364164
rect 512204 364074 512305 364130
rect 512204 364040 512239 364074
rect 512273 364040 512305 364074
rect 512204 363984 512305 364040
rect 512204 363950 512239 363984
rect 512273 363950 512305 363984
rect 513391 364940 513426 364974
rect 513460 364940 513492 364974
rect 513391 364884 513492 364940
rect 513391 364850 513426 364884
rect 513460 364850 513492 364884
rect 513391 364794 513492 364850
rect 513391 364760 513426 364794
rect 513460 364760 513492 364794
rect 513391 364704 513492 364760
rect 513391 364670 513426 364704
rect 513460 364670 513492 364704
rect 513391 364614 513492 364670
rect 513391 364580 513426 364614
rect 513460 364580 513492 364614
rect 513391 364524 513492 364580
rect 513391 364490 513426 364524
rect 513460 364490 513492 364524
rect 513391 364434 513492 364490
rect 513391 364400 513426 364434
rect 513460 364400 513492 364434
rect 513391 364344 513492 364400
rect 513391 364310 513426 364344
rect 513460 364310 513492 364344
rect 513391 364254 513492 364310
rect 513391 364220 513426 364254
rect 513460 364220 513492 364254
rect 513391 364164 513492 364220
rect 513391 364130 513426 364164
rect 513460 364130 513492 364164
rect 516578 365585 516758 365672
rect 516578 365143 516617 365585
rect 516719 365143 516758 365585
rect 516578 365056 516758 365143
rect 520338 365585 520518 365672
rect 520338 365143 520377 365585
rect 520479 365143 520518 365585
rect 520338 365056 520518 365143
rect 527858 367349 528038 367436
rect 527858 366907 527897 367349
rect 527999 366907 528038 367349
rect 527858 366820 528038 366907
rect 531618 367447 531798 367534
rect 531618 367005 531657 367447
rect 531759 367005 531798 367447
rect 531618 366918 531798 367005
rect 535378 369407 535558 369494
rect 535378 368965 535417 369407
rect 535519 368965 535558 369407
rect 535378 368878 535558 368965
rect 513391 364074 513492 364130
rect 513391 364040 513426 364074
rect 513460 364040 513492 364074
rect 513391 363984 513492 364040
rect 512204 363917 512305 363950
rect 513391 363950 513426 363984
rect 513460 363950 513492 363984
rect 513391 363917 513492 363950
rect 512204 363883 513492 363917
rect 512204 363849 512262 363883
rect 512296 363849 512352 363883
rect 512386 363849 512442 363883
rect 512476 363849 512532 363883
rect 512566 363849 512622 363883
rect 512656 363849 512712 363883
rect 512746 363849 512802 363883
rect 512836 363849 512892 363883
rect 512926 363849 512982 363883
rect 513016 363849 513072 363883
rect 513106 363849 513162 363883
rect 513196 363849 513252 363883
rect 513286 363849 513342 363883
rect 513376 363849 513492 363883
rect 512204 363730 513492 363849
rect 512204 363696 512262 363730
rect 512296 363696 512352 363730
rect 512386 363696 512442 363730
rect 512476 363696 512532 363730
rect 512566 363696 512622 363730
rect 512656 363696 512712 363730
rect 512746 363696 512802 363730
rect 512836 363696 512892 363730
rect 512926 363696 512982 363730
rect 513016 363696 513072 363730
rect 513106 363696 513162 363730
rect 513196 363696 513252 363730
rect 513286 363696 513342 363730
rect 513376 363696 513492 363730
rect 512204 363663 513492 363696
rect 512204 363634 512305 363663
rect 512204 363600 512239 363634
rect 512273 363600 512305 363634
rect 513391 363634 513492 363663
rect 512204 363544 512305 363600
rect 512204 363510 512239 363544
rect 512273 363510 512305 363544
rect 512204 363454 512305 363510
rect 512204 363420 512239 363454
rect 512273 363420 512305 363454
rect 512204 363364 512305 363420
rect 512204 363330 512239 363364
rect 512273 363330 512305 363364
rect 512204 363274 512305 363330
rect 512204 363240 512239 363274
rect 512273 363240 512305 363274
rect 512204 363184 512305 363240
rect 512204 363150 512239 363184
rect 512273 363150 512305 363184
rect 512204 363094 512305 363150
rect 512204 363060 512239 363094
rect 512273 363060 512305 363094
rect 512204 363004 512305 363060
rect 512204 362970 512239 363004
rect 512273 362970 512305 363004
rect 512204 362914 512305 362970
rect 512204 362880 512239 362914
rect 512273 362880 512305 362914
rect 512204 362824 512305 362880
rect 512204 362790 512239 362824
rect 512273 362790 512305 362824
rect 512204 362734 512305 362790
rect 512204 362700 512239 362734
rect 512273 362700 512305 362734
rect 512204 362644 512305 362700
rect 512204 362610 512239 362644
rect 512273 362610 512305 362644
rect 513391 363600 513426 363634
rect 513460 363600 513492 363634
rect 513391 363544 513492 363600
rect 513391 363510 513426 363544
rect 513460 363510 513492 363544
rect 513391 363454 513492 363510
rect 513391 363420 513426 363454
rect 513460 363420 513492 363454
rect 513391 363364 513492 363420
rect 513391 363330 513426 363364
rect 513460 363330 513492 363364
rect 513391 363274 513492 363330
rect 513391 363240 513426 363274
rect 513460 363240 513492 363274
rect 513391 363184 513492 363240
rect 513391 363150 513426 363184
rect 513460 363150 513492 363184
rect 513391 363094 513492 363150
rect 513391 363060 513426 363094
rect 513460 363060 513492 363094
rect 527858 364605 528038 364692
rect 527858 364163 527897 364605
rect 527999 364163 528038 364605
rect 527858 364076 528038 364163
rect 531618 364703 531798 364790
rect 531618 364261 531657 364703
rect 531759 364261 531798 364703
rect 531618 364174 531798 364261
rect 535378 366663 535558 366750
rect 535378 366221 535417 366663
rect 535519 366221 535558 366663
rect 535378 366134 535558 366221
rect 513391 363004 513492 363060
rect 513391 362970 513426 363004
rect 513460 362970 513492 363004
rect 513391 362914 513492 362970
rect 513391 362880 513426 362914
rect 513460 362880 513492 362914
rect 513391 362824 513492 362880
rect 513391 362790 513426 362824
rect 513460 362790 513492 362824
rect 513391 362734 513492 362790
rect 513391 362700 513426 362734
rect 513460 362700 513492 362734
rect 513391 362644 513492 362700
rect 512204 362577 512305 362610
rect 513391 362610 513426 362644
rect 513460 362610 513492 362644
rect 513391 362577 513492 362610
rect 512204 362543 513492 362577
rect 512204 362509 512262 362543
rect 512296 362509 512352 362543
rect 512386 362509 512442 362543
rect 512476 362509 512532 362543
rect 512566 362509 512622 362543
rect 512656 362509 512712 362543
rect 512746 362509 512802 362543
rect 512836 362509 512892 362543
rect 512926 362509 512982 362543
rect 513016 362509 513072 362543
rect 513106 362509 513162 362543
rect 513196 362509 513252 362543
rect 513286 362509 513342 362543
rect 513376 362509 513492 362543
rect 535378 363919 535558 364006
rect 535378 363477 535417 363919
rect 535519 363477 535558 363919
rect 535378 363390 535558 363477
rect 512204 362476 513492 362509
rect 565778 357640 565818 357680
rect 562040 357608 562160 357610
rect 562040 357572 562076 357608
rect 562120 357572 562160 357608
rect 562040 357560 562160 357572
rect 563340 357608 563460 357610
rect 563340 357572 563376 357608
rect 563420 357572 563460 357608
rect 563340 357560 563460 357572
rect 564640 357608 564760 357610
rect 564640 357572 564676 357608
rect 564720 357572 564760 357608
rect 564640 357560 564760 357572
rect 565778 357560 565818 357600
rect 565640 311332 565680 311372
rect 561902 311300 562022 311302
rect 561902 311264 561938 311300
rect 561982 311264 562022 311300
rect 561902 311252 562022 311264
rect 563202 311300 563322 311302
rect 563202 311264 563238 311300
rect 563282 311264 563322 311300
rect 563202 311252 563322 311264
rect 564502 311300 564622 311302
rect 564502 311264 564538 311300
rect 564582 311264 564622 311300
rect 564502 311252 564622 311264
rect 565640 311252 565680 311292
<< nsubdiff >>
rect 576740 493522 576860 493524
rect 576740 493486 576776 493522
rect 576820 493486 576860 493522
rect 576740 493484 576860 493486
rect 578040 493522 578160 493524
rect 578040 493486 578076 493522
rect 578120 493486 578160 493522
rect 578040 493484 578160 493486
rect 579340 493522 579460 493524
rect 579340 493486 579376 493522
rect 579420 493486 579460 493522
rect 579340 493484 579460 493486
rect 580478 493474 580518 493514
rect 580478 493394 580518 493434
rect 576018 404646 576138 404648
rect 576018 404610 576054 404646
rect 576098 404610 576138 404646
rect 576018 404608 576138 404610
rect 577318 404646 577438 404648
rect 577318 404610 577354 404646
rect 577398 404610 577438 404646
rect 577318 404608 577438 404610
rect 578618 404646 578738 404648
rect 578618 404610 578654 404646
rect 578698 404610 578738 404646
rect 578618 404608 578738 404610
rect 579756 404598 579796 404638
rect 579756 404518 579796 404558
rect 504847 402754 505809 402773
rect 504847 402720 504923 402754
rect 504957 402720 505013 402754
rect 505047 402720 505103 402754
rect 505137 402720 505193 402754
rect 505227 402720 505283 402754
rect 505317 402720 505373 402754
rect 505407 402720 505463 402754
rect 505497 402720 505553 402754
rect 505587 402720 505643 402754
rect 505677 402720 505809 402754
rect 504847 402701 505809 402720
rect 504847 402642 504919 402701
rect 504847 402608 504866 402642
rect 504900 402608 504919 402642
rect 505737 402676 505809 402701
rect 505737 402642 505756 402676
rect 505790 402642 505809 402676
rect 504847 402552 504919 402608
rect 504847 402518 504866 402552
rect 504900 402518 504919 402552
rect 504847 402462 504919 402518
rect 504847 402428 504866 402462
rect 504900 402428 504919 402462
rect 504847 402372 504919 402428
rect 504847 402338 504866 402372
rect 504900 402338 504919 402372
rect 504847 402282 504919 402338
rect 504847 402248 504866 402282
rect 504900 402248 504919 402282
rect 504847 402192 504919 402248
rect 504847 402158 504866 402192
rect 504900 402158 504919 402192
rect 504847 402102 504919 402158
rect 504847 402068 504866 402102
rect 504900 402068 504919 402102
rect 504847 402012 504919 402068
rect 504847 401978 504866 402012
rect 504900 401978 504919 402012
rect 504847 401922 504919 401978
rect 505737 402586 505809 402642
rect 505737 402552 505756 402586
rect 505790 402552 505809 402586
rect 505737 402496 505809 402552
rect 505737 402462 505756 402496
rect 505790 402462 505809 402496
rect 505737 402406 505809 402462
rect 505737 402372 505756 402406
rect 505790 402372 505809 402406
rect 505737 402316 505809 402372
rect 505737 402282 505756 402316
rect 505790 402282 505809 402316
rect 505737 402226 505809 402282
rect 505737 402192 505756 402226
rect 505790 402192 505809 402226
rect 505737 402136 505809 402192
rect 505737 402102 505756 402136
rect 505790 402102 505809 402136
rect 505737 402046 505809 402102
rect 505737 402012 505756 402046
rect 505790 402012 505809 402046
rect 505737 401956 505809 402012
rect 504847 401888 504866 401922
rect 504900 401888 504919 401922
rect 504847 401883 504919 401888
rect 505737 401922 505756 401956
rect 505790 401922 505809 401956
rect 505737 401883 505809 401922
rect 504847 401864 505809 401883
rect 504847 401830 504942 401864
rect 504976 401830 505032 401864
rect 505066 401830 505122 401864
rect 505156 401830 505212 401864
rect 505246 401830 505302 401864
rect 505336 401830 505392 401864
rect 505426 401830 505482 401864
rect 505516 401830 505572 401864
rect 505606 401830 505662 401864
rect 505696 401830 505809 401864
rect 504847 401811 505809 401830
rect 496948 399981 497068 399984
rect 496948 399947 496991 399981
rect 497025 399947 497068 399981
rect 496948 399944 497068 399947
rect 496938 398881 496978 398926
rect 496938 398847 496941 398881
rect 496975 398847 496978 398881
rect 496938 398806 496978 398847
rect 496938 397581 496978 397626
rect 496938 397547 496941 397581
rect 496975 397547 496978 397581
rect 496938 397506 496978 397547
rect 496938 396281 496978 396326
rect 496938 396247 496941 396281
rect 496975 396247 496978 396281
rect 496938 396206 496978 396247
rect 496938 394981 496978 395026
rect 496938 394947 496941 394981
rect 496975 394947 496978 394981
rect 496938 394906 496978 394947
rect 496938 393681 496978 393726
rect 496938 393647 496941 393681
rect 496975 393647 496978 393681
rect 496938 393606 496978 393647
rect 496938 392381 496978 392426
rect 496938 392347 496941 392381
rect 496975 392347 496978 392381
rect 496938 392306 496978 392347
rect 500708 392337 500828 392340
rect 500708 392303 500751 392337
rect 500785 392303 500828 392337
rect 500708 392300 500828 392303
rect 496938 391081 496978 391126
rect 496938 391047 496941 391081
rect 496975 391047 496978 391081
rect 496938 391006 496978 391047
rect 500698 391237 500738 391282
rect 500698 391203 500701 391237
rect 500735 391203 500738 391237
rect 500698 391162 500738 391203
rect 493188 390181 493308 390184
rect 493188 390147 493231 390181
rect 493265 390147 493308 390181
rect 493188 390144 493308 390147
rect 496938 389781 496978 389826
rect 496938 389747 496941 389781
rect 496975 389747 496978 389781
rect 496938 389706 496978 389747
rect 500698 389937 500738 389982
rect 500698 389903 500701 389937
rect 500735 389903 500738 389937
rect 500698 389862 500738 389903
rect 493178 389081 493218 389126
rect 493178 389047 493181 389081
rect 493215 389047 493218 389081
rect 493178 389006 493218 389047
rect 496938 388481 496978 388526
rect 496938 388447 496941 388481
rect 496975 388447 496978 388481
rect 496938 388406 496978 388447
rect 500698 388637 500738 388682
rect 500698 388603 500701 388637
rect 500735 388603 500738 388637
rect 500698 388562 500738 388603
rect 493178 387781 493218 387826
rect 493178 387747 493181 387781
rect 493215 387747 493218 387781
rect 493178 387706 493218 387747
rect 523268 390181 523388 390184
rect 523268 390147 523311 390181
rect 523345 390147 523388 390181
rect 523268 390144 523388 390147
rect 523258 389081 523298 389126
rect 523258 389047 523261 389081
rect 523295 389047 523298 389081
rect 523258 389006 523298 389047
rect 496938 387181 496978 387226
rect 496938 387147 496941 387181
rect 496975 387147 496978 387181
rect 496938 387106 496978 387147
rect 493178 386481 493218 386526
rect 493178 386447 493181 386481
rect 493215 386447 493218 386481
rect 493178 386406 493218 386447
rect 496938 385881 496978 385926
rect 496938 385847 496941 385881
rect 496975 385847 496978 385881
rect 496938 385806 496978 385847
rect 493178 385181 493218 385226
rect 493178 385147 493181 385181
rect 493215 385147 493218 385181
rect 493178 385106 493218 385147
rect 500708 385673 500828 385676
rect 500708 385639 500751 385673
rect 500785 385639 500828 385673
rect 500708 385636 500828 385639
rect 523258 387781 523298 387826
rect 523258 387747 523261 387781
rect 523295 387747 523298 387781
rect 523258 387706 523298 387747
rect 523258 386481 523298 386526
rect 523258 386447 523261 386481
rect 523295 386447 523298 386481
rect 523258 386406 523298 386447
rect 496938 384581 496978 384626
rect 496938 384547 496941 384581
rect 496975 384547 496978 384581
rect 496938 384506 496978 384547
rect 523258 385181 523298 385226
rect 523258 385147 523261 385181
rect 523295 385147 523298 385181
rect 523258 385106 523298 385147
rect 493178 383881 493218 383926
rect 493178 383847 493181 383881
rect 493215 383847 493218 383881
rect 493178 383806 493218 383847
rect 500698 384573 500738 384618
rect 500698 384539 500701 384573
rect 500735 384539 500738 384573
rect 500698 384498 500738 384539
rect 496938 383281 496978 383326
rect 496938 383247 496941 383281
rect 496975 383247 496978 383281
rect 496938 383206 496978 383247
rect 500698 383273 500738 383318
rect 500698 383239 500701 383273
rect 500735 383239 500738 383273
rect 500698 383198 500738 383239
rect 493178 382581 493218 382626
rect 493178 382547 493181 382581
rect 493215 382547 493218 382581
rect 493178 382506 493218 382547
rect 523258 383881 523298 383926
rect 523258 383847 523261 383881
rect 523295 383847 523298 383881
rect 523258 383806 523298 383847
rect 523258 382581 523298 382626
rect 496938 381981 496978 382026
rect 496938 381947 496941 381981
rect 496975 381947 496978 381981
rect 496938 381906 496978 381947
rect 500698 381973 500738 382018
rect 500698 381939 500701 381973
rect 500735 381939 500738 381973
rect 500698 381898 500738 381939
rect 523258 382547 523261 382581
rect 523295 382547 523298 382581
rect 523258 382506 523298 382547
rect 493178 381281 493218 381326
rect 493178 381247 493181 381281
rect 493215 381247 493218 381281
rect 493178 381206 493218 381247
rect 493178 379981 493218 380026
rect 496938 380681 496978 380726
rect 496938 380647 496941 380681
rect 496975 380647 496978 380681
rect 496938 380606 496978 380647
rect 493178 379947 493181 379981
rect 493215 379947 493218 379981
rect 493178 379906 493218 379947
rect 496938 379381 496978 379426
rect 496938 379347 496941 379381
rect 496975 379347 496978 379381
rect 496938 379306 496978 379347
rect 523258 381281 523298 381326
rect 523258 381247 523261 381281
rect 523295 381247 523298 381281
rect 523258 381206 523298 381247
rect 523258 379981 523298 380026
rect 523258 379947 523261 379981
rect 523295 379947 523298 379981
rect 523258 379906 523298 379947
rect 493178 378681 493218 378726
rect 493178 378647 493181 378681
rect 493215 378647 493218 378681
rect 493178 378606 493218 378647
rect 523258 378681 523298 378726
rect 523258 378647 523261 378681
rect 523295 378647 523298 378681
rect 523258 378606 523298 378647
rect 496938 378081 496978 378126
rect 496938 378047 496941 378081
rect 496975 378047 496978 378081
rect 496938 378006 496978 378047
rect 493178 377381 493218 377426
rect 493178 377347 493181 377381
rect 493215 377347 493218 377381
rect 493178 377306 493218 377347
rect 504468 377539 504588 377542
rect 504468 377505 504511 377539
rect 504545 377505 504588 377539
rect 504468 377502 504588 377505
rect 511988 377539 512108 377542
rect 511988 377505 512031 377539
rect 512065 377505 512108 377539
rect 511988 377502 512108 377505
rect 496938 376781 496978 376826
rect 496938 376747 496941 376781
rect 496975 376747 496978 376781
rect 496938 376706 496978 376747
rect 493178 376081 493218 376126
rect 493178 376047 493181 376081
rect 493215 376047 493218 376081
rect 493178 376006 493218 376047
rect 504458 376439 504498 376484
rect 504458 376405 504461 376439
rect 504495 376405 504498 376439
rect 504458 376364 504498 376405
rect 511978 376439 512018 376484
rect 511978 376405 511981 376439
rect 512015 376405 512018 376439
rect 511978 376364 512018 376405
rect 496938 375481 496978 375526
rect 496938 375447 496941 375481
rect 496975 375447 496978 375481
rect 496938 375406 496978 375447
rect 493178 374781 493218 374826
rect 493178 374747 493181 374781
rect 493215 374747 493218 374781
rect 493178 374706 493218 374747
rect 496938 374181 496978 374226
rect 496938 374147 496941 374181
rect 496975 374147 496978 374181
rect 496938 374106 496978 374147
rect 493178 373481 493218 373526
rect 493178 373447 493181 373481
rect 493215 373447 493218 373481
rect 493178 373406 493218 373447
rect 523258 377381 523298 377426
rect 523258 377347 523261 377381
rect 523295 377347 523298 377381
rect 523258 377306 523298 377347
rect 523258 376081 523298 376126
rect 523258 376047 523261 376081
rect 523295 376047 523298 376081
rect 523258 376006 523298 376047
rect 493178 372181 493218 372226
rect 493178 372147 493181 372181
rect 493215 372147 493218 372181
rect 493178 372106 493218 372147
rect 501087 372962 502049 372981
rect 501087 372928 501163 372962
rect 501197 372928 501253 372962
rect 501287 372928 501343 372962
rect 501377 372928 501433 372962
rect 501467 372928 501523 372962
rect 501557 372928 501613 372962
rect 501647 372928 501703 372962
rect 501737 372928 501793 372962
rect 501827 372928 501883 372962
rect 501917 372928 502049 372962
rect 501087 372909 502049 372928
rect 501087 372850 501159 372909
rect 501087 372816 501106 372850
rect 501140 372816 501159 372850
rect 501977 372884 502049 372909
rect 501977 372850 501996 372884
rect 502030 372850 502049 372884
rect 501087 372760 501159 372816
rect 501087 372726 501106 372760
rect 501140 372726 501159 372760
rect 501087 372670 501159 372726
rect 501087 372636 501106 372670
rect 501140 372636 501159 372670
rect 501087 372580 501159 372636
rect 501087 372546 501106 372580
rect 501140 372546 501159 372580
rect 501087 372490 501159 372546
rect 501087 372456 501106 372490
rect 501140 372456 501159 372490
rect 501087 372400 501159 372456
rect 501087 372366 501106 372400
rect 501140 372366 501159 372400
rect 501087 372310 501159 372366
rect 501087 372276 501106 372310
rect 501140 372276 501159 372310
rect 501087 372220 501159 372276
rect 501087 372186 501106 372220
rect 501140 372186 501159 372220
rect 501087 372130 501159 372186
rect 501977 372794 502049 372850
rect 501977 372760 501996 372794
rect 502030 372760 502049 372794
rect 501977 372704 502049 372760
rect 501977 372670 501996 372704
rect 502030 372670 502049 372704
rect 501977 372614 502049 372670
rect 501977 372580 501996 372614
rect 502030 372580 502049 372614
rect 501977 372524 502049 372580
rect 501977 372490 501996 372524
rect 502030 372490 502049 372524
rect 501977 372434 502049 372490
rect 501977 372400 501996 372434
rect 502030 372400 502049 372434
rect 501977 372344 502049 372400
rect 501977 372310 501996 372344
rect 502030 372310 502049 372344
rect 501977 372254 502049 372310
rect 501977 372220 501996 372254
rect 502030 372220 502049 372254
rect 501977 372164 502049 372220
rect 501087 372096 501106 372130
rect 501140 372096 501159 372130
rect 501087 372091 501159 372096
rect 501977 372130 501996 372164
rect 502030 372130 502049 372164
rect 501977 372091 502049 372130
rect 501087 372072 502049 372091
rect 501087 372038 501182 372072
rect 501216 372038 501272 372072
rect 501306 372038 501362 372072
rect 501396 372038 501452 372072
rect 501486 372038 501542 372072
rect 501576 372038 501632 372072
rect 501666 372038 501722 372072
rect 501756 372038 501812 372072
rect 501846 372038 501902 372072
rect 501936 372038 502049 372072
rect 501087 372019 502049 372038
rect 493178 370881 493218 370926
rect 493178 370847 493181 370881
rect 493215 370847 493218 370881
rect 493178 370806 493218 370847
rect 493178 369581 493218 369626
rect 493178 369547 493181 369581
rect 493215 369547 493218 369581
rect 493178 369506 493218 369547
rect 493178 368281 493218 368326
rect 493178 368247 493181 368281
rect 493215 368247 493218 368281
rect 493178 368206 493218 368247
rect 493178 366981 493218 367026
rect 493178 366947 493181 366981
rect 493215 366947 493218 366981
rect 493178 366906 493218 366947
rect 493178 365681 493218 365726
rect 493178 365647 493181 365681
rect 493215 365647 493218 365681
rect 493178 365606 493218 365647
rect 493178 364381 493218 364426
rect 493178 364347 493181 364381
rect 493215 364347 493218 364381
rect 493178 364306 493218 364347
rect 497327 371786 498289 371805
rect 497327 371752 497403 371786
rect 497437 371752 497493 371786
rect 497527 371752 497583 371786
rect 497617 371752 497673 371786
rect 497707 371752 497763 371786
rect 497797 371752 497853 371786
rect 497887 371752 497943 371786
rect 497977 371752 498033 371786
rect 498067 371752 498123 371786
rect 498157 371752 498289 371786
rect 497327 371733 498289 371752
rect 497327 371674 497399 371733
rect 497327 371640 497346 371674
rect 497380 371640 497399 371674
rect 498217 371708 498289 371733
rect 498217 371674 498236 371708
rect 498270 371674 498289 371708
rect 497327 371584 497399 371640
rect 497327 371550 497346 371584
rect 497380 371550 497399 371584
rect 497327 371494 497399 371550
rect 497327 371460 497346 371494
rect 497380 371460 497399 371494
rect 497327 371404 497399 371460
rect 497327 371370 497346 371404
rect 497380 371370 497399 371404
rect 497327 371314 497399 371370
rect 497327 371280 497346 371314
rect 497380 371280 497399 371314
rect 497327 371224 497399 371280
rect 497327 371190 497346 371224
rect 497380 371190 497399 371224
rect 497327 371134 497399 371190
rect 497327 371100 497346 371134
rect 497380 371100 497399 371134
rect 497327 371044 497399 371100
rect 497327 371010 497346 371044
rect 497380 371010 497399 371044
rect 497327 370954 497399 371010
rect 498217 371618 498289 371674
rect 498217 371584 498236 371618
rect 498270 371584 498289 371618
rect 498217 371528 498289 371584
rect 498217 371494 498236 371528
rect 498270 371494 498289 371528
rect 498217 371438 498289 371494
rect 498217 371404 498236 371438
rect 498270 371404 498289 371438
rect 498217 371348 498289 371404
rect 498217 371314 498236 371348
rect 498270 371314 498289 371348
rect 498217 371258 498289 371314
rect 498217 371224 498236 371258
rect 498270 371224 498289 371258
rect 498217 371168 498289 371224
rect 498217 371134 498236 371168
rect 498270 371134 498289 371168
rect 498217 371078 498289 371134
rect 498217 371044 498236 371078
rect 498270 371044 498289 371078
rect 498217 370988 498289 371044
rect 497327 370920 497346 370954
rect 497380 370920 497399 370954
rect 497327 370915 497399 370920
rect 498217 370954 498236 370988
rect 498270 370954 498289 370988
rect 498217 370915 498289 370954
rect 497327 370896 498289 370915
rect 497327 370862 497422 370896
rect 497456 370862 497512 370896
rect 497546 370862 497602 370896
rect 497636 370862 497692 370896
rect 497726 370862 497782 370896
rect 497816 370862 497872 370896
rect 497906 370862 497962 370896
rect 497996 370862 498052 370896
rect 498086 370862 498142 370896
rect 498176 370862 498289 370896
rect 497327 370843 498289 370862
rect 497327 370446 498289 370465
rect 497327 370412 497403 370446
rect 497437 370412 497493 370446
rect 497527 370412 497583 370446
rect 497617 370412 497673 370446
rect 497707 370412 497763 370446
rect 497797 370412 497853 370446
rect 497887 370412 497943 370446
rect 497977 370412 498033 370446
rect 498067 370412 498123 370446
rect 498157 370412 498289 370446
rect 497327 370393 498289 370412
rect 497327 370334 497399 370393
rect 497327 370300 497346 370334
rect 497380 370300 497399 370334
rect 498217 370368 498289 370393
rect 498217 370334 498236 370368
rect 498270 370334 498289 370368
rect 497327 370244 497399 370300
rect 497327 370210 497346 370244
rect 497380 370210 497399 370244
rect 497327 370154 497399 370210
rect 497327 370120 497346 370154
rect 497380 370120 497399 370154
rect 497327 370064 497399 370120
rect 497327 370030 497346 370064
rect 497380 370030 497399 370064
rect 497327 369974 497399 370030
rect 497327 369940 497346 369974
rect 497380 369940 497399 369974
rect 497327 369884 497399 369940
rect 497327 369850 497346 369884
rect 497380 369850 497399 369884
rect 497327 369794 497399 369850
rect 497327 369760 497346 369794
rect 497380 369760 497399 369794
rect 497327 369704 497399 369760
rect 497327 369670 497346 369704
rect 497380 369670 497399 369704
rect 497327 369614 497399 369670
rect 498217 370278 498289 370334
rect 498217 370244 498236 370278
rect 498270 370244 498289 370278
rect 498217 370188 498289 370244
rect 498217 370154 498236 370188
rect 498270 370154 498289 370188
rect 498217 370098 498289 370154
rect 498217 370064 498236 370098
rect 498270 370064 498289 370098
rect 498217 370008 498289 370064
rect 498217 369974 498236 370008
rect 498270 369974 498289 370008
rect 498217 369918 498289 369974
rect 498217 369884 498236 369918
rect 498270 369884 498289 369918
rect 498217 369828 498289 369884
rect 498217 369794 498236 369828
rect 498270 369794 498289 369828
rect 498217 369738 498289 369794
rect 498217 369704 498236 369738
rect 498270 369704 498289 369738
rect 498217 369648 498289 369704
rect 497327 369580 497346 369614
rect 497380 369580 497399 369614
rect 497327 369575 497399 369580
rect 498217 369614 498236 369648
rect 498270 369614 498289 369648
rect 498217 369575 498289 369614
rect 497327 369556 498289 369575
rect 497327 369522 497422 369556
rect 497456 369522 497512 369556
rect 497546 369522 497602 369556
rect 497636 369522 497692 369556
rect 497726 369522 497782 369556
rect 497816 369522 497872 369556
rect 497906 369522 497962 369556
rect 497996 369522 498052 369556
rect 498086 369522 498142 369556
rect 498176 369522 498289 369556
rect 497327 369503 498289 369522
rect 497327 369106 498289 369125
rect 497327 369072 497403 369106
rect 497437 369072 497493 369106
rect 497527 369072 497583 369106
rect 497617 369072 497673 369106
rect 497707 369072 497763 369106
rect 497797 369072 497853 369106
rect 497887 369072 497943 369106
rect 497977 369072 498033 369106
rect 498067 369072 498123 369106
rect 498157 369072 498289 369106
rect 497327 369053 498289 369072
rect 497327 368994 497399 369053
rect 497327 368960 497346 368994
rect 497380 368960 497399 368994
rect 498217 369028 498289 369053
rect 498217 368994 498236 369028
rect 498270 368994 498289 369028
rect 497327 368904 497399 368960
rect 497327 368870 497346 368904
rect 497380 368870 497399 368904
rect 497327 368814 497399 368870
rect 497327 368780 497346 368814
rect 497380 368780 497399 368814
rect 497327 368724 497399 368780
rect 497327 368690 497346 368724
rect 497380 368690 497399 368724
rect 497327 368634 497399 368690
rect 497327 368600 497346 368634
rect 497380 368600 497399 368634
rect 497327 368544 497399 368600
rect 497327 368510 497346 368544
rect 497380 368510 497399 368544
rect 497327 368454 497399 368510
rect 497327 368420 497346 368454
rect 497380 368420 497399 368454
rect 497327 368364 497399 368420
rect 497327 368330 497346 368364
rect 497380 368330 497399 368364
rect 497327 368274 497399 368330
rect 498217 368938 498289 368994
rect 498217 368904 498236 368938
rect 498270 368904 498289 368938
rect 498217 368848 498289 368904
rect 498217 368814 498236 368848
rect 498270 368814 498289 368848
rect 498217 368758 498289 368814
rect 498217 368724 498236 368758
rect 498270 368724 498289 368758
rect 498217 368668 498289 368724
rect 498217 368634 498236 368668
rect 498270 368634 498289 368668
rect 498217 368578 498289 368634
rect 498217 368544 498236 368578
rect 498270 368544 498289 368578
rect 498217 368488 498289 368544
rect 498217 368454 498236 368488
rect 498270 368454 498289 368488
rect 498217 368398 498289 368454
rect 498217 368364 498236 368398
rect 498270 368364 498289 368398
rect 498217 368308 498289 368364
rect 497327 368240 497346 368274
rect 497380 368240 497399 368274
rect 497327 368235 497399 368240
rect 498217 368274 498236 368308
rect 498270 368274 498289 368308
rect 498217 368235 498289 368274
rect 497327 368216 498289 368235
rect 497327 368182 497422 368216
rect 497456 368182 497512 368216
rect 497546 368182 497602 368216
rect 497636 368182 497692 368216
rect 497726 368182 497782 368216
rect 497816 368182 497872 368216
rect 497906 368182 497962 368216
rect 497996 368182 498052 368216
rect 498086 368182 498142 368216
rect 498176 368182 498289 368216
rect 497327 368163 498289 368182
rect 497327 367766 498289 367785
rect 497327 367732 497403 367766
rect 497437 367732 497493 367766
rect 497527 367732 497583 367766
rect 497617 367732 497673 367766
rect 497707 367732 497763 367766
rect 497797 367732 497853 367766
rect 497887 367732 497943 367766
rect 497977 367732 498033 367766
rect 498067 367732 498123 367766
rect 498157 367732 498289 367766
rect 497327 367713 498289 367732
rect 497327 367654 497399 367713
rect 497327 367620 497346 367654
rect 497380 367620 497399 367654
rect 498217 367688 498289 367713
rect 498217 367654 498236 367688
rect 498270 367654 498289 367688
rect 497327 367564 497399 367620
rect 497327 367530 497346 367564
rect 497380 367530 497399 367564
rect 497327 367474 497399 367530
rect 497327 367440 497346 367474
rect 497380 367440 497399 367474
rect 497327 367384 497399 367440
rect 497327 367350 497346 367384
rect 497380 367350 497399 367384
rect 497327 367294 497399 367350
rect 497327 367260 497346 367294
rect 497380 367260 497399 367294
rect 497327 367204 497399 367260
rect 497327 367170 497346 367204
rect 497380 367170 497399 367204
rect 497327 367114 497399 367170
rect 497327 367080 497346 367114
rect 497380 367080 497399 367114
rect 497327 367024 497399 367080
rect 497327 366990 497346 367024
rect 497380 366990 497399 367024
rect 497327 366934 497399 366990
rect 498217 367598 498289 367654
rect 498217 367564 498236 367598
rect 498270 367564 498289 367598
rect 498217 367508 498289 367564
rect 498217 367474 498236 367508
rect 498270 367474 498289 367508
rect 498217 367418 498289 367474
rect 498217 367384 498236 367418
rect 498270 367384 498289 367418
rect 498217 367328 498289 367384
rect 498217 367294 498236 367328
rect 498270 367294 498289 367328
rect 498217 367238 498289 367294
rect 498217 367204 498236 367238
rect 498270 367204 498289 367238
rect 498217 367148 498289 367204
rect 498217 367114 498236 367148
rect 498270 367114 498289 367148
rect 498217 367058 498289 367114
rect 498217 367024 498236 367058
rect 498270 367024 498289 367058
rect 498217 366968 498289 367024
rect 497327 366900 497346 366934
rect 497380 366900 497399 366934
rect 497327 366895 497399 366900
rect 498217 366934 498236 366968
rect 498270 366934 498289 366968
rect 498217 366895 498289 366934
rect 497327 366876 498289 366895
rect 497327 366842 497422 366876
rect 497456 366842 497512 366876
rect 497546 366842 497602 366876
rect 497636 366842 497692 366876
rect 497726 366842 497782 366876
rect 497816 366842 497872 366876
rect 497906 366842 497962 366876
rect 497996 366842 498052 366876
rect 498086 366842 498142 366876
rect 498176 366842 498289 366876
rect 497327 366823 498289 366842
rect 497327 366426 498289 366445
rect 497327 366392 497403 366426
rect 497437 366392 497493 366426
rect 497527 366392 497583 366426
rect 497617 366392 497673 366426
rect 497707 366392 497763 366426
rect 497797 366392 497853 366426
rect 497887 366392 497943 366426
rect 497977 366392 498033 366426
rect 498067 366392 498123 366426
rect 498157 366392 498289 366426
rect 497327 366373 498289 366392
rect 497327 366314 497399 366373
rect 497327 366280 497346 366314
rect 497380 366280 497399 366314
rect 498217 366348 498289 366373
rect 498217 366314 498236 366348
rect 498270 366314 498289 366348
rect 497327 366224 497399 366280
rect 497327 366190 497346 366224
rect 497380 366190 497399 366224
rect 497327 366134 497399 366190
rect 497327 366100 497346 366134
rect 497380 366100 497399 366134
rect 497327 366044 497399 366100
rect 497327 366010 497346 366044
rect 497380 366010 497399 366044
rect 497327 365954 497399 366010
rect 497327 365920 497346 365954
rect 497380 365920 497399 365954
rect 497327 365864 497399 365920
rect 497327 365830 497346 365864
rect 497380 365830 497399 365864
rect 497327 365774 497399 365830
rect 497327 365740 497346 365774
rect 497380 365740 497399 365774
rect 497327 365684 497399 365740
rect 497327 365650 497346 365684
rect 497380 365650 497399 365684
rect 497327 365594 497399 365650
rect 498217 366258 498289 366314
rect 498217 366224 498236 366258
rect 498270 366224 498289 366258
rect 498217 366168 498289 366224
rect 498217 366134 498236 366168
rect 498270 366134 498289 366168
rect 498217 366078 498289 366134
rect 498217 366044 498236 366078
rect 498270 366044 498289 366078
rect 498217 365988 498289 366044
rect 498217 365954 498236 365988
rect 498270 365954 498289 365988
rect 498217 365898 498289 365954
rect 498217 365864 498236 365898
rect 498270 365864 498289 365898
rect 498217 365808 498289 365864
rect 498217 365774 498236 365808
rect 498270 365774 498289 365808
rect 498217 365718 498289 365774
rect 498217 365684 498236 365718
rect 498270 365684 498289 365718
rect 498217 365628 498289 365684
rect 497327 365560 497346 365594
rect 497380 365560 497399 365594
rect 497327 365555 497399 365560
rect 498217 365594 498236 365628
rect 498270 365594 498289 365628
rect 498217 365555 498289 365594
rect 497327 365536 498289 365555
rect 497327 365502 497422 365536
rect 497456 365502 497512 365536
rect 497546 365502 497602 365536
rect 497636 365502 497692 365536
rect 497726 365502 497782 365536
rect 497816 365502 497872 365536
rect 497906 365502 497962 365536
rect 497996 365502 498052 365536
rect 498086 365502 498142 365536
rect 498176 365502 498289 365536
rect 497327 365483 498289 365502
rect 497327 365086 498289 365105
rect 497327 365052 497403 365086
rect 497437 365052 497493 365086
rect 497527 365052 497583 365086
rect 497617 365052 497673 365086
rect 497707 365052 497763 365086
rect 497797 365052 497853 365086
rect 497887 365052 497943 365086
rect 497977 365052 498033 365086
rect 498067 365052 498123 365086
rect 498157 365052 498289 365086
rect 497327 365033 498289 365052
rect 497327 364974 497399 365033
rect 497327 364940 497346 364974
rect 497380 364940 497399 364974
rect 498217 365008 498289 365033
rect 498217 364974 498236 365008
rect 498270 364974 498289 365008
rect 497327 364884 497399 364940
rect 497327 364850 497346 364884
rect 497380 364850 497399 364884
rect 497327 364794 497399 364850
rect 497327 364760 497346 364794
rect 497380 364760 497399 364794
rect 497327 364704 497399 364760
rect 497327 364670 497346 364704
rect 497380 364670 497399 364704
rect 497327 364614 497399 364670
rect 497327 364580 497346 364614
rect 497380 364580 497399 364614
rect 497327 364524 497399 364580
rect 497327 364490 497346 364524
rect 497380 364490 497399 364524
rect 497327 364434 497399 364490
rect 497327 364400 497346 364434
rect 497380 364400 497399 364434
rect 497327 364344 497399 364400
rect 497327 364310 497346 364344
rect 497380 364310 497399 364344
rect 497327 364254 497399 364310
rect 498217 364918 498289 364974
rect 498217 364884 498236 364918
rect 498270 364884 498289 364918
rect 498217 364828 498289 364884
rect 498217 364794 498236 364828
rect 498270 364794 498289 364828
rect 498217 364738 498289 364794
rect 498217 364704 498236 364738
rect 498270 364704 498289 364738
rect 498217 364648 498289 364704
rect 498217 364614 498236 364648
rect 498270 364614 498289 364648
rect 498217 364558 498289 364614
rect 498217 364524 498236 364558
rect 498270 364524 498289 364558
rect 498217 364468 498289 364524
rect 498217 364434 498236 364468
rect 498270 364434 498289 364468
rect 498217 364378 498289 364434
rect 498217 364344 498236 364378
rect 498270 364344 498289 364378
rect 498217 364288 498289 364344
rect 497327 364220 497346 364254
rect 497380 364220 497399 364254
rect 497327 364215 497399 364220
rect 498217 364254 498236 364288
rect 498270 364254 498289 364288
rect 498217 364215 498289 364254
rect 497327 364196 498289 364215
rect 497327 364162 497422 364196
rect 497456 364162 497512 364196
rect 497546 364162 497602 364196
rect 497636 364162 497692 364196
rect 497726 364162 497782 364196
rect 497816 364162 497872 364196
rect 497906 364162 497962 364196
rect 497996 364162 498052 364196
rect 498086 364162 498142 364196
rect 498176 364162 498289 364196
rect 497327 364143 498289 364162
rect 497327 363746 498289 363765
rect 497327 363712 497403 363746
rect 497437 363712 497493 363746
rect 497527 363712 497583 363746
rect 497617 363712 497673 363746
rect 497707 363712 497763 363746
rect 497797 363712 497853 363746
rect 497887 363712 497943 363746
rect 497977 363712 498033 363746
rect 498067 363712 498123 363746
rect 498157 363712 498289 363746
rect 497327 363693 498289 363712
rect 497327 363634 497399 363693
rect 497327 363600 497346 363634
rect 497380 363600 497399 363634
rect 498217 363668 498289 363693
rect 498217 363634 498236 363668
rect 498270 363634 498289 363668
rect 497327 363544 497399 363600
rect 497327 363510 497346 363544
rect 497380 363510 497399 363544
rect 497327 363454 497399 363510
rect 497327 363420 497346 363454
rect 497380 363420 497399 363454
rect 497327 363364 497399 363420
rect 497327 363330 497346 363364
rect 497380 363330 497399 363364
rect 497327 363274 497399 363330
rect 497327 363240 497346 363274
rect 497380 363240 497399 363274
rect 497327 363184 497399 363240
rect 497327 363150 497346 363184
rect 497380 363150 497399 363184
rect 497327 363094 497399 363150
rect 497327 363060 497346 363094
rect 497380 363060 497399 363094
rect 497327 363004 497399 363060
rect 497327 362970 497346 363004
rect 497380 362970 497399 363004
rect 497327 362914 497399 362970
rect 498217 363578 498289 363634
rect 498217 363544 498236 363578
rect 498270 363544 498289 363578
rect 498217 363488 498289 363544
rect 498217 363454 498236 363488
rect 498270 363454 498289 363488
rect 498217 363398 498289 363454
rect 498217 363364 498236 363398
rect 498270 363364 498289 363398
rect 498217 363308 498289 363364
rect 498217 363274 498236 363308
rect 498270 363274 498289 363308
rect 498217 363218 498289 363274
rect 498217 363184 498236 363218
rect 498270 363184 498289 363218
rect 498217 363128 498289 363184
rect 498217 363094 498236 363128
rect 498270 363094 498289 363128
rect 498217 363038 498289 363094
rect 498217 363004 498236 363038
rect 498270 363004 498289 363038
rect 498217 362948 498289 363004
rect 497327 362880 497346 362914
rect 497380 362880 497399 362914
rect 497327 362875 497399 362880
rect 498217 362914 498236 362948
rect 498270 362914 498289 362948
rect 498217 362875 498289 362914
rect 497327 362856 498289 362875
rect 497327 362822 497422 362856
rect 497456 362822 497512 362856
rect 497546 362822 497602 362856
rect 497636 362822 497692 362856
rect 497726 362822 497782 362856
rect 497816 362822 497872 362856
rect 497906 362822 497962 362856
rect 497996 362822 498052 362856
rect 498086 362822 498142 362856
rect 498176 362822 498289 362856
rect 497327 362803 498289 362822
rect 501087 371622 502049 371641
rect 501087 371588 501163 371622
rect 501197 371588 501253 371622
rect 501287 371588 501343 371622
rect 501377 371588 501433 371622
rect 501467 371588 501523 371622
rect 501557 371588 501613 371622
rect 501647 371588 501703 371622
rect 501737 371588 501793 371622
rect 501827 371588 501883 371622
rect 501917 371588 502049 371622
rect 501087 371569 502049 371588
rect 501087 371510 501159 371569
rect 501087 371476 501106 371510
rect 501140 371476 501159 371510
rect 501977 371544 502049 371569
rect 501977 371510 501996 371544
rect 502030 371510 502049 371544
rect 501087 371420 501159 371476
rect 501087 371386 501106 371420
rect 501140 371386 501159 371420
rect 501087 371330 501159 371386
rect 501087 371296 501106 371330
rect 501140 371296 501159 371330
rect 501087 371240 501159 371296
rect 501087 371206 501106 371240
rect 501140 371206 501159 371240
rect 501087 371150 501159 371206
rect 501087 371116 501106 371150
rect 501140 371116 501159 371150
rect 501087 371060 501159 371116
rect 501087 371026 501106 371060
rect 501140 371026 501159 371060
rect 501087 370970 501159 371026
rect 501087 370936 501106 370970
rect 501140 370936 501159 370970
rect 501087 370880 501159 370936
rect 501087 370846 501106 370880
rect 501140 370846 501159 370880
rect 501087 370790 501159 370846
rect 501977 371454 502049 371510
rect 501977 371420 501996 371454
rect 502030 371420 502049 371454
rect 501977 371364 502049 371420
rect 501977 371330 501996 371364
rect 502030 371330 502049 371364
rect 501977 371274 502049 371330
rect 501977 371240 501996 371274
rect 502030 371240 502049 371274
rect 501977 371184 502049 371240
rect 501977 371150 501996 371184
rect 502030 371150 502049 371184
rect 501977 371094 502049 371150
rect 501977 371060 501996 371094
rect 502030 371060 502049 371094
rect 501977 371004 502049 371060
rect 501977 370970 501996 371004
rect 502030 370970 502049 371004
rect 501977 370914 502049 370970
rect 501977 370880 501996 370914
rect 502030 370880 502049 370914
rect 501977 370824 502049 370880
rect 501087 370756 501106 370790
rect 501140 370756 501159 370790
rect 501087 370751 501159 370756
rect 501977 370790 501996 370824
rect 502030 370790 502049 370824
rect 501977 370751 502049 370790
rect 501087 370732 502049 370751
rect 501087 370698 501182 370732
rect 501216 370698 501272 370732
rect 501306 370698 501362 370732
rect 501396 370698 501452 370732
rect 501486 370698 501542 370732
rect 501576 370698 501632 370732
rect 501666 370698 501722 370732
rect 501756 370698 501812 370732
rect 501846 370698 501902 370732
rect 501936 370698 502049 370732
rect 501087 370679 502049 370698
rect 501087 370282 502049 370301
rect 501087 370248 501163 370282
rect 501197 370248 501253 370282
rect 501287 370248 501343 370282
rect 501377 370248 501433 370282
rect 501467 370248 501523 370282
rect 501557 370248 501613 370282
rect 501647 370248 501703 370282
rect 501737 370248 501793 370282
rect 501827 370248 501883 370282
rect 501917 370248 502049 370282
rect 501087 370229 502049 370248
rect 501087 370170 501159 370229
rect 501087 370136 501106 370170
rect 501140 370136 501159 370170
rect 501977 370204 502049 370229
rect 501977 370170 501996 370204
rect 502030 370170 502049 370204
rect 501087 370080 501159 370136
rect 501087 370046 501106 370080
rect 501140 370046 501159 370080
rect 501087 369990 501159 370046
rect 501087 369956 501106 369990
rect 501140 369956 501159 369990
rect 501087 369900 501159 369956
rect 501087 369866 501106 369900
rect 501140 369866 501159 369900
rect 501087 369810 501159 369866
rect 501087 369776 501106 369810
rect 501140 369776 501159 369810
rect 501087 369720 501159 369776
rect 501087 369686 501106 369720
rect 501140 369686 501159 369720
rect 501087 369630 501159 369686
rect 501087 369596 501106 369630
rect 501140 369596 501159 369630
rect 501087 369540 501159 369596
rect 501087 369506 501106 369540
rect 501140 369506 501159 369540
rect 501087 369450 501159 369506
rect 501977 370114 502049 370170
rect 501977 370080 501996 370114
rect 502030 370080 502049 370114
rect 501977 370024 502049 370080
rect 501977 369990 501996 370024
rect 502030 369990 502049 370024
rect 501977 369934 502049 369990
rect 501977 369900 501996 369934
rect 502030 369900 502049 369934
rect 501977 369844 502049 369900
rect 501977 369810 501996 369844
rect 502030 369810 502049 369844
rect 501977 369754 502049 369810
rect 501977 369720 501996 369754
rect 502030 369720 502049 369754
rect 501977 369664 502049 369720
rect 501977 369630 501996 369664
rect 502030 369630 502049 369664
rect 501977 369574 502049 369630
rect 501977 369540 501996 369574
rect 502030 369540 502049 369574
rect 501977 369484 502049 369540
rect 501087 369416 501106 369450
rect 501140 369416 501159 369450
rect 501087 369411 501159 369416
rect 501977 369450 501996 369484
rect 502030 369450 502049 369484
rect 501977 369411 502049 369450
rect 501087 369392 502049 369411
rect 501087 369358 501182 369392
rect 501216 369358 501272 369392
rect 501306 369358 501362 369392
rect 501396 369358 501452 369392
rect 501486 369358 501542 369392
rect 501576 369358 501632 369392
rect 501666 369358 501722 369392
rect 501756 369358 501812 369392
rect 501846 369358 501902 369392
rect 501936 369358 502049 369392
rect 501087 369339 502049 369358
rect 501087 368942 502049 368961
rect 501087 368908 501163 368942
rect 501197 368908 501253 368942
rect 501287 368908 501343 368942
rect 501377 368908 501433 368942
rect 501467 368908 501523 368942
rect 501557 368908 501613 368942
rect 501647 368908 501703 368942
rect 501737 368908 501793 368942
rect 501827 368908 501883 368942
rect 501917 368908 502049 368942
rect 501087 368889 502049 368908
rect 501087 368830 501159 368889
rect 501087 368796 501106 368830
rect 501140 368796 501159 368830
rect 501977 368864 502049 368889
rect 501977 368830 501996 368864
rect 502030 368830 502049 368864
rect 501087 368740 501159 368796
rect 501087 368706 501106 368740
rect 501140 368706 501159 368740
rect 501087 368650 501159 368706
rect 501087 368616 501106 368650
rect 501140 368616 501159 368650
rect 501087 368560 501159 368616
rect 501087 368526 501106 368560
rect 501140 368526 501159 368560
rect 501087 368470 501159 368526
rect 501087 368436 501106 368470
rect 501140 368436 501159 368470
rect 501087 368380 501159 368436
rect 501087 368346 501106 368380
rect 501140 368346 501159 368380
rect 501087 368290 501159 368346
rect 501087 368256 501106 368290
rect 501140 368256 501159 368290
rect 501087 368200 501159 368256
rect 501087 368166 501106 368200
rect 501140 368166 501159 368200
rect 501087 368110 501159 368166
rect 501977 368774 502049 368830
rect 501977 368740 501996 368774
rect 502030 368740 502049 368774
rect 501977 368684 502049 368740
rect 501977 368650 501996 368684
rect 502030 368650 502049 368684
rect 501977 368594 502049 368650
rect 501977 368560 501996 368594
rect 502030 368560 502049 368594
rect 501977 368504 502049 368560
rect 501977 368470 501996 368504
rect 502030 368470 502049 368504
rect 501977 368414 502049 368470
rect 501977 368380 501996 368414
rect 502030 368380 502049 368414
rect 501977 368324 502049 368380
rect 501977 368290 501996 368324
rect 502030 368290 502049 368324
rect 501977 368234 502049 368290
rect 501977 368200 501996 368234
rect 502030 368200 502049 368234
rect 501977 368144 502049 368200
rect 501087 368076 501106 368110
rect 501140 368076 501159 368110
rect 501087 368071 501159 368076
rect 501977 368110 501996 368144
rect 502030 368110 502049 368144
rect 501977 368071 502049 368110
rect 501087 368052 502049 368071
rect 501087 368018 501182 368052
rect 501216 368018 501272 368052
rect 501306 368018 501362 368052
rect 501396 368018 501452 368052
rect 501486 368018 501542 368052
rect 501576 368018 501632 368052
rect 501666 368018 501722 368052
rect 501756 368018 501812 368052
rect 501846 368018 501902 368052
rect 501936 368018 502049 368052
rect 501087 367999 502049 368018
rect 501087 367602 502049 367621
rect 501087 367568 501163 367602
rect 501197 367568 501253 367602
rect 501287 367568 501343 367602
rect 501377 367568 501433 367602
rect 501467 367568 501523 367602
rect 501557 367568 501613 367602
rect 501647 367568 501703 367602
rect 501737 367568 501793 367602
rect 501827 367568 501883 367602
rect 501917 367568 502049 367602
rect 501087 367549 502049 367568
rect 501087 367490 501159 367549
rect 501087 367456 501106 367490
rect 501140 367456 501159 367490
rect 501977 367524 502049 367549
rect 501977 367490 501996 367524
rect 502030 367490 502049 367524
rect 501087 367400 501159 367456
rect 501087 367366 501106 367400
rect 501140 367366 501159 367400
rect 501087 367310 501159 367366
rect 501087 367276 501106 367310
rect 501140 367276 501159 367310
rect 501087 367220 501159 367276
rect 501087 367186 501106 367220
rect 501140 367186 501159 367220
rect 501087 367130 501159 367186
rect 501087 367096 501106 367130
rect 501140 367096 501159 367130
rect 501087 367040 501159 367096
rect 501087 367006 501106 367040
rect 501140 367006 501159 367040
rect 501087 366950 501159 367006
rect 501087 366916 501106 366950
rect 501140 366916 501159 366950
rect 501087 366860 501159 366916
rect 501087 366826 501106 366860
rect 501140 366826 501159 366860
rect 501087 366770 501159 366826
rect 501977 367434 502049 367490
rect 501977 367400 501996 367434
rect 502030 367400 502049 367434
rect 501977 367344 502049 367400
rect 501977 367310 501996 367344
rect 502030 367310 502049 367344
rect 501977 367254 502049 367310
rect 501977 367220 501996 367254
rect 502030 367220 502049 367254
rect 501977 367164 502049 367220
rect 501977 367130 501996 367164
rect 502030 367130 502049 367164
rect 501977 367074 502049 367130
rect 501977 367040 501996 367074
rect 502030 367040 502049 367074
rect 501977 366984 502049 367040
rect 501977 366950 501996 366984
rect 502030 366950 502049 366984
rect 501977 366894 502049 366950
rect 501977 366860 501996 366894
rect 502030 366860 502049 366894
rect 501977 366804 502049 366860
rect 501087 366736 501106 366770
rect 501140 366736 501159 366770
rect 501087 366731 501159 366736
rect 501977 366770 501996 366804
rect 502030 366770 502049 366804
rect 501977 366731 502049 366770
rect 501087 366712 502049 366731
rect 501087 366678 501182 366712
rect 501216 366678 501272 366712
rect 501306 366678 501362 366712
rect 501396 366678 501452 366712
rect 501486 366678 501542 366712
rect 501576 366678 501632 366712
rect 501666 366678 501722 366712
rect 501756 366678 501812 366712
rect 501846 366678 501902 366712
rect 501936 366678 502049 366712
rect 501087 366659 502049 366678
rect 501087 366262 502049 366281
rect 501087 366228 501163 366262
rect 501197 366228 501253 366262
rect 501287 366228 501343 366262
rect 501377 366228 501433 366262
rect 501467 366228 501523 366262
rect 501557 366228 501613 366262
rect 501647 366228 501703 366262
rect 501737 366228 501793 366262
rect 501827 366228 501883 366262
rect 501917 366228 502049 366262
rect 501087 366209 502049 366228
rect 501087 366150 501159 366209
rect 501087 366116 501106 366150
rect 501140 366116 501159 366150
rect 501977 366184 502049 366209
rect 501977 366150 501996 366184
rect 502030 366150 502049 366184
rect 501087 366060 501159 366116
rect 501087 366026 501106 366060
rect 501140 366026 501159 366060
rect 501087 365970 501159 366026
rect 501087 365936 501106 365970
rect 501140 365936 501159 365970
rect 501087 365880 501159 365936
rect 501087 365846 501106 365880
rect 501140 365846 501159 365880
rect 501087 365790 501159 365846
rect 501087 365756 501106 365790
rect 501140 365756 501159 365790
rect 501087 365700 501159 365756
rect 501087 365666 501106 365700
rect 501140 365666 501159 365700
rect 501087 365610 501159 365666
rect 501087 365576 501106 365610
rect 501140 365576 501159 365610
rect 501087 365520 501159 365576
rect 501087 365486 501106 365520
rect 501140 365486 501159 365520
rect 501087 365430 501159 365486
rect 501977 366094 502049 366150
rect 501977 366060 501996 366094
rect 502030 366060 502049 366094
rect 501977 366004 502049 366060
rect 501977 365970 501996 366004
rect 502030 365970 502049 366004
rect 501977 365914 502049 365970
rect 501977 365880 501996 365914
rect 502030 365880 502049 365914
rect 501977 365824 502049 365880
rect 501977 365790 501996 365824
rect 502030 365790 502049 365824
rect 501977 365734 502049 365790
rect 501977 365700 501996 365734
rect 502030 365700 502049 365734
rect 501977 365644 502049 365700
rect 501977 365610 501996 365644
rect 502030 365610 502049 365644
rect 501977 365554 502049 365610
rect 501977 365520 501996 365554
rect 502030 365520 502049 365554
rect 501977 365464 502049 365520
rect 501087 365396 501106 365430
rect 501140 365396 501159 365430
rect 501087 365391 501159 365396
rect 501977 365430 501996 365464
rect 502030 365430 502049 365464
rect 501977 365391 502049 365430
rect 501087 365372 502049 365391
rect 501087 365338 501182 365372
rect 501216 365338 501272 365372
rect 501306 365338 501362 365372
rect 501396 365338 501452 365372
rect 501486 365338 501542 365372
rect 501576 365338 501632 365372
rect 501666 365338 501722 365372
rect 501756 365338 501812 365372
rect 501846 365338 501902 365372
rect 501936 365338 502049 365372
rect 501087 365319 502049 365338
rect 501087 364922 502049 364941
rect 501087 364888 501163 364922
rect 501197 364888 501253 364922
rect 501287 364888 501343 364922
rect 501377 364888 501433 364922
rect 501467 364888 501523 364922
rect 501557 364888 501613 364922
rect 501647 364888 501703 364922
rect 501737 364888 501793 364922
rect 501827 364888 501883 364922
rect 501917 364888 502049 364922
rect 501087 364869 502049 364888
rect 501087 364810 501159 364869
rect 501087 364776 501106 364810
rect 501140 364776 501159 364810
rect 501977 364844 502049 364869
rect 501977 364810 501996 364844
rect 502030 364810 502049 364844
rect 501087 364720 501159 364776
rect 501087 364686 501106 364720
rect 501140 364686 501159 364720
rect 501087 364630 501159 364686
rect 501087 364596 501106 364630
rect 501140 364596 501159 364630
rect 501087 364540 501159 364596
rect 501087 364506 501106 364540
rect 501140 364506 501159 364540
rect 501087 364450 501159 364506
rect 501087 364416 501106 364450
rect 501140 364416 501159 364450
rect 501087 364360 501159 364416
rect 501087 364326 501106 364360
rect 501140 364326 501159 364360
rect 501087 364270 501159 364326
rect 501087 364236 501106 364270
rect 501140 364236 501159 364270
rect 501087 364180 501159 364236
rect 501087 364146 501106 364180
rect 501140 364146 501159 364180
rect 501087 364090 501159 364146
rect 501977 364754 502049 364810
rect 501977 364720 501996 364754
rect 502030 364720 502049 364754
rect 501977 364664 502049 364720
rect 501977 364630 501996 364664
rect 502030 364630 502049 364664
rect 501977 364574 502049 364630
rect 501977 364540 501996 364574
rect 502030 364540 502049 364574
rect 501977 364484 502049 364540
rect 501977 364450 501996 364484
rect 502030 364450 502049 364484
rect 501977 364394 502049 364450
rect 501977 364360 501996 364394
rect 502030 364360 502049 364394
rect 501977 364304 502049 364360
rect 501977 364270 501996 364304
rect 502030 364270 502049 364304
rect 501977 364214 502049 364270
rect 501977 364180 501996 364214
rect 502030 364180 502049 364214
rect 501977 364124 502049 364180
rect 501087 364056 501106 364090
rect 501140 364056 501159 364090
rect 501087 364051 501159 364056
rect 501977 364090 501996 364124
rect 502030 364090 502049 364124
rect 501977 364051 502049 364090
rect 501087 364032 502049 364051
rect 501087 363998 501182 364032
rect 501216 363998 501272 364032
rect 501306 363998 501362 364032
rect 501396 363998 501452 364032
rect 501486 363998 501542 364032
rect 501576 363998 501632 364032
rect 501666 363998 501722 364032
rect 501756 363998 501812 364032
rect 501846 363998 501902 364032
rect 501936 363998 502049 364032
rect 501087 363979 502049 363998
rect 501087 363582 502049 363601
rect 501087 363548 501163 363582
rect 501197 363548 501253 363582
rect 501287 363548 501343 363582
rect 501377 363548 501433 363582
rect 501467 363548 501523 363582
rect 501557 363548 501613 363582
rect 501647 363548 501703 363582
rect 501737 363548 501793 363582
rect 501827 363548 501883 363582
rect 501917 363548 502049 363582
rect 501087 363529 502049 363548
rect 501087 363470 501159 363529
rect 501087 363436 501106 363470
rect 501140 363436 501159 363470
rect 501977 363504 502049 363529
rect 501977 363470 501996 363504
rect 502030 363470 502049 363504
rect 501087 363380 501159 363436
rect 501087 363346 501106 363380
rect 501140 363346 501159 363380
rect 501087 363290 501159 363346
rect 501087 363256 501106 363290
rect 501140 363256 501159 363290
rect 501087 363200 501159 363256
rect 501087 363166 501106 363200
rect 501140 363166 501159 363200
rect 501087 363110 501159 363166
rect 501087 363076 501106 363110
rect 501140 363076 501159 363110
rect 501087 363020 501159 363076
rect 501087 362986 501106 363020
rect 501140 362986 501159 363020
rect 501087 362930 501159 362986
rect 501087 362896 501106 362930
rect 501140 362896 501159 362930
rect 501087 362840 501159 362896
rect 501087 362806 501106 362840
rect 501140 362806 501159 362840
rect 501087 362750 501159 362806
rect 501977 363414 502049 363470
rect 501977 363380 501996 363414
rect 502030 363380 502049 363414
rect 501977 363324 502049 363380
rect 501977 363290 501996 363324
rect 502030 363290 502049 363324
rect 501977 363234 502049 363290
rect 501977 363200 501996 363234
rect 502030 363200 502049 363234
rect 501977 363144 502049 363200
rect 501977 363110 501996 363144
rect 502030 363110 502049 363144
rect 501977 363054 502049 363110
rect 501977 363020 501996 363054
rect 502030 363020 502049 363054
rect 501977 362964 502049 363020
rect 501977 362930 501996 362964
rect 502030 362930 502049 362964
rect 501977 362874 502049 362930
rect 501977 362840 501996 362874
rect 502030 362840 502049 362874
rect 501977 362784 502049 362840
rect 501087 362716 501106 362750
rect 501140 362716 501159 362750
rect 501087 362711 501159 362716
rect 501977 362750 501996 362784
rect 502030 362750 502049 362784
rect 501977 362711 502049 362750
rect 501087 362692 502049 362711
rect 501087 362658 501182 362692
rect 501216 362658 501272 362692
rect 501306 362658 501362 362692
rect 501396 362658 501452 362692
rect 501486 362658 501542 362692
rect 501576 362658 501632 362692
rect 501666 362658 501722 362692
rect 501756 362658 501812 362692
rect 501846 362658 501902 362692
rect 501936 362658 502049 362692
rect 501087 362639 502049 362658
rect 504847 372962 505809 372981
rect 504847 372928 504923 372962
rect 504957 372928 505013 372962
rect 505047 372928 505103 372962
rect 505137 372928 505193 372962
rect 505227 372928 505283 372962
rect 505317 372928 505373 372962
rect 505407 372928 505463 372962
rect 505497 372928 505553 372962
rect 505587 372928 505643 372962
rect 505677 372928 505809 372962
rect 504847 372909 505809 372928
rect 504847 372850 504919 372909
rect 504847 372816 504866 372850
rect 504900 372816 504919 372850
rect 505737 372884 505809 372909
rect 505737 372850 505756 372884
rect 505790 372850 505809 372884
rect 504847 372760 504919 372816
rect 504847 372726 504866 372760
rect 504900 372726 504919 372760
rect 504847 372670 504919 372726
rect 504847 372636 504866 372670
rect 504900 372636 504919 372670
rect 504847 372580 504919 372636
rect 504847 372546 504866 372580
rect 504900 372546 504919 372580
rect 504847 372490 504919 372546
rect 504847 372456 504866 372490
rect 504900 372456 504919 372490
rect 504847 372400 504919 372456
rect 504847 372366 504866 372400
rect 504900 372366 504919 372400
rect 504847 372310 504919 372366
rect 504847 372276 504866 372310
rect 504900 372276 504919 372310
rect 504847 372220 504919 372276
rect 504847 372186 504866 372220
rect 504900 372186 504919 372220
rect 504847 372130 504919 372186
rect 505737 372794 505809 372850
rect 505737 372760 505756 372794
rect 505790 372760 505809 372794
rect 505737 372704 505809 372760
rect 505737 372670 505756 372704
rect 505790 372670 505809 372704
rect 505737 372614 505809 372670
rect 505737 372580 505756 372614
rect 505790 372580 505809 372614
rect 505737 372524 505809 372580
rect 505737 372490 505756 372524
rect 505790 372490 505809 372524
rect 505737 372434 505809 372490
rect 505737 372400 505756 372434
rect 505790 372400 505809 372434
rect 505737 372344 505809 372400
rect 505737 372310 505756 372344
rect 505790 372310 505809 372344
rect 505737 372254 505809 372310
rect 505737 372220 505756 372254
rect 505790 372220 505809 372254
rect 505737 372164 505809 372220
rect 504847 372096 504866 372130
rect 504900 372096 504919 372130
rect 504847 372091 504919 372096
rect 505737 372130 505756 372164
rect 505790 372130 505809 372164
rect 505737 372091 505809 372130
rect 504847 372072 505809 372091
rect 504847 372038 504942 372072
rect 504976 372038 505032 372072
rect 505066 372038 505122 372072
rect 505156 372038 505212 372072
rect 505246 372038 505302 372072
rect 505336 372038 505392 372072
rect 505426 372038 505482 372072
rect 505516 372038 505572 372072
rect 505606 372038 505662 372072
rect 505696 372038 505809 372072
rect 504847 372019 505809 372038
rect 504847 371622 505809 371641
rect 504847 371588 504923 371622
rect 504957 371588 505013 371622
rect 505047 371588 505103 371622
rect 505137 371588 505193 371622
rect 505227 371588 505283 371622
rect 505317 371588 505373 371622
rect 505407 371588 505463 371622
rect 505497 371588 505553 371622
rect 505587 371588 505643 371622
rect 505677 371588 505809 371622
rect 504847 371569 505809 371588
rect 504847 371510 504919 371569
rect 504847 371476 504866 371510
rect 504900 371476 504919 371510
rect 505737 371544 505809 371569
rect 505737 371510 505756 371544
rect 505790 371510 505809 371544
rect 504847 371420 504919 371476
rect 504847 371386 504866 371420
rect 504900 371386 504919 371420
rect 504847 371330 504919 371386
rect 504847 371296 504866 371330
rect 504900 371296 504919 371330
rect 504847 371240 504919 371296
rect 504847 371206 504866 371240
rect 504900 371206 504919 371240
rect 504847 371150 504919 371206
rect 504847 371116 504866 371150
rect 504900 371116 504919 371150
rect 504847 371060 504919 371116
rect 504847 371026 504866 371060
rect 504900 371026 504919 371060
rect 504847 370970 504919 371026
rect 504847 370936 504866 370970
rect 504900 370936 504919 370970
rect 504847 370880 504919 370936
rect 504847 370846 504866 370880
rect 504900 370846 504919 370880
rect 504847 370790 504919 370846
rect 505737 371454 505809 371510
rect 505737 371420 505756 371454
rect 505790 371420 505809 371454
rect 505737 371364 505809 371420
rect 505737 371330 505756 371364
rect 505790 371330 505809 371364
rect 505737 371274 505809 371330
rect 505737 371240 505756 371274
rect 505790 371240 505809 371274
rect 505737 371184 505809 371240
rect 505737 371150 505756 371184
rect 505790 371150 505809 371184
rect 505737 371094 505809 371150
rect 505737 371060 505756 371094
rect 505790 371060 505809 371094
rect 505737 371004 505809 371060
rect 505737 370970 505756 371004
rect 505790 370970 505809 371004
rect 505737 370914 505809 370970
rect 505737 370880 505756 370914
rect 505790 370880 505809 370914
rect 505737 370824 505809 370880
rect 504847 370756 504866 370790
rect 504900 370756 504919 370790
rect 504847 370751 504919 370756
rect 505737 370790 505756 370824
rect 505790 370790 505809 370824
rect 505737 370751 505809 370790
rect 504847 370732 505809 370751
rect 504847 370698 504942 370732
rect 504976 370698 505032 370732
rect 505066 370698 505122 370732
rect 505156 370698 505212 370732
rect 505246 370698 505302 370732
rect 505336 370698 505392 370732
rect 505426 370698 505482 370732
rect 505516 370698 505572 370732
rect 505606 370698 505662 370732
rect 505696 370698 505809 370732
rect 504847 370679 505809 370698
rect 504847 370282 505809 370301
rect 504847 370248 504923 370282
rect 504957 370248 505013 370282
rect 505047 370248 505103 370282
rect 505137 370248 505193 370282
rect 505227 370248 505283 370282
rect 505317 370248 505373 370282
rect 505407 370248 505463 370282
rect 505497 370248 505553 370282
rect 505587 370248 505643 370282
rect 505677 370248 505809 370282
rect 504847 370229 505809 370248
rect 504847 370170 504919 370229
rect 504847 370136 504866 370170
rect 504900 370136 504919 370170
rect 505737 370204 505809 370229
rect 505737 370170 505756 370204
rect 505790 370170 505809 370204
rect 504847 370080 504919 370136
rect 504847 370046 504866 370080
rect 504900 370046 504919 370080
rect 504847 369990 504919 370046
rect 504847 369956 504866 369990
rect 504900 369956 504919 369990
rect 504847 369900 504919 369956
rect 504847 369866 504866 369900
rect 504900 369866 504919 369900
rect 504847 369810 504919 369866
rect 504847 369776 504866 369810
rect 504900 369776 504919 369810
rect 504847 369720 504919 369776
rect 504847 369686 504866 369720
rect 504900 369686 504919 369720
rect 504847 369630 504919 369686
rect 504847 369596 504866 369630
rect 504900 369596 504919 369630
rect 504847 369540 504919 369596
rect 504847 369506 504866 369540
rect 504900 369506 504919 369540
rect 504847 369450 504919 369506
rect 505737 370114 505809 370170
rect 505737 370080 505756 370114
rect 505790 370080 505809 370114
rect 505737 370024 505809 370080
rect 505737 369990 505756 370024
rect 505790 369990 505809 370024
rect 505737 369934 505809 369990
rect 505737 369900 505756 369934
rect 505790 369900 505809 369934
rect 505737 369844 505809 369900
rect 505737 369810 505756 369844
rect 505790 369810 505809 369844
rect 505737 369754 505809 369810
rect 505737 369720 505756 369754
rect 505790 369720 505809 369754
rect 505737 369664 505809 369720
rect 505737 369630 505756 369664
rect 505790 369630 505809 369664
rect 505737 369574 505809 369630
rect 505737 369540 505756 369574
rect 505790 369540 505809 369574
rect 505737 369484 505809 369540
rect 504847 369416 504866 369450
rect 504900 369416 504919 369450
rect 504847 369411 504919 369416
rect 505737 369450 505756 369484
rect 505790 369450 505809 369484
rect 505737 369411 505809 369450
rect 504847 369392 505809 369411
rect 504847 369358 504942 369392
rect 504976 369358 505032 369392
rect 505066 369358 505122 369392
rect 505156 369358 505212 369392
rect 505246 369358 505302 369392
rect 505336 369358 505392 369392
rect 505426 369358 505482 369392
rect 505516 369358 505572 369392
rect 505606 369358 505662 369392
rect 505696 369358 505809 369392
rect 504847 369339 505809 369358
rect 504847 368942 505809 368961
rect 504847 368908 504923 368942
rect 504957 368908 505013 368942
rect 505047 368908 505103 368942
rect 505137 368908 505193 368942
rect 505227 368908 505283 368942
rect 505317 368908 505373 368942
rect 505407 368908 505463 368942
rect 505497 368908 505553 368942
rect 505587 368908 505643 368942
rect 505677 368908 505809 368942
rect 504847 368889 505809 368908
rect 504847 368830 504919 368889
rect 504847 368796 504866 368830
rect 504900 368796 504919 368830
rect 505737 368864 505809 368889
rect 505737 368830 505756 368864
rect 505790 368830 505809 368864
rect 504847 368740 504919 368796
rect 504847 368706 504866 368740
rect 504900 368706 504919 368740
rect 504847 368650 504919 368706
rect 504847 368616 504866 368650
rect 504900 368616 504919 368650
rect 504847 368560 504919 368616
rect 504847 368526 504866 368560
rect 504900 368526 504919 368560
rect 504847 368470 504919 368526
rect 504847 368436 504866 368470
rect 504900 368436 504919 368470
rect 504847 368380 504919 368436
rect 504847 368346 504866 368380
rect 504900 368346 504919 368380
rect 504847 368290 504919 368346
rect 504847 368256 504866 368290
rect 504900 368256 504919 368290
rect 504847 368200 504919 368256
rect 504847 368166 504866 368200
rect 504900 368166 504919 368200
rect 504847 368110 504919 368166
rect 505737 368774 505809 368830
rect 505737 368740 505756 368774
rect 505790 368740 505809 368774
rect 505737 368684 505809 368740
rect 505737 368650 505756 368684
rect 505790 368650 505809 368684
rect 505737 368594 505809 368650
rect 505737 368560 505756 368594
rect 505790 368560 505809 368594
rect 505737 368504 505809 368560
rect 505737 368470 505756 368504
rect 505790 368470 505809 368504
rect 505737 368414 505809 368470
rect 505737 368380 505756 368414
rect 505790 368380 505809 368414
rect 505737 368324 505809 368380
rect 505737 368290 505756 368324
rect 505790 368290 505809 368324
rect 505737 368234 505809 368290
rect 505737 368200 505756 368234
rect 505790 368200 505809 368234
rect 505737 368144 505809 368200
rect 504847 368076 504866 368110
rect 504900 368076 504919 368110
rect 504847 368071 504919 368076
rect 505737 368110 505756 368144
rect 505790 368110 505809 368144
rect 505737 368071 505809 368110
rect 504847 368052 505809 368071
rect 504847 368018 504942 368052
rect 504976 368018 505032 368052
rect 505066 368018 505122 368052
rect 505156 368018 505212 368052
rect 505246 368018 505302 368052
rect 505336 368018 505392 368052
rect 505426 368018 505482 368052
rect 505516 368018 505572 368052
rect 505606 368018 505662 368052
rect 505696 368018 505809 368052
rect 504847 367999 505809 368018
rect 504847 367602 505809 367621
rect 504847 367568 504923 367602
rect 504957 367568 505013 367602
rect 505047 367568 505103 367602
rect 505137 367568 505193 367602
rect 505227 367568 505283 367602
rect 505317 367568 505373 367602
rect 505407 367568 505463 367602
rect 505497 367568 505553 367602
rect 505587 367568 505643 367602
rect 505677 367568 505809 367602
rect 504847 367549 505809 367568
rect 504847 367490 504919 367549
rect 504847 367456 504866 367490
rect 504900 367456 504919 367490
rect 505737 367524 505809 367549
rect 505737 367490 505756 367524
rect 505790 367490 505809 367524
rect 504847 367400 504919 367456
rect 504847 367366 504866 367400
rect 504900 367366 504919 367400
rect 504847 367310 504919 367366
rect 504847 367276 504866 367310
rect 504900 367276 504919 367310
rect 504847 367220 504919 367276
rect 504847 367186 504866 367220
rect 504900 367186 504919 367220
rect 504847 367130 504919 367186
rect 504847 367096 504866 367130
rect 504900 367096 504919 367130
rect 504847 367040 504919 367096
rect 504847 367006 504866 367040
rect 504900 367006 504919 367040
rect 504847 366950 504919 367006
rect 504847 366916 504866 366950
rect 504900 366916 504919 366950
rect 504847 366860 504919 366916
rect 504847 366826 504866 366860
rect 504900 366826 504919 366860
rect 504847 366770 504919 366826
rect 505737 367434 505809 367490
rect 505737 367400 505756 367434
rect 505790 367400 505809 367434
rect 505737 367344 505809 367400
rect 505737 367310 505756 367344
rect 505790 367310 505809 367344
rect 505737 367254 505809 367310
rect 505737 367220 505756 367254
rect 505790 367220 505809 367254
rect 505737 367164 505809 367220
rect 505737 367130 505756 367164
rect 505790 367130 505809 367164
rect 505737 367074 505809 367130
rect 505737 367040 505756 367074
rect 505790 367040 505809 367074
rect 505737 366984 505809 367040
rect 505737 366950 505756 366984
rect 505790 366950 505809 366984
rect 505737 366894 505809 366950
rect 505737 366860 505756 366894
rect 505790 366860 505809 366894
rect 505737 366804 505809 366860
rect 504847 366736 504866 366770
rect 504900 366736 504919 366770
rect 504847 366731 504919 366736
rect 505737 366770 505756 366804
rect 505790 366770 505809 366804
rect 505737 366731 505809 366770
rect 504847 366712 505809 366731
rect 504847 366678 504942 366712
rect 504976 366678 505032 366712
rect 505066 366678 505122 366712
rect 505156 366678 505212 366712
rect 505246 366678 505302 366712
rect 505336 366678 505392 366712
rect 505426 366678 505482 366712
rect 505516 366678 505572 366712
rect 505606 366678 505662 366712
rect 505696 366678 505809 366712
rect 504847 366659 505809 366678
rect 504847 366262 505809 366281
rect 504847 366228 504923 366262
rect 504957 366228 505013 366262
rect 505047 366228 505103 366262
rect 505137 366228 505193 366262
rect 505227 366228 505283 366262
rect 505317 366228 505373 366262
rect 505407 366228 505463 366262
rect 505497 366228 505553 366262
rect 505587 366228 505643 366262
rect 505677 366228 505809 366262
rect 504847 366209 505809 366228
rect 504847 366150 504919 366209
rect 504847 366116 504866 366150
rect 504900 366116 504919 366150
rect 505737 366184 505809 366209
rect 505737 366150 505756 366184
rect 505790 366150 505809 366184
rect 504847 366060 504919 366116
rect 504847 366026 504866 366060
rect 504900 366026 504919 366060
rect 504847 365970 504919 366026
rect 504847 365936 504866 365970
rect 504900 365936 504919 365970
rect 504847 365880 504919 365936
rect 504847 365846 504866 365880
rect 504900 365846 504919 365880
rect 504847 365790 504919 365846
rect 504847 365756 504866 365790
rect 504900 365756 504919 365790
rect 504847 365700 504919 365756
rect 504847 365666 504866 365700
rect 504900 365666 504919 365700
rect 504847 365610 504919 365666
rect 504847 365576 504866 365610
rect 504900 365576 504919 365610
rect 504847 365520 504919 365576
rect 504847 365486 504866 365520
rect 504900 365486 504919 365520
rect 504847 365430 504919 365486
rect 505737 366094 505809 366150
rect 505737 366060 505756 366094
rect 505790 366060 505809 366094
rect 505737 366004 505809 366060
rect 505737 365970 505756 366004
rect 505790 365970 505809 366004
rect 505737 365914 505809 365970
rect 505737 365880 505756 365914
rect 505790 365880 505809 365914
rect 505737 365824 505809 365880
rect 505737 365790 505756 365824
rect 505790 365790 505809 365824
rect 505737 365734 505809 365790
rect 505737 365700 505756 365734
rect 505790 365700 505809 365734
rect 505737 365644 505809 365700
rect 505737 365610 505756 365644
rect 505790 365610 505809 365644
rect 505737 365554 505809 365610
rect 505737 365520 505756 365554
rect 505790 365520 505809 365554
rect 505737 365464 505809 365520
rect 504847 365396 504866 365430
rect 504900 365396 504919 365430
rect 504847 365391 504919 365396
rect 505737 365430 505756 365464
rect 505790 365430 505809 365464
rect 505737 365391 505809 365430
rect 504847 365372 505809 365391
rect 504847 365338 504942 365372
rect 504976 365338 505032 365372
rect 505066 365338 505122 365372
rect 505156 365338 505212 365372
rect 505246 365338 505302 365372
rect 505336 365338 505392 365372
rect 505426 365338 505482 365372
rect 505516 365338 505572 365372
rect 505606 365338 505662 365372
rect 505696 365338 505809 365372
rect 504847 365319 505809 365338
rect 504847 364922 505809 364941
rect 504847 364888 504923 364922
rect 504957 364888 505013 364922
rect 505047 364888 505103 364922
rect 505137 364888 505193 364922
rect 505227 364888 505283 364922
rect 505317 364888 505373 364922
rect 505407 364888 505463 364922
rect 505497 364888 505553 364922
rect 505587 364888 505643 364922
rect 505677 364888 505809 364922
rect 504847 364869 505809 364888
rect 504847 364810 504919 364869
rect 504847 364776 504866 364810
rect 504900 364776 504919 364810
rect 505737 364844 505809 364869
rect 505737 364810 505756 364844
rect 505790 364810 505809 364844
rect 504847 364720 504919 364776
rect 504847 364686 504866 364720
rect 504900 364686 504919 364720
rect 504847 364630 504919 364686
rect 504847 364596 504866 364630
rect 504900 364596 504919 364630
rect 504847 364540 504919 364596
rect 504847 364506 504866 364540
rect 504900 364506 504919 364540
rect 504847 364450 504919 364506
rect 504847 364416 504866 364450
rect 504900 364416 504919 364450
rect 504847 364360 504919 364416
rect 504847 364326 504866 364360
rect 504900 364326 504919 364360
rect 504847 364270 504919 364326
rect 504847 364236 504866 364270
rect 504900 364236 504919 364270
rect 504847 364180 504919 364236
rect 504847 364146 504866 364180
rect 504900 364146 504919 364180
rect 504847 364090 504919 364146
rect 505737 364754 505809 364810
rect 505737 364720 505756 364754
rect 505790 364720 505809 364754
rect 505737 364664 505809 364720
rect 505737 364630 505756 364664
rect 505790 364630 505809 364664
rect 505737 364574 505809 364630
rect 505737 364540 505756 364574
rect 505790 364540 505809 364574
rect 505737 364484 505809 364540
rect 505737 364450 505756 364484
rect 505790 364450 505809 364484
rect 505737 364394 505809 364450
rect 505737 364360 505756 364394
rect 505790 364360 505809 364394
rect 505737 364304 505809 364360
rect 505737 364270 505756 364304
rect 505790 364270 505809 364304
rect 505737 364214 505809 364270
rect 505737 364180 505756 364214
rect 505790 364180 505809 364214
rect 505737 364124 505809 364180
rect 504847 364056 504866 364090
rect 504900 364056 504919 364090
rect 504847 364051 504919 364056
rect 505737 364090 505756 364124
rect 505790 364090 505809 364124
rect 505737 364051 505809 364090
rect 504847 364032 505809 364051
rect 504847 363998 504942 364032
rect 504976 363998 505032 364032
rect 505066 363998 505122 364032
rect 505156 363998 505212 364032
rect 505246 363998 505302 364032
rect 505336 363998 505392 364032
rect 505426 363998 505482 364032
rect 505516 363998 505572 364032
rect 505606 363998 505662 364032
rect 505696 363998 505809 364032
rect 504847 363979 505809 363998
rect 504847 363582 505809 363601
rect 504847 363548 504923 363582
rect 504957 363548 505013 363582
rect 505047 363548 505103 363582
rect 505137 363548 505193 363582
rect 505227 363548 505283 363582
rect 505317 363548 505373 363582
rect 505407 363548 505463 363582
rect 505497 363548 505553 363582
rect 505587 363548 505643 363582
rect 505677 363548 505809 363582
rect 504847 363529 505809 363548
rect 504847 363470 504919 363529
rect 504847 363436 504866 363470
rect 504900 363436 504919 363470
rect 505737 363504 505809 363529
rect 505737 363470 505756 363504
rect 505790 363470 505809 363504
rect 504847 363380 504919 363436
rect 504847 363346 504866 363380
rect 504900 363346 504919 363380
rect 504847 363290 504919 363346
rect 504847 363256 504866 363290
rect 504900 363256 504919 363290
rect 504847 363200 504919 363256
rect 504847 363166 504866 363200
rect 504900 363166 504919 363200
rect 504847 363110 504919 363166
rect 504847 363076 504866 363110
rect 504900 363076 504919 363110
rect 504847 363020 504919 363076
rect 504847 362986 504866 363020
rect 504900 362986 504919 363020
rect 504847 362930 504919 362986
rect 504847 362896 504866 362930
rect 504900 362896 504919 362930
rect 504847 362840 504919 362896
rect 504847 362806 504866 362840
rect 504900 362806 504919 362840
rect 504847 362750 504919 362806
rect 505737 363414 505809 363470
rect 505737 363380 505756 363414
rect 505790 363380 505809 363414
rect 505737 363324 505809 363380
rect 505737 363290 505756 363324
rect 505790 363290 505809 363324
rect 505737 363234 505809 363290
rect 505737 363200 505756 363234
rect 505790 363200 505809 363234
rect 505737 363144 505809 363200
rect 505737 363110 505756 363144
rect 505790 363110 505809 363144
rect 505737 363054 505809 363110
rect 505737 363020 505756 363054
rect 505790 363020 505809 363054
rect 505737 362964 505809 363020
rect 505737 362930 505756 362964
rect 505790 362930 505809 362964
rect 505737 362874 505809 362930
rect 505737 362840 505756 362874
rect 505790 362840 505809 362874
rect 505737 362784 505809 362840
rect 504847 362716 504866 362750
rect 504900 362716 504919 362750
rect 504847 362711 504919 362716
rect 505737 362750 505756 362784
rect 505790 362750 505809 362784
rect 505737 362711 505809 362750
rect 504847 362692 505809 362711
rect 504847 362658 504942 362692
rect 504976 362658 505032 362692
rect 505066 362658 505122 362692
rect 505156 362658 505212 362692
rect 505246 362658 505302 362692
rect 505336 362658 505392 362692
rect 505426 362658 505482 362692
rect 505516 362658 505572 362692
rect 505606 362658 505662 362692
rect 505696 362658 505809 362692
rect 504847 362639 505809 362658
rect 508607 372962 509569 372981
rect 508607 372928 508683 372962
rect 508717 372928 508773 372962
rect 508807 372928 508863 372962
rect 508897 372928 508953 372962
rect 508987 372928 509043 372962
rect 509077 372928 509133 372962
rect 509167 372928 509223 372962
rect 509257 372928 509313 372962
rect 509347 372928 509403 372962
rect 509437 372928 509569 372962
rect 508607 372909 509569 372928
rect 508607 372850 508679 372909
rect 508607 372816 508626 372850
rect 508660 372816 508679 372850
rect 509497 372884 509569 372909
rect 509497 372850 509516 372884
rect 509550 372850 509569 372884
rect 508607 372760 508679 372816
rect 508607 372726 508626 372760
rect 508660 372726 508679 372760
rect 508607 372670 508679 372726
rect 508607 372636 508626 372670
rect 508660 372636 508679 372670
rect 508607 372580 508679 372636
rect 508607 372546 508626 372580
rect 508660 372546 508679 372580
rect 508607 372490 508679 372546
rect 508607 372456 508626 372490
rect 508660 372456 508679 372490
rect 508607 372400 508679 372456
rect 508607 372366 508626 372400
rect 508660 372366 508679 372400
rect 508607 372310 508679 372366
rect 508607 372276 508626 372310
rect 508660 372276 508679 372310
rect 508607 372220 508679 372276
rect 508607 372186 508626 372220
rect 508660 372186 508679 372220
rect 508607 372130 508679 372186
rect 509497 372794 509569 372850
rect 509497 372760 509516 372794
rect 509550 372760 509569 372794
rect 509497 372704 509569 372760
rect 509497 372670 509516 372704
rect 509550 372670 509569 372704
rect 509497 372614 509569 372670
rect 509497 372580 509516 372614
rect 509550 372580 509569 372614
rect 509497 372524 509569 372580
rect 509497 372490 509516 372524
rect 509550 372490 509569 372524
rect 509497 372434 509569 372490
rect 509497 372400 509516 372434
rect 509550 372400 509569 372434
rect 509497 372344 509569 372400
rect 509497 372310 509516 372344
rect 509550 372310 509569 372344
rect 509497 372254 509569 372310
rect 509497 372220 509516 372254
rect 509550 372220 509569 372254
rect 509497 372164 509569 372220
rect 508607 372096 508626 372130
rect 508660 372096 508679 372130
rect 508607 372091 508679 372096
rect 509497 372130 509516 372164
rect 509550 372130 509569 372164
rect 509497 372091 509569 372130
rect 508607 372072 509569 372091
rect 508607 372038 508702 372072
rect 508736 372038 508792 372072
rect 508826 372038 508882 372072
rect 508916 372038 508972 372072
rect 509006 372038 509062 372072
rect 509096 372038 509152 372072
rect 509186 372038 509242 372072
rect 509276 372038 509332 372072
rect 509366 372038 509422 372072
rect 509456 372038 509569 372072
rect 508607 372019 509569 372038
rect 508607 371622 509569 371641
rect 508607 371588 508683 371622
rect 508717 371588 508773 371622
rect 508807 371588 508863 371622
rect 508897 371588 508953 371622
rect 508987 371588 509043 371622
rect 509077 371588 509133 371622
rect 509167 371588 509223 371622
rect 509257 371588 509313 371622
rect 509347 371588 509403 371622
rect 509437 371588 509569 371622
rect 508607 371569 509569 371588
rect 508607 371510 508679 371569
rect 508607 371476 508626 371510
rect 508660 371476 508679 371510
rect 509497 371544 509569 371569
rect 509497 371510 509516 371544
rect 509550 371510 509569 371544
rect 508607 371420 508679 371476
rect 508607 371386 508626 371420
rect 508660 371386 508679 371420
rect 508607 371330 508679 371386
rect 508607 371296 508626 371330
rect 508660 371296 508679 371330
rect 508607 371240 508679 371296
rect 508607 371206 508626 371240
rect 508660 371206 508679 371240
rect 508607 371150 508679 371206
rect 508607 371116 508626 371150
rect 508660 371116 508679 371150
rect 508607 371060 508679 371116
rect 508607 371026 508626 371060
rect 508660 371026 508679 371060
rect 508607 370970 508679 371026
rect 508607 370936 508626 370970
rect 508660 370936 508679 370970
rect 508607 370880 508679 370936
rect 508607 370846 508626 370880
rect 508660 370846 508679 370880
rect 508607 370790 508679 370846
rect 509497 371454 509569 371510
rect 509497 371420 509516 371454
rect 509550 371420 509569 371454
rect 509497 371364 509569 371420
rect 509497 371330 509516 371364
rect 509550 371330 509569 371364
rect 509497 371274 509569 371330
rect 509497 371240 509516 371274
rect 509550 371240 509569 371274
rect 509497 371184 509569 371240
rect 509497 371150 509516 371184
rect 509550 371150 509569 371184
rect 509497 371094 509569 371150
rect 509497 371060 509516 371094
rect 509550 371060 509569 371094
rect 509497 371004 509569 371060
rect 509497 370970 509516 371004
rect 509550 370970 509569 371004
rect 509497 370914 509569 370970
rect 509497 370880 509516 370914
rect 509550 370880 509569 370914
rect 509497 370824 509569 370880
rect 508607 370756 508626 370790
rect 508660 370756 508679 370790
rect 508607 370751 508679 370756
rect 509497 370790 509516 370824
rect 509550 370790 509569 370824
rect 509497 370751 509569 370790
rect 508607 370732 509569 370751
rect 508607 370698 508702 370732
rect 508736 370698 508792 370732
rect 508826 370698 508882 370732
rect 508916 370698 508972 370732
rect 509006 370698 509062 370732
rect 509096 370698 509152 370732
rect 509186 370698 509242 370732
rect 509276 370698 509332 370732
rect 509366 370698 509422 370732
rect 509456 370698 509569 370732
rect 508607 370679 509569 370698
rect 508607 370282 509569 370301
rect 508607 370248 508683 370282
rect 508717 370248 508773 370282
rect 508807 370248 508863 370282
rect 508897 370248 508953 370282
rect 508987 370248 509043 370282
rect 509077 370248 509133 370282
rect 509167 370248 509223 370282
rect 509257 370248 509313 370282
rect 509347 370248 509403 370282
rect 509437 370248 509569 370282
rect 508607 370229 509569 370248
rect 508607 370170 508679 370229
rect 508607 370136 508626 370170
rect 508660 370136 508679 370170
rect 509497 370204 509569 370229
rect 509497 370170 509516 370204
rect 509550 370170 509569 370204
rect 508607 370080 508679 370136
rect 508607 370046 508626 370080
rect 508660 370046 508679 370080
rect 508607 369990 508679 370046
rect 508607 369956 508626 369990
rect 508660 369956 508679 369990
rect 508607 369900 508679 369956
rect 508607 369866 508626 369900
rect 508660 369866 508679 369900
rect 508607 369810 508679 369866
rect 508607 369776 508626 369810
rect 508660 369776 508679 369810
rect 508607 369720 508679 369776
rect 508607 369686 508626 369720
rect 508660 369686 508679 369720
rect 508607 369630 508679 369686
rect 508607 369596 508626 369630
rect 508660 369596 508679 369630
rect 508607 369540 508679 369596
rect 508607 369506 508626 369540
rect 508660 369506 508679 369540
rect 508607 369450 508679 369506
rect 509497 370114 509569 370170
rect 509497 370080 509516 370114
rect 509550 370080 509569 370114
rect 509497 370024 509569 370080
rect 509497 369990 509516 370024
rect 509550 369990 509569 370024
rect 509497 369934 509569 369990
rect 509497 369900 509516 369934
rect 509550 369900 509569 369934
rect 509497 369844 509569 369900
rect 509497 369810 509516 369844
rect 509550 369810 509569 369844
rect 509497 369754 509569 369810
rect 509497 369720 509516 369754
rect 509550 369720 509569 369754
rect 509497 369664 509569 369720
rect 509497 369630 509516 369664
rect 509550 369630 509569 369664
rect 509497 369574 509569 369630
rect 509497 369540 509516 369574
rect 509550 369540 509569 369574
rect 509497 369484 509569 369540
rect 508607 369416 508626 369450
rect 508660 369416 508679 369450
rect 508607 369411 508679 369416
rect 509497 369450 509516 369484
rect 509550 369450 509569 369484
rect 509497 369411 509569 369450
rect 508607 369392 509569 369411
rect 508607 369358 508702 369392
rect 508736 369358 508792 369392
rect 508826 369358 508882 369392
rect 508916 369358 508972 369392
rect 509006 369358 509062 369392
rect 509096 369358 509152 369392
rect 509186 369358 509242 369392
rect 509276 369358 509332 369392
rect 509366 369358 509422 369392
rect 509456 369358 509569 369392
rect 508607 369339 509569 369358
rect 508607 368942 509569 368961
rect 508607 368908 508683 368942
rect 508717 368908 508773 368942
rect 508807 368908 508863 368942
rect 508897 368908 508953 368942
rect 508987 368908 509043 368942
rect 509077 368908 509133 368942
rect 509167 368908 509223 368942
rect 509257 368908 509313 368942
rect 509347 368908 509403 368942
rect 509437 368908 509569 368942
rect 508607 368889 509569 368908
rect 508607 368830 508679 368889
rect 508607 368796 508626 368830
rect 508660 368796 508679 368830
rect 509497 368864 509569 368889
rect 509497 368830 509516 368864
rect 509550 368830 509569 368864
rect 508607 368740 508679 368796
rect 508607 368706 508626 368740
rect 508660 368706 508679 368740
rect 508607 368650 508679 368706
rect 508607 368616 508626 368650
rect 508660 368616 508679 368650
rect 508607 368560 508679 368616
rect 508607 368526 508626 368560
rect 508660 368526 508679 368560
rect 508607 368470 508679 368526
rect 508607 368436 508626 368470
rect 508660 368436 508679 368470
rect 508607 368380 508679 368436
rect 508607 368346 508626 368380
rect 508660 368346 508679 368380
rect 508607 368290 508679 368346
rect 508607 368256 508626 368290
rect 508660 368256 508679 368290
rect 508607 368200 508679 368256
rect 508607 368166 508626 368200
rect 508660 368166 508679 368200
rect 508607 368110 508679 368166
rect 509497 368774 509569 368830
rect 509497 368740 509516 368774
rect 509550 368740 509569 368774
rect 509497 368684 509569 368740
rect 509497 368650 509516 368684
rect 509550 368650 509569 368684
rect 509497 368594 509569 368650
rect 509497 368560 509516 368594
rect 509550 368560 509569 368594
rect 509497 368504 509569 368560
rect 509497 368470 509516 368504
rect 509550 368470 509569 368504
rect 509497 368414 509569 368470
rect 509497 368380 509516 368414
rect 509550 368380 509569 368414
rect 509497 368324 509569 368380
rect 509497 368290 509516 368324
rect 509550 368290 509569 368324
rect 509497 368234 509569 368290
rect 509497 368200 509516 368234
rect 509550 368200 509569 368234
rect 509497 368144 509569 368200
rect 508607 368076 508626 368110
rect 508660 368076 508679 368110
rect 508607 368071 508679 368076
rect 509497 368110 509516 368144
rect 509550 368110 509569 368144
rect 509497 368071 509569 368110
rect 508607 368052 509569 368071
rect 508607 368018 508702 368052
rect 508736 368018 508792 368052
rect 508826 368018 508882 368052
rect 508916 368018 508972 368052
rect 509006 368018 509062 368052
rect 509096 368018 509152 368052
rect 509186 368018 509242 368052
rect 509276 368018 509332 368052
rect 509366 368018 509422 368052
rect 509456 368018 509569 368052
rect 508607 367999 509569 368018
rect 508607 367602 509569 367621
rect 508607 367568 508683 367602
rect 508717 367568 508773 367602
rect 508807 367568 508863 367602
rect 508897 367568 508953 367602
rect 508987 367568 509043 367602
rect 509077 367568 509133 367602
rect 509167 367568 509223 367602
rect 509257 367568 509313 367602
rect 509347 367568 509403 367602
rect 509437 367568 509569 367602
rect 508607 367549 509569 367568
rect 508607 367490 508679 367549
rect 508607 367456 508626 367490
rect 508660 367456 508679 367490
rect 509497 367524 509569 367549
rect 509497 367490 509516 367524
rect 509550 367490 509569 367524
rect 508607 367400 508679 367456
rect 508607 367366 508626 367400
rect 508660 367366 508679 367400
rect 508607 367310 508679 367366
rect 508607 367276 508626 367310
rect 508660 367276 508679 367310
rect 508607 367220 508679 367276
rect 508607 367186 508626 367220
rect 508660 367186 508679 367220
rect 508607 367130 508679 367186
rect 508607 367096 508626 367130
rect 508660 367096 508679 367130
rect 508607 367040 508679 367096
rect 508607 367006 508626 367040
rect 508660 367006 508679 367040
rect 508607 366950 508679 367006
rect 508607 366916 508626 366950
rect 508660 366916 508679 366950
rect 508607 366860 508679 366916
rect 508607 366826 508626 366860
rect 508660 366826 508679 366860
rect 508607 366770 508679 366826
rect 509497 367434 509569 367490
rect 509497 367400 509516 367434
rect 509550 367400 509569 367434
rect 509497 367344 509569 367400
rect 509497 367310 509516 367344
rect 509550 367310 509569 367344
rect 509497 367254 509569 367310
rect 509497 367220 509516 367254
rect 509550 367220 509569 367254
rect 509497 367164 509569 367220
rect 509497 367130 509516 367164
rect 509550 367130 509569 367164
rect 509497 367074 509569 367130
rect 509497 367040 509516 367074
rect 509550 367040 509569 367074
rect 509497 366984 509569 367040
rect 509497 366950 509516 366984
rect 509550 366950 509569 366984
rect 509497 366894 509569 366950
rect 509497 366860 509516 366894
rect 509550 366860 509569 366894
rect 509497 366804 509569 366860
rect 508607 366736 508626 366770
rect 508660 366736 508679 366770
rect 508607 366731 508679 366736
rect 509497 366770 509516 366804
rect 509550 366770 509569 366804
rect 509497 366731 509569 366770
rect 508607 366712 509569 366731
rect 508607 366678 508702 366712
rect 508736 366678 508792 366712
rect 508826 366678 508882 366712
rect 508916 366678 508972 366712
rect 509006 366678 509062 366712
rect 509096 366678 509152 366712
rect 509186 366678 509242 366712
rect 509276 366678 509332 366712
rect 509366 366678 509422 366712
rect 509456 366678 509569 366712
rect 508607 366659 509569 366678
rect 508607 366262 509569 366281
rect 508607 366228 508683 366262
rect 508717 366228 508773 366262
rect 508807 366228 508863 366262
rect 508897 366228 508953 366262
rect 508987 366228 509043 366262
rect 509077 366228 509133 366262
rect 509167 366228 509223 366262
rect 509257 366228 509313 366262
rect 509347 366228 509403 366262
rect 509437 366228 509569 366262
rect 508607 366209 509569 366228
rect 508607 366150 508679 366209
rect 508607 366116 508626 366150
rect 508660 366116 508679 366150
rect 509497 366184 509569 366209
rect 509497 366150 509516 366184
rect 509550 366150 509569 366184
rect 508607 366060 508679 366116
rect 508607 366026 508626 366060
rect 508660 366026 508679 366060
rect 508607 365970 508679 366026
rect 508607 365936 508626 365970
rect 508660 365936 508679 365970
rect 508607 365880 508679 365936
rect 508607 365846 508626 365880
rect 508660 365846 508679 365880
rect 508607 365790 508679 365846
rect 508607 365756 508626 365790
rect 508660 365756 508679 365790
rect 508607 365700 508679 365756
rect 508607 365666 508626 365700
rect 508660 365666 508679 365700
rect 508607 365610 508679 365666
rect 508607 365576 508626 365610
rect 508660 365576 508679 365610
rect 508607 365520 508679 365576
rect 508607 365486 508626 365520
rect 508660 365486 508679 365520
rect 508607 365430 508679 365486
rect 509497 366094 509569 366150
rect 509497 366060 509516 366094
rect 509550 366060 509569 366094
rect 509497 366004 509569 366060
rect 509497 365970 509516 366004
rect 509550 365970 509569 366004
rect 509497 365914 509569 365970
rect 509497 365880 509516 365914
rect 509550 365880 509569 365914
rect 509497 365824 509569 365880
rect 509497 365790 509516 365824
rect 509550 365790 509569 365824
rect 509497 365734 509569 365790
rect 509497 365700 509516 365734
rect 509550 365700 509569 365734
rect 509497 365644 509569 365700
rect 509497 365610 509516 365644
rect 509550 365610 509569 365644
rect 509497 365554 509569 365610
rect 509497 365520 509516 365554
rect 509550 365520 509569 365554
rect 509497 365464 509569 365520
rect 508607 365396 508626 365430
rect 508660 365396 508679 365430
rect 508607 365391 508679 365396
rect 509497 365430 509516 365464
rect 509550 365430 509569 365464
rect 509497 365391 509569 365430
rect 508607 365372 509569 365391
rect 508607 365338 508702 365372
rect 508736 365338 508792 365372
rect 508826 365338 508882 365372
rect 508916 365338 508972 365372
rect 509006 365338 509062 365372
rect 509096 365338 509152 365372
rect 509186 365338 509242 365372
rect 509276 365338 509332 365372
rect 509366 365338 509422 365372
rect 509456 365338 509569 365372
rect 508607 365319 509569 365338
rect 508607 364922 509569 364941
rect 508607 364888 508683 364922
rect 508717 364888 508773 364922
rect 508807 364888 508863 364922
rect 508897 364888 508953 364922
rect 508987 364888 509043 364922
rect 509077 364888 509133 364922
rect 509167 364888 509223 364922
rect 509257 364888 509313 364922
rect 509347 364888 509403 364922
rect 509437 364888 509569 364922
rect 508607 364869 509569 364888
rect 508607 364810 508679 364869
rect 508607 364776 508626 364810
rect 508660 364776 508679 364810
rect 509497 364844 509569 364869
rect 509497 364810 509516 364844
rect 509550 364810 509569 364844
rect 508607 364720 508679 364776
rect 508607 364686 508626 364720
rect 508660 364686 508679 364720
rect 508607 364630 508679 364686
rect 508607 364596 508626 364630
rect 508660 364596 508679 364630
rect 508607 364540 508679 364596
rect 508607 364506 508626 364540
rect 508660 364506 508679 364540
rect 508607 364450 508679 364506
rect 508607 364416 508626 364450
rect 508660 364416 508679 364450
rect 508607 364360 508679 364416
rect 508607 364326 508626 364360
rect 508660 364326 508679 364360
rect 508607 364270 508679 364326
rect 508607 364236 508626 364270
rect 508660 364236 508679 364270
rect 508607 364180 508679 364236
rect 508607 364146 508626 364180
rect 508660 364146 508679 364180
rect 508607 364090 508679 364146
rect 509497 364754 509569 364810
rect 509497 364720 509516 364754
rect 509550 364720 509569 364754
rect 509497 364664 509569 364720
rect 509497 364630 509516 364664
rect 509550 364630 509569 364664
rect 509497 364574 509569 364630
rect 509497 364540 509516 364574
rect 509550 364540 509569 364574
rect 509497 364484 509569 364540
rect 509497 364450 509516 364484
rect 509550 364450 509569 364484
rect 509497 364394 509569 364450
rect 509497 364360 509516 364394
rect 509550 364360 509569 364394
rect 509497 364304 509569 364360
rect 509497 364270 509516 364304
rect 509550 364270 509569 364304
rect 509497 364214 509569 364270
rect 509497 364180 509516 364214
rect 509550 364180 509569 364214
rect 509497 364124 509569 364180
rect 508607 364056 508626 364090
rect 508660 364056 508679 364090
rect 508607 364051 508679 364056
rect 509497 364090 509516 364124
rect 509550 364090 509569 364124
rect 509497 364051 509569 364090
rect 508607 364032 509569 364051
rect 508607 363998 508702 364032
rect 508736 363998 508792 364032
rect 508826 363998 508882 364032
rect 508916 363998 508972 364032
rect 509006 363998 509062 364032
rect 509096 363998 509152 364032
rect 509186 363998 509242 364032
rect 509276 363998 509332 364032
rect 509366 363998 509422 364032
rect 509456 363998 509569 364032
rect 508607 363979 509569 363998
rect 508607 363582 509569 363601
rect 508607 363548 508683 363582
rect 508717 363548 508773 363582
rect 508807 363548 508863 363582
rect 508897 363548 508953 363582
rect 508987 363548 509043 363582
rect 509077 363548 509133 363582
rect 509167 363548 509223 363582
rect 509257 363548 509313 363582
rect 509347 363548 509403 363582
rect 509437 363548 509569 363582
rect 508607 363529 509569 363548
rect 508607 363470 508679 363529
rect 508607 363436 508626 363470
rect 508660 363436 508679 363470
rect 509497 363504 509569 363529
rect 509497 363470 509516 363504
rect 509550 363470 509569 363504
rect 508607 363380 508679 363436
rect 508607 363346 508626 363380
rect 508660 363346 508679 363380
rect 508607 363290 508679 363346
rect 508607 363256 508626 363290
rect 508660 363256 508679 363290
rect 508607 363200 508679 363256
rect 508607 363166 508626 363200
rect 508660 363166 508679 363200
rect 508607 363110 508679 363166
rect 508607 363076 508626 363110
rect 508660 363076 508679 363110
rect 508607 363020 508679 363076
rect 508607 362986 508626 363020
rect 508660 362986 508679 363020
rect 508607 362930 508679 362986
rect 508607 362896 508626 362930
rect 508660 362896 508679 362930
rect 508607 362840 508679 362896
rect 508607 362806 508626 362840
rect 508660 362806 508679 362840
rect 508607 362750 508679 362806
rect 509497 363414 509569 363470
rect 509497 363380 509516 363414
rect 509550 363380 509569 363414
rect 509497 363324 509569 363380
rect 509497 363290 509516 363324
rect 509550 363290 509569 363324
rect 509497 363234 509569 363290
rect 509497 363200 509516 363234
rect 509550 363200 509569 363234
rect 509497 363144 509569 363200
rect 509497 363110 509516 363144
rect 509550 363110 509569 363144
rect 509497 363054 509569 363110
rect 509497 363020 509516 363054
rect 509550 363020 509569 363054
rect 509497 362964 509569 363020
rect 509497 362930 509516 362964
rect 509550 362930 509569 362964
rect 509497 362874 509569 362930
rect 509497 362840 509516 362874
rect 509550 362840 509569 362874
rect 509497 362784 509569 362840
rect 508607 362716 508626 362750
rect 508660 362716 508679 362750
rect 508607 362711 508679 362716
rect 509497 362750 509516 362784
rect 509550 362750 509569 362784
rect 509497 362711 509569 362750
rect 508607 362692 509569 362711
rect 508607 362658 508702 362692
rect 508736 362658 508792 362692
rect 508826 362658 508882 362692
rect 508916 362658 508972 362692
rect 509006 362658 509062 362692
rect 509096 362658 509152 362692
rect 509186 362658 509242 362692
rect 509276 362658 509332 362692
rect 509366 362658 509422 362692
rect 509456 362658 509569 362692
rect 508607 362639 509569 362658
rect 512367 372962 513329 372981
rect 512367 372928 512443 372962
rect 512477 372928 512533 372962
rect 512567 372928 512623 372962
rect 512657 372928 512713 372962
rect 512747 372928 512803 372962
rect 512837 372928 512893 372962
rect 512927 372928 512983 372962
rect 513017 372928 513073 372962
rect 513107 372928 513163 372962
rect 513197 372928 513329 372962
rect 512367 372909 513329 372928
rect 512367 372850 512439 372909
rect 512367 372816 512386 372850
rect 512420 372816 512439 372850
rect 513257 372884 513329 372909
rect 513257 372850 513276 372884
rect 513310 372850 513329 372884
rect 512367 372760 512439 372816
rect 512367 372726 512386 372760
rect 512420 372726 512439 372760
rect 512367 372670 512439 372726
rect 512367 372636 512386 372670
rect 512420 372636 512439 372670
rect 512367 372580 512439 372636
rect 512367 372546 512386 372580
rect 512420 372546 512439 372580
rect 512367 372490 512439 372546
rect 512367 372456 512386 372490
rect 512420 372456 512439 372490
rect 512367 372400 512439 372456
rect 512367 372366 512386 372400
rect 512420 372366 512439 372400
rect 512367 372310 512439 372366
rect 512367 372276 512386 372310
rect 512420 372276 512439 372310
rect 512367 372220 512439 372276
rect 512367 372186 512386 372220
rect 512420 372186 512439 372220
rect 512367 372130 512439 372186
rect 513257 372794 513329 372850
rect 513257 372760 513276 372794
rect 513310 372760 513329 372794
rect 513257 372704 513329 372760
rect 513257 372670 513276 372704
rect 513310 372670 513329 372704
rect 513257 372614 513329 372670
rect 513257 372580 513276 372614
rect 513310 372580 513329 372614
rect 513257 372524 513329 372580
rect 513257 372490 513276 372524
rect 513310 372490 513329 372524
rect 513257 372434 513329 372490
rect 513257 372400 513276 372434
rect 513310 372400 513329 372434
rect 513257 372344 513329 372400
rect 513257 372310 513276 372344
rect 513310 372310 513329 372344
rect 513257 372254 513329 372310
rect 513257 372220 513276 372254
rect 513310 372220 513329 372254
rect 513257 372164 513329 372220
rect 512367 372096 512386 372130
rect 512420 372096 512439 372130
rect 512367 372091 512439 372096
rect 513257 372130 513276 372164
rect 513310 372130 513329 372164
rect 513257 372091 513329 372130
rect 512367 372072 513329 372091
rect 512367 372038 512462 372072
rect 512496 372038 512552 372072
rect 512586 372038 512642 372072
rect 512676 372038 512732 372072
rect 512766 372038 512822 372072
rect 512856 372038 512912 372072
rect 512946 372038 513002 372072
rect 513036 372038 513092 372072
rect 513126 372038 513182 372072
rect 513216 372038 513329 372072
rect 512367 372019 513329 372038
rect 523258 374781 523298 374826
rect 523258 374747 523261 374781
rect 523295 374747 523298 374781
rect 523258 374706 523298 374747
rect 523258 373481 523298 373526
rect 523258 373447 523261 373481
rect 523295 373447 523298 373481
rect 523258 373406 523298 373447
rect 523258 372181 523298 372226
rect 523258 372147 523261 372181
rect 523295 372147 523298 372181
rect 523258 372106 523298 372147
rect 512367 371622 513329 371641
rect 512367 371588 512443 371622
rect 512477 371588 512533 371622
rect 512567 371588 512623 371622
rect 512657 371588 512713 371622
rect 512747 371588 512803 371622
rect 512837 371588 512893 371622
rect 512927 371588 512983 371622
rect 513017 371588 513073 371622
rect 513107 371588 513163 371622
rect 513197 371588 513329 371622
rect 512367 371569 513329 371588
rect 512367 371510 512439 371569
rect 512367 371476 512386 371510
rect 512420 371476 512439 371510
rect 513257 371544 513329 371569
rect 513257 371510 513276 371544
rect 513310 371510 513329 371544
rect 512367 371420 512439 371476
rect 512367 371386 512386 371420
rect 512420 371386 512439 371420
rect 512367 371330 512439 371386
rect 512367 371296 512386 371330
rect 512420 371296 512439 371330
rect 512367 371240 512439 371296
rect 512367 371206 512386 371240
rect 512420 371206 512439 371240
rect 512367 371150 512439 371206
rect 512367 371116 512386 371150
rect 512420 371116 512439 371150
rect 512367 371060 512439 371116
rect 512367 371026 512386 371060
rect 512420 371026 512439 371060
rect 512367 370970 512439 371026
rect 512367 370936 512386 370970
rect 512420 370936 512439 370970
rect 512367 370880 512439 370936
rect 512367 370846 512386 370880
rect 512420 370846 512439 370880
rect 512367 370790 512439 370846
rect 513257 371454 513329 371510
rect 513257 371420 513276 371454
rect 513310 371420 513329 371454
rect 513257 371364 513329 371420
rect 513257 371330 513276 371364
rect 513310 371330 513329 371364
rect 513257 371274 513329 371330
rect 513257 371240 513276 371274
rect 513310 371240 513329 371274
rect 513257 371184 513329 371240
rect 513257 371150 513276 371184
rect 513310 371150 513329 371184
rect 513257 371094 513329 371150
rect 513257 371060 513276 371094
rect 513310 371060 513329 371094
rect 513257 371004 513329 371060
rect 513257 370970 513276 371004
rect 513310 370970 513329 371004
rect 513257 370914 513329 370970
rect 513257 370880 513276 370914
rect 513310 370880 513329 370914
rect 513257 370824 513329 370880
rect 512367 370756 512386 370790
rect 512420 370756 512439 370790
rect 512367 370751 512439 370756
rect 513257 370790 513276 370824
rect 513310 370790 513329 370824
rect 513257 370751 513329 370790
rect 512367 370732 513329 370751
rect 512367 370698 512462 370732
rect 512496 370698 512552 370732
rect 512586 370698 512642 370732
rect 512676 370698 512732 370732
rect 512766 370698 512822 370732
rect 512856 370698 512912 370732
rect 512946 370698 513002 370732
rect 513036 370698 513092 370732
rect 513126 370698 513182 370732
rect 513216 370698 513329 370732
rect 512367 370679 513329 370698
rect 512367 370282 513329 370301
rect 512367 370248 512443 370282
rect 512477 370248 512533 370282
rect 512567 370248 512623 370282
rect 512657 370248 512713 370282
rect 512747 370248 512803 370282
rect 512837 370248 512893 370282
rect 512927 370248 512983 370282
rect 513017 370248 513073 370282
rect 513107 370248 513163 370282
rect 513197 370248 513329 370282
rect 512367 370229 513329 370248
rect 512367 370170 512439 370229
rect 512367 370136 512386 370170
rect 512420 370136 512439 370170
rect 513257 370204 513329 370229
rect 513257 370170 513276 370204
rect 513310 370170 513329 370204
rect 512367 370080 512439 370136
rect 512367 370046 512386 370080
rect 512420 370046 512439 370080
rect 512367 369990 512439 370046
rect 512367 369956 512386 369990
rect 512420 369956 512439 369990
rect 512367 369900 512439 369956
rect 512367 369866 512386 369900
rect 512420 369866 512439 369900
rect 512367 369810 512439 369866
rect 512367 369776 512386 369810
rect 512420 369776 512439 369810
rect 512367 369720 512439 369776
rect 512367 369686 512386 369720
rect 512420 369686 512439 369720
rect 512367 369630 512439 369686
rect 512367 369596 512386 369630
rect 512420 369596 512439 369630
rect 512367 369540 512439 369596
rect 512367 369506 512386 369540
rect 512420 369506 512439 369540
rect 512367 369450 512439 369506
rect 513257 370114 513329 370170
rect 513257 370080 513276 370114
rect 513310 370080 513329 370114
rect 513257 370024 513329 370080
rect 513257 369990 513276 370024
rect 513310 369990 513329 370024
rect 513257 369934 513329 369990
rect 513257 369900 513276 369934
rect 513310 369900 513329 369934
rect 513257 369844 513329 369900
rect 513257 369810 513276 369844
rect 513310 369810 513329 369844
rect 513257 369754 513329 369810
rect 513257 369720 513276 369754
rect 513310 369720 513329 369754
rect 513257 369664 513329 369720
rect 513257 369630 513276 369664
rect 513310 369630 513329 369664
rect 513257 369574 513329 369630
rect 513257 369540 513276 369574
rect 513310 369540 513329 369574
rect 513257 369484 513329 369540
rect 512367 369416 512386 369450
rect 512420 369416 512439 369450
rect 512367 369411 512439 369416
rect 513257 369450 513276 369484
rect 513310 369450 513329 369484
rect 513257 369411 513329 369450
rect 512367 369392 513329 369411
rect 512367 369358 512462 369392
rect 512496 369358 512552 369392
rect 512586 369358 512642 369392
rect 512676 369358 512732 369392
rect 512766 369358 512822 369392
rect 512856 369358 512912 369392
rect 512946 369358 513002 369392
rect 513036 369358 513092 369392
rect 513126 369358 513182 369392
rect 513216 369358 513329 369392
rect 512367 369339 513329 369358
rect 523258 370881 523298 370926
rect 523258 370847 523261 370881
rect 523295 370847 523298 370881
rect 523258 370806 523298 370847
rect 523258 369581 523298 369626
rect 523258 369547 523261 369581
rect 523295 369547 523298 369581
rect 523258 369506 523298 369547
rect 512367 368942 513329 368961
rect 512367 368908 512443 368942
rect 512477 368908 512533 368942
rect 512567 368908 512623 368942
rect 512657 368908 512713 368942
rect 512747 368908 512803 368942
rect 512837 368908 512893 368942
rect 512927 368908 512983 368942
rect 513017 368908 513073 368942
rect 513107 368908 513163 368942
rect 513197 368908 513329 368942
rect 512367 368889 513329 368908
rect 512367 368830 512439 368889
rect 512367 368796 512386 368830
rect 512420 368796 512439 368830
rect 513257 368864 513329 368889
rect 513257 368830 513276 368864
rect 513310 368830 513329 368864
rect 512367 368740 512439 368796
rect 512367 368706 512386 368740
rect 512420 368706 512439 368740
rect 512367 368650 512439 368706
rect 512367 368616 512386 368650
rect 512420 368616 512439 368650
rect 512367 368560 512439 368616
rect 512367 368526 512386 368560
rect 512420 368526 512439 368560
rect 512367 368470 512439 368526
rect 512367 368436 512386 368470
rect 512420 368436 512439 368470
rect 512367 368380 512439 368436
rect 512367 368346 512386 368380
rect 512420 368346 512439 368380
rect 512367 368290 512439 368346
rect 512367 368256 512386 368290
rect 512420 368256 512439 368290
rect 512367 368200 512439 368256
rect 512367 368166 512386 368200
rect 512420 368166 512439 368200
rect 512367 368110 512439 368166
rect 513257 368774 513329 368830
rect 513257 368740 513276 368774
rect 513310 368740 513329 368774
rect 513257 368684 513329 368740
rect 513257 368650 513276 368684
rect 513310 368650 513329 368684
rect 513257 368594 513329 368650
rect 513257 368560 513276 368594
rect 513310 368560 513329 368594
rect 513257 368504 513329 368560
rect 513257 368470 513276 368504
rect 513310 368470 513329 368504
rect 513257 368414 513329 368470
rect 513257 368380 513276 368414
rect 513310 368380 513329 368414
rect 513257 368324 513329 368380
rect 513257 368290 513276 368324
rect 513310 368290 513329 368324
rect 513257 368234 513329 368290
rect 513257 368200 513276 368234
rect 513310 368200 513329 368234
rect 513257 368144 513329 368200
rect 512367 368076 512386 368110
rect 512420 368076 512439 368110
rect 512367 368071 512439 368076
rect 513257 368110 513276 368144
rect 513310 368110 513329 368144
rect 513257 368071 513329 368110
rect 512367 368052 513329 368071
rect 512367 368018 512462 368052
rect 512496 368018 512552 368052
rect 512586 368018 512642 368052
rect 512676 368018 512732 368052
rect 512766 368018 512822 368052
rect 512856 368018 512912 368052
rect 512946 368018 513002 368052
rect 513036 368018 513092 368052
rect 513126 368018 513182 368052
rect 513216 368018 513329 368052
rect 512367 367999 513329 368018
rect 512367 367602 513329 367621
rect 512367 367568 512443 367602
rect 512477 367568 512533 367602
rect 512567 367568 512623 367602
rect 512657 367568 512713 367602
rect 512747 367568 512803 367602
rect 512837 367568 512893 367602
rect 512927 367568 512983 367602
rect 513017 367568 513073 367602
rect 513107 367568 513163 367602
rect 513197 367568 513329 367602
rect 512367 367549 513329 367568
rect 512367 367490 512439 367549
rect 512367 367456 512386 367490
rect 512420 367456 512439 367490
rect 513257 367524 513329 367549
rect 513257 367490 513276 367524
rect 513310 367490 513329 367524
rect 512367 367400 512439 367456
rect 512367 367366 512386 367400
rect 512420 367366 512439 367400
rect 512367 367310 512439 367366
rect 512367 367276 512386 367310
rect 512420 367276 512439 367310
rect 512367 367220 512439 367276
rect 512367 367186 512386 367220
rect 512420 367186 512439 367220
rect 512367 367130 512439 367186
rect 512367 367096 512386 367130
rect 512420 367096 512439 367130
rect 512367 367040 512439 367096
rect 512367 367006 512386 367040
rect 512420 367006 512439 367040
rect 512367 366950 512439 367006
rect 512367 366916 512386 366950
rect 512420 366916 512439 366950
rect 512367 366860 512439 366916
rect 512367 366826 512386 366860
rect 512420 366826 512439 366860
rect 512367 366770 512439 366826
rect 513257 367434 513329 367490
rect 513257 367400 513276 367434
rect 513310 367400 513329 367434
rect 513257 367344 513329 367400
rect 513257 367310 513276 367344
rect 513310 367310 513329 367344
rect 513257 367254 513329 367310
rect 513257 367220 513276 367254
rect 513310 367220 513329 367254
rect 513257 367164 513329 367220
rect 513257 367130 513276 367164
rect 513310 367130 513329 367164
rect 513257 367074 513329 367130
rect 513257 367040 513276 367074
rect 513310 367040 513329 367074
rect 513257 366984 513329 367040
rect 513257 366950 513276 366984
rect 513310 366950 513329 366984
rect 513257 366894 513329 366950
rect 513257 366860 513276 366894
rect 513310 366860 513329 366894
rect 513257 366804 513329 366860
rect 512367 366736 512386 366770
rect 512420 366736 512439 366770
rect 512367 366731 512439 366736
rect 513257 366770 513276 366804
rect 513310 366770 513329 366804
rect 513257 366731 513329 366770
rect 512367 366712 513329 366731
rect 512367 366678 512462 366712
rect 512496 366678 512552 366712
rect 512586 366678 512642 366712
rect 512676 366678 512732 366712
rect 512766 366678 512822 366712
rect 512856 366678 512912 366712
rect 512946 366678 513002 366712
rect 513036 366678 513092 366712
rect 513126 366678 513182 366712
rect 513216 366678 513329 366712
rect 512367 366659 513329 366678
rect 523258 368281 523298 368326
rect 523258 368247 523261 368281
rect 523295 368247 523298 368281
rect 523258 368206 523298 368247
rect 523258 366981 523298 367026
rect 523258 366947 523261 366981
rect 523295 366947 523298 366981
rect 523258 366906 523298 366947
rect 512367 366262 513329 366281
rect 512367 366228 512443 366262
rect 512477 366228 512533 366262
rect 512567 366228 512623 366262
rect 512657 366228 512713 366262
rect 512747 366228 512803 366262
rect 512837 366228 512893 366262
rect 512927 366228 512983 366262
rect 513017 366228 513073 366262
rect 513107 366228 513163 366262
rect 513197 366228 513329 366262
rect 512367 366209 513329 366228
rect 512367 366150 512439 366209
rect 512367 366116 512386 366150
rect 512420 366116 512439 366150
rect 513257 366184 513329 366209
rect 513257 366150 513276 366184
rect 513310 366150 513329 366184
rect 512367 366060 512439 366116
rect 512367 366026 512386 366060
rect 512420 366026 512439 366060
rect 512367 365970 512439 366026
rect 512367 365936 512386 365970
rect 512420 365936 512439 365970
rect 512367 365880 512439 365936
rect 512367 365846 512386 365880
rect 512420 365846 512439 365880
rect 512367 365790 512439 365846
rect 512367 365756 512386 365790
rect 512420 365756 512439 365790
rect 512367 365700 512439 365756
rect 512367 365666 512386 365700
rect 512420 365666 512439 365700
rect 512367 365610 512439 365666
rect 512367 365576 512386 365610
rect 512420 365576 512439 365610
rect 512367 365520 512439 365576
rect 512367 365486 512386 365520
rect 512420 365486 512439 365520
rect 512367 365430 512439 365486
rect 513257 366094 513329 366150
rect 513257 366060 513276 366094
rect 513310 366060 513329 366094
rect 513257 366004 513329 366060
rect 513257 365970 513276 366004
rect 513310 365970 513329 366004
rect 513257 365914 513329 365970
rect 513257 365880 513276 365914
rect 513310 365880 513329 365914
rect 513257 365824 513329 365880
rect 513257 365790 513276 365824
rect 513310 365790 513329 365824
rect 513257 365734 513329 365790
rect 513257 365700 513276 365734
rect 513310 365700 513329 365734
rect 513257 365644 513329 365700
rect 513257 365610 513276 365644
rect 513310 365610 513329 365644
rect 513257 365554 513329 365610
rect 513257 365520 513276 365554
rect 513310 365520 513329 365554
rect 513257 365464 513329 365520
rect 512367 365396 512386 365430
rect 512420 365396 512439 365430
rect 512367 365391 512439 365396
rect 513257 365430 513276 365464
rect 513310 365430 513329 365464
rect 513257 365391 513329 365430
rect 512367 365372 513329 365391
rect 512367 365338 512462 365372
rect 512496 365338 512552 365372
rect 512586 365338 512642 365372
rect 512676 365338 512732 365372
rect 512766 365338 512822 365372
rect 512856 365338 512912 365372
rect 512946 365338 513002 365372
rect 513036 365338 513092 365372
rect 513126 365338 513182 365372
rect 513216 365338 513329 365372
rect 512367 365319 513329 365338
rect 512367 364922 513329 364941
rect 512367 364888 512443 364922
rect 512477 364888 512533 364922
rect 512567 364888 512623 364922
rect 512657 364888 512713 364922
rect 512747 364888 512803 364922
rect 512837 364888 512893 364922
rect 512927 364888 512983 364922
rect 513017 364888 513073 364922
rect 513107 364888 513163 364922
rect 513197 364888 513329 364922
rect 512367 364869 513329 364888
rect 512367 364810 512439 364869
rect 512367 364776 512386 364810
rect 512420 364776 512439 364810
rect 513257 364844 513329 364869
rect 513257 364810 513276 364844
rect 513310 364810 513329 364844
rect 512367 364720 512439 364776
rect 512367 364686 512386 364720
rect 512420 364686 512439 364720
rect 512367 364630 512439 364686
rect 512367 364596 512386 364630
rect 512420 364596 512439 364630
rect 512367 364540 512439 364596
rect 512367 364506 512386 364540
rect 512420 364506 512439 364540
rect 512367 364450 512439 364506
rect 512367 364416 512386 364450
rect 512420 364416 512439 364450
rect 512367 364360 512439 364416
rect 512367 364326 512386 364360
rect 512420 364326 512439 364360
rect 512367 364270 512439 364326
rect 512367 364236 512386 364270
rect 512420 364236 512439 364270
rect 512367 364180 512439 364236
rect 512367 364146 512386 364180
rect 512420 364146 512439 364180
rect 512367 364090 512439 364146
rect 513257 364754 513329 364810
rect 513257 364720 513276 364754
rect 513310 364720 513329 364754
rect 513257 364664 513329 364720
rect 513257 364630 513276 364664
rect 513310 364630 513329 364664
rect 513257 364574 513329 364630
rect 513257 364540 513276 364574
rect 513310 364540 513329 364574
rect 513257 364484 513329 364540
rect 513257 364450 513276 364484
rect 513310 364450 513329 364484
rect 513257 364394 513329 364450
rect 513257 364360 513276 364394
rect 513310 364360 513329 364394
rect 513257 364304 513329 364360
rect 513257 364270 513276 364304
rect 513310 364270 513329 364304
rect 513257 364214 513329 364270
rect 513257 364180 513276 364214
rect 513310 364180 513329 364214
rect 513257 364124 513329 364180
rect 512367 364056 512386 364090
rect 512420 364056 512439 364090
rect 512367 364051 512439 364056
rect 513257 364090 513276 364124
rect 513310 364090 513329 364124
rect 513257 364051 513329 364090
rect 512367 364032 513329 364051
rect 512367 363998 512462 364032
rect 512496 363998 512552 364032
rect 512586 363998 512642 364032
rect 512676 363998 512732 364032
rect 512766 363998 512822 364032
rect 512856 363998 512912 364032
rect 512946 363998 513002 364032
rect 513036 363998 513092 364032
rect 513126 363998 513182 364032
rect 513216 363998 513329 364032
rect 512367 363979 513329 363998
rect 523258 365681 523298 365726
rect 523258 365647 523261 365681
rect 523295 365647 523298 365681
rect 523258 365606 523298 365647
rect 523258 364381 523298 364426
rect 523258 364347 523261 364381
rect 523295 364347 523298 364381
rect 523258 364306 523298 364347
rect 512367 363582 513329 363601
rect 512367 363548 512443 363582
rect 512477 363548 512533 363582
rect 512567 363548 512623 363582
rect 512657 363548 512713 363582
rect 512747 363548 512803 363582
rect 512837 363548 512893 363582
rect 512927 363548 512983 363582
rect 513017 363548 513073 363582
rect 513107 363548 513163 363582
rect 513197 363548 513329 363582
rect 512367 363529 513329 363548
rect 512367 363470 512439 363529
rect 512367 363436 512386 363470
rect 512420 363436 512439 363470
rect 513257 363504 513329 363529
rect 513257 363470 513276 363504
rect 513310 363470 513329 363504
rect 512367 363380 512439 363436
rect 512367 363346 512386 363380
rect 512420 363346 512439 363380
rect 512367 363290 512439 363346
rect 512367 363256 512386 363290
rect 512420 363256 512439 363290
rect 512367 363200 512439 363256
rect 512367 363166 512386 363200
rect 512420 363166 512439 363200
rect 512367 363110 512439 363166
rect 512367 363076 512386 363110
rect 512420 363076 512439 363110
rect 512367 363020 512439 363076
rect 512367 362986 512386 363020
rect 512420 362986 512439 363020
rect 512367 362930 512439 362986
rect 512367 362896 512386 362930
rect 512420 362896 512439 362930
rect 512367 362840 512439 362896
rect 512367 362806 512386 362840
rect 512420 362806 512439 362840
rect 512367 362750 512439 362806
rect 513257 363414 513329 363470
rect 513257 363380 513276 363414
rect 513310 363380 513329 363414
rect 513257 363324 513329 363380
rect 513257 363290 513276 363324
rect 513310 363290 513329 363324
rect 513257 363234 513329 363290
rect 513257 363200 513276 363234
rect 513310 363200 513329 363234
rect 513257 363144 513329 363200
rect 513257 363110 513276 363144
rect 513310 363110 513329 363144
rect 513257 363054 513329 363110
rect 513257 363020 513276 363054
rect 513310 363020 513329 363054
rect 513257 362964 513329 363020
rect 513257 362930 513276 362964
rect 513310 362930 513329 362964
rect 513257 362874 513329 362930
rect 513257 362840 513276 362874
rect 513310 362840 513329 362874
rect 513257 362784 513329 362840
rect 512367 362716 512386 362750
rect 512420 362716 512439 362750
rect 512367 362711 512439 362716
rect 513257 362750 513276 362784
rect 513310 362750 513329 362784
rect 513257 362711 513329 362750
rect 512367 362692 513329 362711
rect 512367 362658 512462 362692
rect 512496 362658 512552 362692
rect 512586 362658 512642 362692
rect 512676 362658 512732 362692
rect 512766 362658 512822 362692
rect 512856 362658 512912 362692
rect 512946 362658 513002 362692
rect 513036 362658 513092 362692
rect 513126 362658 513182 362692
rect 513216 362658 513329 362692
rect 512367 362639 513329 362658
rect 576214 359218 576334 359220
rect 576214 359182 576250 359218
rect 576294 359182 576334 359218
rect 576214 359180 576334 359182
rect 577514 359218 577634 359220
rect 577514 359182 577550 359218
rect 577594 359182 577634 359218
rect 577514 359180 577634 359182
rect 578814 359218 578934 359220
rect 578814 359182 578850 359218
rect 578894 359182 578934 359218
rect 578814 359180 578934 359182
rect 579952 359170 579992 359210
rect 579952 359090 579992 359130
rect 576662 313050 576782 313052
rect 576662 313014 576698 313050
rect 576742 313014 576782 313050
rect 576662 313012 576782 313014
rect 577962 313050 578082 313052
rect 577962 313014 577998 313050
rect 578042 313014 578082 313050
rect 577962 313012 578082 313014
rect 579262 313050 579382 313052
rect 579262 313014 579298 313050
rect 579342 313014 579382 313050
rect 579262 313012 579382 313014
rect 580400 313002 580440 313042
rect 580400 312922 580440 312962
<< psubdiffcont >>
rect 562184 492032 562228 492068
rect 563484 492032 563528 492068
rect 564784 492032 564828 492068
rect 565886 492060 565926 492100
rect 504742 402868 504776 402902
rect 504832 402868 504866 402902
rect 504922 402868 504956 402902
rect 505012 402868 505046 402902
rect 505102 402868 505136 402902
rect 505192 402868 505226 402902
rect 505282 402868 505316 402902
rect 505372 402868 505406 402902
rect 505462 402868 505496 402902
rect 505552 402868 505586 402902
rect 505642 402868 505676 402902
rect 505732 402868 505766 402902
rect 505822 402868 505856 402902
rect 560630 402918 560670 402958
rect 561728 402890 561772 402926
rect 563028 402890 563072 402926
rect 564328 402890 564372 402926
rect 504719 402772 504753 402806
rect 504719 402682 504753 402716
rect 504719 402592 504753 402626
rect 504719 402502 504753 402536
rect 504719 402412 504753 402446
rect 504719 402322 504753 402356
rect 504719 402232 504753 402266
rect 504719 402142 504753 402176
rect 504719 402052 504753 402086
rect 504719 401962 504753 401996
rect 504719 401872 504753 401906
rect 504719 401782 504753 401816
rect 505906 402772 505940 402806
rect 505906 402682 505940 402716
rect 505906 402592 505940 402626
rect 505906 402502 505940 402536
rect 505906 402412 505940 402446
rect 505906 402322 505940 402356
rect 505906 402232 505940 402266
rect 505906 402142 505940 402176
rect 505906 402052 505940 402086
rect 505906 401962 505940 401996
rect 505906 401872 505940 401906
rect 505906 401782 505940 401816
rect 504742 401681 504776 401715
rect 504832 401681 504866 401715
rect 504922 401681 504956 401715
rect 505012 401681 505046 401715
rect 505102 401681 505136 401715
rect 505192 401681 505226 401715
rect 505282 401681 505316 401715
rect 505372 401681 505406 401715
rect 505462 401681 505496 401715
rect 505552 401681 505586 401715
rect 505642 401681 505676 401715
rect 505732 401681 505766 401715
rect 505822 401681 505856 401715
rect 498591 400859 498625 400893
rect 505337 399835 505439 400277
rect 505337 397091 505439 397533
rect 512857 396993 512959 397435
rect 494057 392681 494159 393123
rect 505337 394059 505439 394501
rect 509097 394249 509199 394691
rect 512857 394249 512959 394691
rect 494831 391059 494865 391093
rect 505337 391015 505439 391457
rect 509097 391217 509199 391659
rect 512857 391505 512959 391947
rect 516617 391113 516719 391555
rect 506111 389559 506145 389593
rect 517391 389559 517425 389593
rect 506141 388457 506175 388491
rect 520377 389643 520479 390085
rect 517421 388457 517455 388491
rect 506141 387157 506175 387191
rect 512857 386311 512959 386753
rect 517421 387157 517455 387191
rect 520377 386311 520479 386753
rect 520377 383567 520479 384009
rect 520377 380333 520479 380775
rect 502351 377701 502385 377735
rect 502381 376599 502415 376633
rect 502381 375299 502415 375333
rect 516617 376119 516719 376561
rect 520377 376119 520479 376561
rect 500982 373076 501016 373110
rect 501072 373076 501106 373110
rect 501162 373076 501196 373110
rect 501252 373076 501286 373110
rect 501342 373076 501376 373110
rect 501432 373076 501466 373110
rect 501522 373076 501556 373110
rect 501612 373076 501646 373110
rect 501702 373076 501736 373110
rect 501792 373076 501826 373110
rect 501882 373076 501916 373110
rect 501972 373076 502006 373110
rect 502062 373076 502096 373110
rect 500959 372980 500993 373014
rect 500959 372890 500993 372924
rect 500959 372800 500993 372834
rect 500959 372710 500993 372744
rect 500959 372620 500993 372654
rect 500959 372530 500993 372564
rect 500959 372440 500993 372474
rect 500959 372350 500993 372384
rect 500959 372260 500993 372294
rect 500959 372170 500993 372204
rect 500959 372080 500993 372114
rect 500959 371990 500993 372024
rect 502146 372980 502180 373014
rect 502146 372890 502180 372924
rect 502146 372800 502180 372834
rect 502146 372710 502180 372744
rect 502146 372620 502180 372654
rect 502146 372530 502180 372564
rect 502146 372440 502180 372474
rect 502146 372350 502180 372384
rect 502146 372260 502180 372294
rect 502146 372170 502180 372204
rect 502146 372080 502180 372114
rect 497222 371900 497256 371934
rect 497312 371900 497346 371934
rect 497402 371900 497436 371934
rect 497492 371900 497526 371934
rect 497582 371900 497616 371934
rect 497672 371900 497706 371934
rect 497762 371900 497796 371934
rect 497852 371900 497886 371934
rect 497942 371900 497976 371934
rect 498032 371900 498066 371934
rect 498122 371900 498156 371934
rect 498212 371900 498246 371934
rect 498302 371900 498336 371934
rect 497199 371804 497233 371838
rect 497199 371714 497233 371748
rect 497199 371624 497233 371658
rect 497199 371534 497233 371568
rect 497199 371444 497233 371478
rect 497199 371354 497233 371388
rect 497199 371264 497233 371298
rect 497199 371174 497233 371208
rect 497199 371084 497233 371118
rect 497199 370994 497233 371028
rect 497199 370904 497233 370938
rect 497199 370814 497233 370848
rect 498386 371804 498420 371838
rect 498386 371714 498420 371748
rect 498386 371624 498420 371658
rect 498386 371534 498420 371568
rect 498386 371444 498420 371478
rect 498386 371354 498420 371388
rect 498386 371264 498420 371298
rect 498386 371174 498420 371208
rect 498386 371084 498420 371118
rect 498386 370994 498420 371028
rect 498386 370904 498420 370938
rect 498386 370814 498420 370848
rect 497222 370713 497256 370747
rect 497312 370713 497346 370747
rect 497402 370713 497436 370747
rect 497492 370713 497526 370747
rect 497582 370713 497616 370747
rect 497672 370713 497706 370747
rect 497762 370713 497796 370747
rect 497852 370713 497886 370747
rect 497942 370713 497976 370747
rect 498032 370713 498066 370747
rect 498122 370713 498156 370747
rect 498212 370713 498246 370747
rect 498302 370713 498336 370747
rect 497222 370560 497256 370594
rect 497312 370560 497346 370594
rect 497402 370560 497436 370594
rect 497492 370560 497526 370594
rect 497582 370560 497616 370594
rect 497672 370560 497706 370594
rect 497762 370560 497796 370594
rect 497852 370560 497886 370594
rect 497942 370560 497976 370594
rect 498032 370560 498066 370594
rect 498122 370560 498156 370594
rect 498212 370560 498246 370594
rect 498302 370560 498336 370594
rect 497199 370464 497233 370498
rect 497199 370374 497233 370408
rect 497199 370284 497233 370318
rect 497199 370194 497233 370228
rect 497199 370104 497233 370138
rect 497199 370014 497233 370048
rect 497199 369924 497233 369958
rect 497199 369834 497233 369868
rect 497199 369744 497233 369778
rect 497199 369654 497233 369688
rect 497199 369564 497233 369598
rect 497199 369474 497233 369508
rect 498386 370464 498420 370498
rect 498386 370374 498420 370408
rect 498386 370284 498420 370318
rect 498386 370194 498420 370228
rect 498386 370104 498420 370138
rect 498386 370014 498420 370048
rect 498386 369924 498420 369958
rect 498386 369834 498420 369868
rect 498386 369744 498420 369778
rect 498386 369654 498420 369688
rect 498386 369564 498420 369598
rect 498386 369474 498420 369508
rect 497222 369373 497256 369407
rect 497312 369373 497346 369407
rect 497402 369373 497436 369407
rect 497492 369373 497526 369407
rect 497582 369373 497616 369407
rect 497672 369373 497706 369407
rect 497762 369373 497796 369407
rect 497852 369373 497886 369407
rect 497942 369373 497976 369407
rect 498032 369373 498066 369407
rect 498122 369373 498156 369407
rect 498212 369373 498246 369407
rect 498302 369373 498336 369407
rect 497222 369220 497256 369254
rect 497312 369220 497346 369254
rect 497402 369220 497436 369254
rect 497492 369220 497526 369254
rect 497582 369220 497616 369254
rect 497672 369220 497706 369254
rect 497762 369220 497796 369254
rect 497852 369220 497886 369254
rect 497942 369220 497976 369254
rect 498032 369220 498066 369254
rect 498122 369220 498156 369254
rect 498212 369220 498246 369254
rect 498302 369220 498336 369254
rect 497199 369124 497233 369158
rect 497199 369034 497233 369068
rect 497199 368944 497233 368978
rect 497199 368854 497233 368888
rect 497199 368764 497233 368798
rect 497199 368674 497233 368708
rect 497199 368584 497233 368618
rect 497199 368494 497233 368528
rect 497199 368404 497233 368438
rect 497199 368314 497233 368348
rect 497199 368224 497233 368258
rect 497199 368134 497233 368168
rect 498386 369124 498420 369158
rect 498386 369034 498420 369068
rect 498386 368944 498420 368978
rect 498386 368854 498420 368888
rect 498386 368764 498420 368798
rect 498386 368674 498420 368708
rect 498386 368584 498420 368618
rect 498386 368494 498420 368528
rect 498386 368404 498420 368438
rect 498386 368314 498420 368348
rect 498386 368224 498420 368258
rect 498386 368134 498420 368168
rect 497222 368033 497256 368067
rect 497312 368033 497346 368067
rect 497402 368033 497436 368067
rect 497492 368033 497526 368067
rect 497582 368033 497616 368067
rect 497672 368033 497706 368067
rect 497762 368033 497796 368067
rect 497852 368033 497886 368067
rect 497942 368033 497976 368067
rect 498032 368033 498066 368067
rect 498122 368033 498156 368067
rect 498212 368033 498246 368067
rect 498302 368033 498336 368067
rect 497222 367880 497256 367914
rect 497312 367880 497346 367914
rect 497402 367880 497436 367914
rect 497492 367880 497526 367914
rect 497582 367880 497616 367914
rect 497672 367880 497706 367914
rect 497762 367880 497796 367914
rect 497852 367880 497886 367914
rect 497942 367880 497976 367914
rect 498032 367880 498066 367914
rect 498122 367880 498156 367914
rect 498212 367880 498246 367914
rect 498302 367880 498336 367914
rect 497199 367784 497233 367818
rect 497199 367694 497233 367728
rect 497199 367604 497233 367638
rect 497199 367514 497233 367548
rect 497199 367424 497233 367458
rect 497199 367334 497233 367368
rect 497199 367244 497233 367278
rect 497199 367154 497233 367188
rect 497199 367064 497233 367098
rect 497199 366974 497233 367008
rect 497199 366884 497233 366918
rect 497199 366794 497233 366828
rect 498386 367784 498420 367818
rect 498386 367694 498420 367728
rect 498386 367604 498420 367638
rect 498386 367514 498420 367548
rect 498386 367424 498420 367458
rect 498386 367334 498420 367368
rect 498386 367244 498420 367278
rect 498386 367154 498420 367188
rect 498386 367064 498420 367098
rect 498386 366974 498420 367008
rect 498386 366884 498420 366918
rect 498386 366794 498420 366828
rect 497222 366693 497256 366727
rect 497312 366693 497346 366727
rect 497402 366693 497436 366727
rect 497492 366693 497526 366727
rect 497582 366693 497616 366727
rect 497672 366693 497706 366727
rect 497762 366693 497796 366727
rect 497852 366693 497886 366727
rect 497942 366693 497976 366727
rect 498032 366693 498066 366727
rect 498122 366693 498156 366727
rect 498212 366693 498246 366727
rect 498302 366693 498336 366727
rect 497222 366540 497256 366574
rect 497312 366540 497346 366574
rect 497402 366540 497436 366574
rect 497492 366540 497526 366574
rect 497582 366540 497616 366574
rect 497672 366540 497706 366574
rect 497762 366540 497796 366574
rect 497852 366540 497886 366574
rect 497942 366540 497976 366574
rect 498032 366540 498066 366574
rect 498122 366540 498156 366574
rect 498212 366540 498246 366574
rect 498302 366540 498336 366574
rect 497199 366444 497233 366478
rect 497199 366354 497233 366388
rect 497199 366264 497233 366298
rect 497199 366174 497233 366208
rect 497199 366084 497233 366118
rect 497199 365994 497233 366028
rect 497199 365904 497233 365938
rect 497199 365814 497233 365848
rect 497199 365724 497233 365758
rect 497199 365634 497233 365668
rect 497199 365544 497233 365578
rect 497199 365454 497233 365488
rect 498386 366444 498420 366478
rect 498386 366354 498420 366388
rect 498386 366264 498420 366298
rect 498386 366174 498420 366208
rect 498386 366084 498420 366118
rect 498386 365994 498420 366028
rect 498386 365904 498420 365938
rect 498386 365814 498420 365848
rect 498386 365724 498420 365758
rect 498386 365634 498420 365668
rect 498386 365544 498420 365578
rect 498386 365454 498420 365488
rect 497222 365353 497256 365387
rect 497312 365353 497346 365387
rect 497402 365353 497436 365387
rect 497492 365353 497526 365387
rect 497582 365353 497616 365387
rect 497672 365353 497706 365387
rect 497762 365353 497796 365387
rect 497852 365353 497886 365387
rect 497942 365353 497976 365387
rect 498032 365353 498066 365387
rect 498122 365353 498156 365387
rect 498212 365353 498246 365387
rect 498302 365353 498336 365387
rect 497222 365200 497256 365234
rect 497312 365200 497346 365234
rect 497402 365200 497436 365234
rect 497492 365200 497526 365234
rect 497582 365200 497616 365234
rect 497672 365200 497706 365234
rect 497762 365200 497796 365234
rect 497852 365200 497886 365234
rect 497942 365200 497976 365234
rect 498032 365200 498066 365234
rect 498122 365200 498156 365234
rect 498212 365200 498246 365234
rect 498302 365200 498336 365234
rect 497199 365104 497233 365138
rect 497199 365014 497233 365048
rect 497199 364924 497233 364958
rect 497199 364834 497233 364868
rect 497199 364744 497233 364778
rect 497199 364654 497233 364688
rect 497199 364564 497233 364598
rect 497199 364474 497233 364508
rect 497199 364384 497233 364418
rect 497199 364294 497233 364328
rect 497199 364204 497233 364238
rect 497199 364114 497233 364148
rect 498386 365104 498420 365138
rect 498386 365014 498420 365048
rect 498386 364924 498420 364958
rect 498386 364834 498420 364868
rect 498386 364744 498420 364778
rect 498386 364654 498420 364688
rect 498386 364564 498420 364598
rect 498386 364474 498420 364508
rect 498386 364384 498420 364418
rect 498386 364294 498420 364328
rect 498386 364204 498420 364238
rect 498386 364114 498420 364148
rect 497222 364013 497256 364047
rect 497312 364013 497346 364047
rect 497402 364013 497436 364047
rect 497492 364013 497526 364047
rect 497582 364013 497616 364047
rect 497672 364013 497706 364047
rect 497762 364013 497796 364047
rect 497852 364013 497886 364047
rect 497942 364013 497976 364047
rect 498032 364013 498066 364047
rect 498122 364013 498156 364047
rect 498212 364013 498246 364047
rect 498302 364013 498336 364047
rect 497222 363860 497256 363894
rect 497312 363860 497346 363894
rect 497402 363860 497436 363894
rect 497492 363860 497526 363894
rect 497582 363860 497616 363894
rect 497672 363860 497706 363894
rect 497762 363860 497796 363894
rect 497852 363860 497886 363894
rect 497942 363860 497976 363894
rect 498032 363860 498066 363894
rect 498122 363860 498156 363894
rect 498212 363860 498246 363894
rect 498302 363860 498336 363894
rect 497199 363764 497233 363798
rect 497199 363674 497233 363708
rect 497199 363584 497233 363618
rect 497199 363494 497233 363528
rect 497199 363404 497233 363438
rect 497199 363314 497233 363348
rect 497199 363224 497233 363258
rect 497199 363134 497233 363168
rect 497199 363044 497233 363078
rect 497199 362954 497233 362988
rect 497199 362864 497233 362898
rect 497199 362774 497233 362808
rect 498386 363764 498420 363798
rect 498386 363674 498420 363708
rect 498386 363584 498420 363618
rect 498386 363494 498420 363528
rect 498386 363404 498420 363438
rect 498386 363314 498420 363348
rect 498386 363224 498420 363258
rect 498386 363134 498420 363168
rect 498386 363044 498420 363078
rect 498386 362954 498420 362988
rect 498386 362864 498420 362898
rect 498386 362774 498420 362808
rect 497222 362673 497256 362707
rect 497312 362673 497346 362707
rect 497402 362673 497436 362707
rect 497492 362673 497526 362707
rect 497582 362673 497616 362707
rect 497672 362673 497706 362707
rect 497762 362673 497796 362707
rect 497852 362673 497886 362707
rect 497942 362673 497976 362707
rect 498032 362673 498066 362707
rect 498122 362673 498156 362707
rect 498212 362673 498246 362707
rect 498302 362673 498336 362707
rect 502146 371990 502180 372024
rect 500982 371889 501016 371923
rect 501072 371889 501106 371923
rect 501162 371889 501196 371923
rect 501252 371889 501286 371923
rect 501342 371889 501376 371923
rect 501432 371889 501466 371923
rect 501522 371889 501556 371923
rect 501612 371889 501646 371923
rect 501702 371889 501736 371923
rect 501792 371889 501826 371923
rect 501882 371889 501916 371923
rect 501972 371889 502006 371923
rect 502062 371889 502096 371923
rect 500982 371736 501016 371770
rect 501072 371736 501106 371770
rect 501162 371736 501196 371770
rect 501252 371736 501286 371770
rect 501342 371736 501376 371770
rect 501432 371736 501466 371770
rect 501522 371736 501556 371770
rect 501612 371736 501646 371770
rect 501702 371736 501736 371770
rect 501792 371736 501826 371770
rect 501882 371736 501916 371770
rect 501972 371736 502006 371770
rect 502062 371736 502096 371770
rect 500959 371640 500993 371674
rect 500959 371550 500993 371584
rect 500959 371460 500993 371494
rect 500959 371370 500993 371404
rect 500959 371280 500993 371314
rect 500959 371190 500993 371224
rect 500959 371100 500993 371134
rect 500959 371010 500993 371044
rect 500959 370920 500993 370954
rect 500959 370830 500993 370864
rect 500959 370740 500993 370774
rect 500959 370650 500993 370684
rect 502146 371640 502180 371674
rect 502146 371550 502180 371584
rect 502146 371460 502180 371494
rect 502146 371370 502180 371404
rect 502146 371280 502180 371314
rect 502146 371190 502180 371224
rect 502146 371100 502180 371134
rect 502146 371010 502180 371044
rect 502146 370920 502180 370954
rect 502146 370830 502180 370864
rect 502146 370740 502180 370774
rect 502146 370650 502180 370684
rect 500982 370549 501016 370583
rect 501072 370549 501106 370583
rect 501162 370549 501196 370583
rect 501252 370549 501286 370583
rect 501342 370549 501376 370583
rect 501432 370549 501466 370583
rect 501522 370549 501556 370583
rect 501612 370549 501646 370583
rect 501702 370549 501736 370583
rect 501792 370549 501826 370583
rect 501882 370549 501916 370583
rect 501972 370549 502006 370583
rect 502062 370549 502096 370583
rect 500982 370396 501016 370430
rect 501072 370396 501106 370430
rect 501162 370396 501196 370430
rect 501252 370396 501286 370430
rect 501342 370396 501376 370430
rect 501432 370396 501466 370430
rect 501522 370396 501556 370430
rect 501612 370396 501646 370430
rect 501702 370396 501736 370430
rect 501792 370396 501826 370430
rect 501882 370396 501916 370430
rect 501972 370396 502006 370430
rect 502062 370396 502096 370430
rect 500959 370300 500993 370334
rect 500959 370210 500993 370244
rect 500959 370120 500993 370154
rect 500959 370030 500993 370064
rect 500959 369940 500993 369974
rect 500959 369850 500993 369884
rect 500959 369760 500993 369794
rect 500959 369670 500993 369704
rect 500959 369580 500993 369614
rect 500959 369490 500993 369524
rect 500959 369400 500993 369434
rect 500959 369310 500993 369344
rect 502146 370300 502180 370334
rect 502146 370210 502180 370244
rect 502146 370120 502180 370154
rect 502146 370030 502180 370064
rect 502146 369940 502180 369974
rect 502146 369850 502180 369884
rect 502146 369760 502180 369794
rect 502146 369670 502180 369704
rect 502146 369580 502180 369614
rect 502146 369490 502180 369524
rect 502146 369400 502180 369434
rect 502146 369310 502180 369344
rect 500982 369209 501016 369243
rect 501072 369209 501106 369243
rect 501162 369209 501196 369243
rect 501252 369209 501286 369243
rect 501342 369209 501376 369243
rect 501432 369209 501466 369243
rect 501522 369209 501556 369243
rect 501612 369209 501646 369243
rect 501702 369209 501736 369243
rect 501792 369209 501826 369243
rect 501882 369209 501916 369243
rect 501972 369209 502006 369243
rect 502062 369209 502096 369243
rect 500982 369056 501016 369090
rect 501072 369056 501106 369090
rect 501162 369056 501196 369090
rect 501252 369056 501286 369090
rect 501342 369056 501376 369090
rect 501432 369056 501466 369090
rect 501522 369056 501556 369090
rect 501612 369056 501646 369090
rect 501702 369056 501736 369090
rect 501792 369056 501826 369090
rect 501882 369056 501916 369090
rect 501972 369056 502006 369090
rect 502062 369056 502096 369090
rect 500959 368960 500993 368994
rect 500959 368870 500993 368904
rect 500959 368780 500993 368814
rect 500959 368690 500993 368724
rect 500959 368600 500993 368634
rect 500959 368510 500993 368544
rect 500959 368420 500993 368454
rect 500959 368330 500993 368364
rect 500959 368240 500993 368274
rect 500959 368150 500993 368184
rect 500959 368060 500993 368094
rect 500959 367970 500993 368004
rect 502146 368960 502180 368994
rect 502146 368870 502180 368904
rect 502146 368780 502180 368814
rect 502146 368690 502180 368724
rect 502146 368600 502180 368634
rect 502146 368510 502180 368544
rect 502146 368420 502180 368454
rect 502146 368330 502180 368364
rect 502146 368240 502180 368274
rect 502146 368150 502180 368184
rect 502146 368060 502180 368094
rect 502146 367970 502180 368004
rect 500982 367869 501016 367903
rect 501072 367869 501106 367903
rect 501162 367869 501196 367903
rect 501252 367869 501286 367903
rect 501342 367869 501376 367903
rect 501432 367869 501466 367903
rect 501522 367869 501556 367903
rect 501612 367869 501646 367903
rect 501702 367869 501736 367903
rect 501792 367869 501826 367903
rect 501882 367869 501916 367903
rect 501972 367869 502006 367903
rect 502062 367869 502096 367903
rect 500982 367716 501016 367750
rect 501072 367716 501106 367750
rect 501162 367716 501196 367750
rect 501252 367716 501286 367750
rect 501342 367716 501376 367750
rect 501432 367716 501466 367750
rect 501522 367716 501556 367750
rect 501612 367716 501646 367750
rect 501702 367716 501736 367750
rect 501792 367716 501826 367750
rect 501882 367716 501916 367750
rect 501972 367716 502006 367750
rect 502062 367716 502096 367750
rect 500959 367620 500993 367654
rect 500959 367530 500993 367564
rect 500959 367440 500993 367474
rect 500959 367350 500993 367384
rect 500959 367260 500993 367294
rect 500959 367170 500993 367204
rect 500959 367080 500993 367114
rect 500959 366990 500993 367024
rect 500959 366900 500993 366934
rect 500959 366810 500993 366844
rect 500959 366720 500993 366754
rect 500959 366630 500993 366664
rect 502146 367620 502180 367654
rect 502146 367530 502180 367564
rect 502146 367440 502180 367474
rect 502146 367350 502180 367384
rect 502146 367260 502180 367294
rect 502146 367170 502180 367204
rect 502146 367080 502180 367114
rect 502146 366990 502180 367024
rect 502146 366900 502180 366934
rect 502146 366810 502180 366844
rect 502146 366720 502180 366754
rect 502146 366630 502180 366664
rect 500982 366529 501016 366563
rect 501072 366529 501106 366563
rect 501162 366529 501196 366563
rect 501252 366529 501286 366563
rect 501342 366529 501376 366563
rect 501432 366529 501466 366563
rect 501522 366529 501556 366563
rect 501612 366529 501646 366563
rect 501702 366529 501736 366563
rect 501792 366529 501826 366563
rect 501882 366529 501916 366563
rect 501972 366529 502006 366563
rect 502062 366529 502096 366563
rect 500982 366376 501016 366410
rect 501072 366376 501106 366410
rect 501162 366376 501196 366410
rect 501252 366376 501286 366410
rect 501342 366376 501376 366410
rect 501432 366376 501466 366410
rect 501522 366376 501556 366410
rect 501612 366376 501646 366410
rect 501702 366376 501736 366410
rect 501792 366376 501826 366410
rect 501882 366376 501916 366410
rect 501972 366376 502006 366410
rect 502062 366376 502096 366410
rect 500959 366280 500993 366314
rect 500959 366190 500993 366224
rect 500959 366100 500993 366134
rect 500959 366010 500993 366044
rect 500959 365920 500993 365954
rect 500959 365830 500993 365864
rect 500959 365740 500993 365774
rect 500959 365650 500993 365684
rect 500959 365560 500993 365594
rect 500959 365470 500993 365504
rect 500959 365380 500993 365414
rect 500959 365290 500993 365324
rect 502146 366280 502180 366314
rect 502146 366190 502180 366224
rect 502146 366100 502180 366134
rect 502146 366010 502180 366044
rect 502146 365920 502180 365954
rect 502146 365830 502180 365864
rect 502146 365740 502180 365774
rect 502146 365650 502180 365684
rect 502146 365560 502180 365594
rect 502146 365470 502180 365504
rect 502146 365380 502180 365414
rect 502146 365290 502180 365324
rect 500982 365189 501016 365223
rect 501072 365189 501106 365223
rect 501162 365189 501196 365223
rect 501252 365189 501286 365223
rect 501342 365189 501376 365223
rect 501432 365189 501466 365223
rect 501522 365189 501556 365223
rect 501612 365189 501646 365223
rect 501702 365189 501736 365223
rect 501792 365189 501826 365223
rect 501882 365189 501916 365223
rect 501972 365189 502006 365223
rect 502062 365189 502096 365223
rect 500982 365036 501016 365070
rect 501072 365036 501106 365070
rect 501162 365036 501196 365070
rect 501252 365036 501286 365070
rect 501342 365036 501376 365070
rect 501432 365036 501466 365070
rect 501522 365036 501556 365070
rect 501612 365036 501646 365070
rect 501702 365036 501736 365070
rect 501792 365036 501826 365070
rect 501882 365036 501916 365070
rect 501972 365036 502006 365070
rect 502062 365036 502096 365070
rect 500959 364940 500993 364974
rect 500959 364850 500993 364884
rect 500959 364760 500993 364794
rect 500959 364670 500993 364704
rect 500959 364580 500993 364614
rect 500959 364490 500993 364524
rect 500959 364400 500993 364434
rect 500959 364310 500993 364344
rect 500959 364220 500993 364254
rect 500959 364130 500993 364164
rect 500959 364040 500993 364074
rect 500959 363950 500993 363984
rect 502146 364940 502180 364974
rect 502146 364850 502180 364884
rect 502146 364760 502180 364794
rect 502146 364670 502180 364704
rect 502146 364580 502180 364614
rect 502146 364490 502180 364524
rect 502146 364400 502180 364434
rect 502146 364310 502180 364344
rect 502146 364220 502180 364254
rect 502146 364130 502180 364164
rect 502146 364040 502180 364074
rect 502146 363950 502180 363984
rect 500982 363849 501016 363883
rect 501072 363849 501106 363883
rect 501162 363849 501196 363883
rect 501252 363849 501286 363883
rect 501342 363849 501376 363883
rect 501432 363849 501466 363883
rect 501522 363849 501556 363883
rect 501612 363849 501646 363883
rect 501702 363849 501736 363883
rect 501792 363849 501826 363883
rect 501882 363849 501916 363883
rect 501972 363849 502006 363883
rect 502062 363849 502096 363883
rect 500982 363696 501016 363730
rect 501072 363696 501106 363730
rect 501162 363696 501196 363730
rect 501252 363696 501286 363730
rect 501342 363696 501376 363730
rect 501432 363696 501466 363730
rect 501522 363696 501556 363730
rect 501612 363696 501646 363730
rect 501702 363696 501736 363730
rect 501792 363696 501826 363730
rect 501882 363696 501916 363730
rect 501972 363696 502006 363730
rect 502062 363696 502096 363730
rect 500959 363600 500993 363634
rect 500959 363510 500993 363544
rect 500959 363420 500993 363454
rect 500959 363330 500993 363364
rect 500959 363240 500993 363274
rect 500959 363150 500993 363184
rect 500959 363060 500993 363094
rect 500959 362970 500993 363004
rect 500959 362880 500993 362914
rect 500959 362790 500993 362824
rect 500959 362700 500993 362734
rect 500959 362610 500993 362644
rect 502146 363600 502180 363634
rect 502146 363510 502180 363544
rect 502146 363420 502180 363454
rect 502146 363330 502180 363364
rect 502146 363240 502180 363274
rect 502146 363150 502180 363184
rect 502146 363060 502180 363094
rect 502146 362970 502180 363004
rect 502146 362880 502180 362914
rect 502146 362790 502180 362824
rect 502146 362700 502180 362734
rect 502146 362610 502180 362644
rect 500982 362509 501016 362543
rect 501072 362509 501106 362543
rect 501162 362509 501196 362543
rect 501252 362509 501286 362543
rect 501342 362509 501376 362543
rect 501432 362509 501466 362543
rect 501522 362509 501556 362543
rect 501612 362509 501646 362543
rect 501702 362509 501736 362543
rect 501792 362509 501826 362543
rect 501882 362509 501916 362543
rect 501972 362509 502006 362543
rect 502062 362509 502096 362543
rect 504742 373076 504776 373110
rect 504832 373076 504866 373110
rect 504922 373076 504956 373110
rect 505012 373076 505046 373110
rect 505102 373076 505136 373110
rect 505192 373076 505226 373110
rect 505282 373076 505316 373110
rect 505372 373076 505406 373110
rect 505462 373076 505496 373110
rect 505552 373076 505586 373110
rect 505642 373076 505676 373110
rect 505732 373076 505766 373110
rect 505822 373076 505856 373110
rect 504719 372980 504753 373014
rect 504719 372890 504753 372924
rect 504719 372800 504753 372834
rect 504719 372710 504753 372744
rect 504719 372620 504753 372654
rect 504719 372530 504753 372564
rect 504719 372440 504753 372474
rect 504719 372350 504753 372384
rect 504719 372260 504753 372294
rect 504719 372170 504753 372204
rect 504719 372080 504753 372114
rect 504719 371990 504753 372024
rect 505906 372980 505940 373014
rect 505906 372890 505940 372924
rect 505906 372800 505940 372834
rect 505906 372710 505940 372744
rect 505906 372620 505940 372654
rect 505906 372530 505940 372564
rect 505906 372440 505940 372474
rect 505906 372350 505940 372384
rect 505906 372260 505940 372294
rect 505906 372170 505940 372204
rect 505906 372080 505940 372114
rect 505906 371990 505940 372024
rect 504742 371889 504776 371923
rect 504832 371889 504866 371923
rect 504922 371889 504956 371923
rect 505012 371889 505046 371923
rect 505102 371889 505136 371923
rect 505192 371889 505226 371923
rect 505282 371889 505316 371923
rect 505372 371889 505406 371923
rect 505462 371889 505496 371923
rect 505552 371889 505586 371923
rect 505642 371889 505676 371923
rect 505732 371889 505766 371923
rect 505822 371889 505856 371923
rect 504742 371736 504776 371770
rect 504832 371736 504866 371770
rect 504922 371736 504956 371770
rect 505012 371736 505046 371770
rect 505102 371736 505136 371770
rect 505192 371736 505226 371770
rect 505282 371736 505316 371770
rect 505372 371736 505406 371770
rect 505462 371736 505496 371770
rect 505552 371736 505586 371770
rect 505642 371736 505676 371770
rect 505732 371736 505766 371770
rect 505822 371736 505856 371770
rect 504719 371640 504753 371674
rect 504719 371550 504753 371584
rect 504719 371460 504753 371494
rect 504719 371370 504753 371404
rect 504719 371280 504753 371314
rect 504719 371190 504753 371224
rect 504719 371100 504753 371134
rect 504719 371010 504753 371044
rect 504719 370920 504753 370954
rect 504719 370830 504753 370864
rect 504719 370740 504753 370774
rect 504719 370650 504753 370684
rect 505906 371640 505940 371674
rect 505906 371550 505940 371584
rect 505906 371460 505940 371494
rect 505906 371370 505940 371404
rect 505906 371280 505940 371314
rect 505906 371190 505940 371224
rect 505906 371100 505940 371134
rect 505906 371010 505940 371044
rect 505906 370920 505940 370954
rect 505906 370830 505940 370864
rect 505906 370740 505940 370774
rect 505906 370650 505940 370684
rect 504742 370549 504776 370583
rect 504832 370549 504866 370583
rect 504922 370549 504956 370583
rect 505012 370549 505046 370583
rect 505102 370549 505136 370583
rect 505192 370549 505226 370583
rect 505282 370549 505316 370583
rect 505372 370549 505406 370583
rect 505462 370549 505496 370583
rect 505552 370549 505586 370583
rect 505642 370549 505676 370583
rect 505732 370549 505766 370583
rect 505822 370549 505856 370583
rect 504742 370396 504776 370430
rect 504832 370396 504866 370430
rect 504922 370396 504956 370430
rect 505012 370396 505046 370430
rect 505102 370396 505136 370430
rect 505192 370396 505226 370430
rect 505282 370396 505316 370430
rect 505372 370396 505406 370430
rect 505462 370396 505496 370430
rect 505552 370396 505586 370430
rect 505642 370396 505676 370430
rect 505732 370396 505766 370430
rect 505822 370396 505856 370430
rect 504719 370300 504753 370334
rect 504719 370210 504753 370244
rect 504719 370120 504753 370154
rect 504719 370030 504753 370064
rect 504719 369940 504753 369974
rect 504719 369850 504753 369884
rect 504719 369760 504753 369794
rect 504719 369670 504753 369704
rect 504719 369580 504753 369614
rect 504719 369490 504753 369524
rect 504719 369400 504753 369434
rect 504719 369310 504753 369344
rect 505906 370300 505940 370334
rect 505906 370210 505940 370244
rect 505906 370120 505940 370154
rect 505906 370030 505940 370064
rect 505906 369940 505940 369974
rect 505906 369850 505940 369884
rect 505906 369760 505940 369794
rect 505906 369670 505940 369704
rect 505906 369580 505940 369614
rect 505906 369490 505940 369524
rect 505906 369400 505940 369434
rect 505906 369310 505940 369344
rect 504742 369209 504776 369243
rect 504832 369209 504866 369243
rect 504922 369209 504956 369243
rect 505012 369209 505046 369243
rect 505102 369209 505136 369243
rect 505192 369209 505226 369243
rect 505282 369209 505316 369243
rect 505372 369209 505406 369243
rect 505462 369209 505496 369243
rect 505552 369209 505586 369243
rect 505642 369209 505676 369243
rect 505732 369209 505766 369243
rect 505822 369209 505856 369243
rect 504742 369056 504776 369090
rect 504832 369056 504866 369090
rect 504922 369056 504956 369090
rect 505012 369056 505046 369090
rect 505102 369056 505136 369090
rect 505192 369056 505226 369090
rect 505282 369056 505316 369090
rect 505372 369056 505406 369090
rect 505462 369056 505496 369090
rect 505552 369056 505586 369090
rect 505642 369056 505676 369090
rect 505732 369056 505766 369090
rect 505822 369056 505856 369090
rect 504719 368960 504753 368994
rect 504719 368870 504753 368904
rect 504719 368780 504753 368814
rect 504719 368690 504753 368724
rect 504719 368600 504753 368634
rect 504719 368510 504753 368544
rect 504719 368420 504753 368454
rect 504719 368330 504753 368364
rect 504719 368240 504753 368274
rect 504719 368150 504753 368184
rect 504719 368060 504753 368094
rect 504719 367970 504753 368004
rect 505906 368960 505940 368994
rect 505906 368870 505940 368904
rect 505906 368780 505940 368814
rect 505906 368690 505940 368724
rect 505906 368600 505940 368634
rect 505906 368510 505940 368544
rect 505906 368420 505940 368454
rect 505906 368330 505940 368364
rect 505906 368240 505940 368274
rect 505906 368150 505940 368184
rect 505906 368060 505940 368094
rect 505906 367970 505940 368004
rect 504742 367869 504776 367903
rect 504832 367869 504866 367903
rect 504922 367869 504956 367903
rect 505012 367869 505046 367903
rect 505102 367869 505136 367903
rect 505192 367869 505226 367903
rect 505282 367869 505316 367903
rect 505372 367869 505406 367903
rect 505462 367869 505496 367903
rect 505552 367869 505586 367903
rect 505642 367869 505676 367903
rect 505732 367869 505766 367903
rect 505822 367869 505856 367903
rect 504742 367716 504776 367750
rect 504832 367716 504866 367750
rect 504922 367716 504956 367750
rect 505012 367716 505046 367750
rect 505102 367716 505136 367750
rect 505192 367716 505226 367750
rect 505282 367716 505316 367750
rect 505372 367716 505406 367750
rect 505462 367716 505496 367750
rect 505552 367716 505586 367750
rect 505642 367716 505676 367750
rect 505732 367716 505766 367750
rect 505822 367716 505856 367750
rect 504719 367620 504753 367654
rect 504719 367530 504753 367564
rect 504719 367440 504753 367474
rect 504719 367350 504753 367384
rect 504719 367260 504753 367294
rect 504719 367170 504753 367204
rect 504719 367080 504753 367114
rect 504719 366990 504753 367024
rect 504719 366900 504753 366934
rect 504719 366810 504753 366844
rect 504719 366720 504753 366754
rect 504719 366630 504753 366664
rect 505906 367620 505940 367654
rect 505906 367530 505940 367564
rect 505906 367440 505940 367474
rect 505906 367350 505940 367384
rect 505906 367260 505940 367294
rect 505906 367170 505940 367204
rect 505906 367080 505940 367114
rect 505906 366990 505940 367024
rect 505906 366900 505940 366934
rect 505906 366810 505940 366844
rect 505906 366720 505940 366754
rect 505906 366630 505940 366664
rect 504742 366529 504776 366563
rect 504832 366529 504866 366563
rect 504922 366529 504956 366563
rect 505012 366529 505046 366563
rect 505102 366529 505136 366563
rect 505192 366529 505226 366563
rect 505282 366529 505316 366563
rect 505372 366529 505406 366563
rect 505462 366529 505496 366563
rect 505552 366529 505586 366563
rect 505642 366529 505676 366563
rect 505732 366529 505766 366563
rect 505822 366529 505856 366563
rect 504742 366376 504776 366410
rect 504832 366376 504866 366410
rect 504922 366376 504956 366410
rect 505012 366376 505046 366410
rect 505102 366376 505136 366410
rect 505192 366376 505226 366410
rect 505282 366376 505316 366410
rect 505372 366376 505406 366410
rect 505462 366376 505496 366410
rect 505552 366376 505586 366410
rect 505642 366376 505676 366410
rect 505732 366376 505766 366410
rect 505822 366376 505856 366410
rect 504719 366280 504753 366314
rect 504719 366190 504753 366224
rect 504719 366100 504753 366134
rect 504719 366010 504753 366044
rect 504719 365920 504753 365954
rect 504719 365830 504753 365864
rect 504719 365740 504753 365774
rect 504719 365650 504753 365684
rect 504719 365560 504753 365594
rect 504719 365470 504753 365504
rect 504719 365380 504753 365414
rect 504719 365290 504753 365324
rect 505906 366280 505940 366314
rect 505906 366190 505940 366224
rect 505906 366100 505940 366134
rect 505906 366010 505940 366044
rect 505906 365920 505940 365954
rect 505906 365830 505940 365864
rect 505906 365740 505940 365774
rect 505906 365650 505940 365684
rect 505906 365560 505940 365594
rect 505906 365470 505940 365504
rect 505906 365380 505940 365414
rect 505906 365290 505940 365324
rect 504742 365189 504776 365223
rect 504832 365189 504866 365223
rect 504922 365189 504956 365223
rect 505012 365189 505046 365223
rect 505102 365189 505136 365223
rect 505192 365189 505226 365223
rect 505282 365189 505316 365223
rect 505372 365189 505406 365223
rect 505462 365189 505496 365223
rect 505552 365189 505586 365223
rect 505642 365189 505676 365223
rect 505732 365189 505766 365223
rect 505822 365189 505856 365223
rect 504742 365036 504776 365070
rect 504832 365036 504866 365070
rect 504922 365036 504956 365070
rect 505012 365036 505046 365070
rect 505102 365036 505136 365070
rect 505192 365036 505226 365070
rect 505282 365036 505316 365070
rect 505372 365036 505406 365070
rect 505462 365036 505496 365070
rect 505552 365036 505586 365070
rect 505642 365036 505676 365070
rect 505732 365036 505766 365070
rect 505822 365036 505856 365070
rect 504719 364940 504753 364974
rect 504719 364850 504753 364884
rect 504719 364760 504753 364794
rect 504719 364670 504753 364704
rect 504719 364580 504753 364614
rect 504719 364490 504753 364524
rect 504719 364400 504753 364434
rect 504719 364310 504753 364344
rect 504719 364220 504753 364254
rect 504719 364130 504753 364164
rect 504719 364040 504753 364074
rect 504719 363950 504753 363984
rect 505906 364940 505940 364974
rect 505906 364850 505940 364884
rect 505906 364760 505940 364794
rect 505906 364670 505940 364704
rect 505906 364580 505940 364614
rect 505906 364490 505940 364524
rect 505906 364400 505940 364434
rect 505906 364310 505940 364344
rect 505906 364220 505940 364254
rect 505906 364130 505940 364164
rect 505906 364040 505940 364074
rect 505906 363950 505940 363984
rect 504742 363849 504776 363883
rect 504832 363849 504866 363883
rect 504922 363849 504956 363883
rect 505012 363849 505046 363883
rect 505102 363849 505136 363883
rect 505192 363849 505226 363883
rect 505282 363849 505316 363883
rect 505372 363849 505406 363883
rect 505462 363849 505496 363883
rect 505552 363849 505586 363883
rect 505642 363849 505676 363883
rect 505732 363849 505766 363883
rect 505822 363849 505856 363883
rect 504742 363696 504776 363730
rect 504832 363696 504866 363730
rect 504922 363696 504956 363730
rect 505012 363696 505046 363730
rect 505102 363696 505136 363730
rect 505192 363696 505226 363730
rect 505282 363696 505316 363730
rect 505372 363696 505406 363730
rect 505462 363696 505496 363730
rect 505552 363696 505586 363730
rect 505642 363696 505676 363730
rect 505732 363696 505766 363730
rect 505822 363696 505856 363730
rect 504719 363600 504753 363634
rect 504719 363510 504753 363544
rect 504719 363420 504753 363454
rect 504719 363330 504753 363364
rect 504719 363240 504753 363274
rect 504719 363150 504753 363184
rect 504719 363060 504753 363094
rect 504719 362970 504753 363004
rect 504719 362880 504753 362914
rect 504719 362790 504753 362824
rect 504719 362700 504753 362734
rect 504719 362610 504753 362644
rect 505906 363600 505940 363634
rect 505906 363510 505940 363544
rect 505906 363420 505940 363454
rect 505906 363330 505940 363364
rect 505906 363240 505940 363274
rect 505906 363150 505940 363184
rect 505906 363060 505940 363094
rect 505906 362970 505940 363004
rect 505906 362880 505940 362914
rect 505906 362790 505940 362824
rect 505906 362700 505940 362734
rect 505906 362610 505940 362644
rect 504742 362509 504776 362543
rect 504832 362509 504866 362543
rect 504922 362509 504956 362543
rect 505012 362509 505046 362543
rect 505102 362509 505136 362543
rect 505192 362509 505226 362543
rect 505282 362509 505316 362543
rect 505372 362509 505406 362543
rect 505462 362509 505496 362543
rect 505552 362509 505586 362543
rect 505642 362509 505676 362543
rect 505732 362509 505766 362543
rect 505822 362509 505856 362543
rect 508502 373076 508536 373110
rect 508592 373076 508626 373110
rect 508682 373076 508716 373110
rect 508772 373076 508806 373110
rect 508862 373076 508896 373110
rect 508952 373076 508986 373110
rect 509042 373076 509076 373110
rect 509132 373076 509166 373110
rect 509222 373076 509256 373110
rect 509312 373076 509346 373110
rect 509402 373076 509436 373110
rect 509492 373076 509526 373110
rect 509582 373076 509616 373110
rect 508479 372980 508513 373014
rect 508479 372890 508513 372924
rect 508479 372800 508513 372834
rect 508479 372710 508513 372744
rect 508479 372620 508513 372654
rect 508479 372530 508513 372564
rect 508479 372440 508513 372474
rect 508479 372350 508513 372384
rect 508479 372260 508513 372294
rect 508479 372170 508513 372204
rect 508479 372080 508513 372114
rect 508479 371990 508513 372024
rect 509666 372980 509700 373014
rect 509666 372890 509700 372924
rect 509666 372800 509700 372834
rect 509666 372710 509700 372744
rect 509666 372620 509700 372654
rect 509666 372530 509700 372564
rect 509666 372440 509700 372474
rect 509666 372350 509700 372384
rect 509666 372260 509700 372294
rect 509666 372170 509700 372204
rect 509666 372080 509700 372114
rect 509666 371990 509700 372024
rect 508502 371889 508536 371923
rect 508592 371889 508626 371923
rect 508682 371889 508716 371923
rect 508772 371889 508806 371923
rect 508862 371889 508896 371923
rect 508952 371889 508986 371923
rect 509042 371889 509076 371923
rect 509132 371889 509166 371923
rect 509222 371889 509256 371923
rect 509312 371889 509346 371923
rect 509402 371889 509436 371923
rect 509492 371889 509526 371923
rect 509582 371889 509616 371923
rect 508502 371736 508536 371770
rect 508592 371736 508626 371770
rect 508682 371736 508716 371770
rect 508772 371736 508806 371770
rect 508862 371736 508896 371770
rect 508952 371736 508986 371770
rect 509042 371736 509076 371770
rect 509132 371736 509166 371770
rect 509222 371736 509256 371770
rect 509312 371736 509346 371770
rect 509402 371736 509436 371770
rect 509492 371736 509526 371770
rect 509582 371736 509616 371770
rect 508479 371640 508513 371674
rect 508479 371550 508513 371584
rect 508479 371460 508513 371494
rect 508479 371370 508513 371404
rect 508479 371280 508513 371314
rect 508479 371190 508513 371224
rect 508479 371100 508513 371134
rect 508479 371010 508513 371044
rect 508479 370920 508513 370954
rect 508479 370830 508513 370864
rect 508479 370740 508513 370774
rect 508479 370650 508513 370684
rect 509666 371640 509700 371674
rect 509666 371550 509700 371584
rect 509666 371460 509700 371494
rect 509666 371370 509700 371404
rect 509666 371280 509700 371314
rect 509666 371190 509700 371224
rect 509666 371100 509700 371134
rect 509666 371010 509700 371044
rect 509666 370920 509700 370954
rect 509666 370830 509700 370864
rect 509666 370740 509700 370774
rect 509666 370650 509700 370684
rect 508502 370549 508536 370583
rect 508592 370549 508626 370583
rect 508682 370549 508716 370583
rect 508772 370549 508806 370583
rect 508862 370549 508896 370583
rect 508952 370549 508986 370583
rect 509042 370549 509076 370583
rect 509132 370549 509166 370583
rect 509222 370549 509256 370583
rect 509312 370549 509346 370583
rect 509402 370549 509436 370583
rect 509492 370549 509526 370583
rect 509582 370549 509616 370583
rect 508502 370396 508536 370430
rect 508592 370396 508626 370430
rect 508682 370396 508716 370430
rect 508772 370396 508806 370430
rect 508862 370396 508896 370430
rect 508952 370396 508986 370430
rect 509042 370396 509076 370430
rect 509132 370396 509166 370430
rect 509222 370396 509256 370430
rect 509312 370396 509346 370430
rect 509402 370396 509436 370430
rect 509492 370396 509526 370430
rect 509582 370396 509616 370430
rect 508479 370300 508513 370334
rect 508479 370210 508513 370244
rect 508479 370120 508513 370154
rect 508479 370030 508513 370064
rect 508479 369940 508513 369974
rect 508479 369850 508513 369884
rect 508479 369760 508513 369794
rect 508479 369670 508513 369704
rect 508479 369580 508513 369614
rect 508479 369490 508513 369524
rect 508479 369400 508513 369434
rect 508479 369310 508513 369344
rect 509666 370300 509700 370334
rect 509666 370210 509700 370244
rect 509666 370120 509700 370154
rect 509666 370030 509700 370064
rect 509666 369940 509700 369974
rect 509666 369850 509700 369884
rect 509666 369760 509700 369794
rect 509666 369670 509700 369704
rect 509666 369580 509700 369614
rect 509666 369490 509700 369524
rect 509666 369400 509700 369434
rect 509666 369310 509700 369344
rect 508502 369209 508536 369243
rect 508592 369209 508626 369243
rect 508682 369209 508716 369243
rect 508772 369209 508806 369243
rect 508862 369209 508896 369243
rect 508952 369209 508986 369243
rect 509042 369209 509076 369243
rect 509132 369209 509166 369243
rect 509222 369209 509256 369243
rect 509312 369209 509346 369243
rect 509402 369209 509436 369243
rect 509492 369209 509526 369243
rect 509582 369209 509616 369243
rect 508502 369056 508536 369090
rect 508592 369056 508626 369090
rect 508682 369056 508716 369090
rect 508772 369056 508806 369090
rect 508862 369056 508896 369090
rect 508952 369056 508986 369090
rect 509042 369056 509076 369090
rect 509132 369056 509166 369090
rect 509222 369056 509256 369090
rect 509312 369056 509346 369090
rect 509402 369056 509436 369090
rect 509492 369056 509526 369090
rect 509582 369056 509616 369090
rect 508479 368960 508513 368994
rect 508479 368870 508513 368904
rect 508479 368780 508513 368814
rect 508479 368690 508513 368724
rect 508479 368600 508513 368634
rect 508479 368510 508513 368544
rect 508479 368420 508513 368454
rect 508479 368330 508513 368364
rect 508479 368240 508513 368274
rect 508479 368150 508513 368184
rect 508479 368060 508513 368094
rect 508479 367970 508513 368004
rect 509666 368960 509700 368994
rect 509666 368870 509700 368904
rect 509666 368780 509700 368814
rect 509666 368690 509700 368724
rect 509666 368600 509700 368634
rect 509666 368510 509700 368544
rect 509666 368420 509700 368454
rect 509666 368330 509700 368364
rect 509666 368240 509700 368274
rect 509666 368150 509700 368184
rect 509666 368060 509700 368094
rect 509666 367970 509700 368004
rect 508502 367869 508536 367903
rect 508592 367869 508626 367903
rect 508682 367869 508716 367903
rect 508772 367869 508806 367903
rect 508862 367869 508896 367903
rect 508952 367869 508986 367903
rect 509042 367869 509076 367903
rect 509132 367869 509166 367903
rect 509222 367869 509256 367903
rect 509312 367869 509346 367903
rect 509402 367869 509436 367903
rect 509492 367869 509526 367903
rect 509582 367869 509616 367903
rect 508502 367716 508536 367750
rect 508592 367716 508626 367750
rect 508682 367716 508716 367750
rect 508772 367716 508806 367750
rect 508862 367716 508896 367750
rect 508952 367716 508986 367750
rect 509042 367716 509076 367750
rect 509132 367716 509166 367750
rect 509222 367716 509256 367750
rect 509312 367716 509346 367750
rect 509402 367716 509436 367750
rect 509492 367716 509526 367750
rect 509582 367716 509616 367750
rect 508479 367620 508513 367654
rect 508479 367530 508513 367564
rect 508479 367440 508513 367474
rect 508479 367350 508513 367384
rect 508479 367260 508513 367294
rect 508479 367170 508513 367204
rect 508479 367080 508513 367114
rect 508479 366990 508513 367024
rect 508479 366900 508513 366934
rect 508479 366810 508513 366844
rect 508479 366720 508513 366754
rect 508479 366630 508513 366664
rect 509666 367620 509700 367654
rect 509666 367530 509700 367564
rect 509666 367440 509700 367474
rect 509666 367350 509700 367384
rect 509666 367260 509700 367294
rect 509666 367170 509700 367204
rect 509666 367080 509700 367114
rect 509666 366990 509700 367024
rect 509666 366900 509700 366934
rect 509666 366810 509700 366844
rect 509666 366720 509700 366754
rect 509666 366630 509700 366664
rect 508502 366529 508536 366563
rect 508592 366529 508626 366563
rect 508682 366529 508716 366563
rect 508772 366529 508806 366563
rect 508862 366529 508896 366563
rect 508952 366529 508986 366563
rect 509042 366529 509076 366563
rect 509132 366529 509166 366563
rect 509222 366529 509256 366563
rect 509312 366529 509346 366563
rect 509402 366529 509436 366563
rect 509492 366529 509526 366563
rect 509582 366529 509616 366563
rect 508502 366376 508536 366410
rect 508592 366376 508626 366410
rect 508682 366376 508716 366410
rect 508772 366376 508806 366410
rect 508862 366376 508896 366410
rect 508952 366376 508986 366410
rect 509042 366376 509076 366410
rect 509132 366376 509166 366410
rect 509222 366376 509256 366410
rect 509312 366376 509346 366410
rect 509402 366376 509436 366410
rect 509492 366376 509526 366410
rect 509582 366376 509616 366410
rect 508479 366280 508513 366314
rect 508479 366190 508513 366224
rect 508479 366100 508513 366134
rect 508479 366010 508513 366044
rect 508479 365920 508513 365954
rect 508479 365830 508513 365864
rect 508479 365740 508513 365774
rect 508479 365650 508513 365684
rect 508479 365560 508513 365594
rect 508479 365470 508513 365504
rect 508479 365380 508513 365414
rect 508479 365290 508513 365324
rect 509666 366280 509700 366314
rect 509666 366190 509700 366224
rect 509666 366100 509700 366134
rect 509666 366010 509700 366044
rect 509666 365920 509700 365954
rect 509666 365830 509700 365864
rect 509666 365740 509700 365774
rect 509666 365650 509700 365684
rect 509666 365560 509700 365594
rect 509666 365470 509700 365504
rect 509666 365380 509700 365414
rect 509666 365290 509700 365324
rect 508502 365189 508536 365223
rect 508592 365189 508626 365223
rect 508682 365189 508716 365223
rect 508772 365189 508806 365223
rect 508862 365189 508896 365223
rect 508952 365189 508986 365223
rect 509042 365189 509076 365223
rect 509132 365189 509166 365223
rect 509222 365189 509256 365223
rect 509312 365189 509346 365223
rect 509402 365189 509436 365223
rect 509492 365189 509526 365223
rect 509582 365189 509616 365223
rect 508502 365036 508536 365070
rect 508592 365036 508626 365070
rect 508682 365036 508716 365070
rect 508772 365036 508806 365070
rect 508862 365036 508896 365070
rect 508952 365036 508986 365070
rect 509042 365036 509076 365070
rect 509132 365036 509166 365070
rect 509222 365036 509256 365070
rect 509312 365036 509346 365070
rect 509402 365036 509436 365070
rect 509492 365036 509526 365070
rect 509582 365036 509616 365070
rect 508479 364940 508513 364974
rect 508479 364850 508513 364884
rect 508479 364760 508513 364794
rect 508479 364670 508513 364704
rect 508479 364580 508513 364614
rect 508479 364490 508513 364524
rect 508479 364400 508513 364434
rect 508479 364310 508513 364344
rect 508479 364220 508513 364254
rect 508479 364130 508513 364164
rect 508479 364040 508513 364074
rect 508479 363950 508513 363984
rect 509666 364940 509700 364974
rect 509666 364850 509700 364884
rect 509666 364760 509700 364794
rect 509666 364670 509700 364704
rect 509666 364580 509700 364614
rect 509666 364490 509700 364524
rect 509666 364400 509700 364434
rect 509666 364310 509700 364344
rect 509666 364220 509700 364254
rect 509666 364130 509700 364164
rect 509666 364040 509700 364074
rect 509666 363950 509700 363984
rect 508502 363849 508536 363883
rect 508592 363849 508626 363883
rect 508682 363849 508716 363883
rect 508772 363849 508806 363883
rect 508862 363849 508896 363883
rect 508952 363849 508986 363883
rect 509042 363849 509076 363883
rect 509132 363849 509166 363883
rect 509222 363849 509256 363883
rect 509312 363849 509346 363883
rect 509402 363849 509436 363883
rect 509492 363849 509526 363883
rect 509582 363849 509616 363883
rect 508502 363696 508536 363730
rect 508592 363696 508626 363730
rect 508682 363696 508716 363730
rect 508772 363696 508806 363730
rect 508862 363696 508896 363730
rect 508952 363696 508986 363730
rect 509042 363696 509076 363730
rect 509132 363696 509166 363730
rect 509222 363696 509256 363730
rect 509312 363696 509346 363730
rect 509402 363696 509436 363730
rect 509492 363696 509526 363730
rect 509582 363696 509616 363730
rect 508479 363600 508513 363634
rect 508479 363510 508513 363544
rect 508479 363420 508513 363454
rect 508479 363330 508513 363364
rect 508479 363240 508513 363274
rect 508479 363150 508513 363184
rect 508479 363060 508513 363094
rect 508479 362970 508513 363004
rect 508479 362880 508513 362914
rect 508479 362790 508513 362824
rect 508479 362700 508513 362734
rect 508479 362610 508513 362644
rect 509666 363600 509700 363634
rect 509666 363510 509700 363544
rect 509666 363420 509700 363454
rect 509666 363330 509700 363364
rect 509666 363240 509700 363274
rect 509666 363150 509700 363184
rect 509666 363060 509700 363094
rect 509666 362970 509700 363004
rect 509666 362880 509700 362914
rect 509666 362790 509700 362824
rect 509666 362700 509700 362734
rect 509666 362610 509700 362644
rect 508502 362509 508536 362543
rect 508592 362509 508626 362543
rect 508682 362509 508716 362543
rect 508772 362509 508806 362543
rect 508862 362509 508896 362543
rect 508952 362509 508986 362543
rect 509042 362509 509076 362543
rect 509132 362509 509166 362543
rect 509222 362509 509256 362543
rect 509312 362509 509346 362543
rect 509402 362509 509436 362543
rect 509492 362509 509526 362543
rect 509582 362509 509616 362543
rect 512262 373076 512296 373110
rect 512352 373076 512386 373110
rect 512442 373076 512476 373110
rect 512532 373076 512566 373110
rect 512622 373076 512656 373110
rect 512712 373076 512746 373110
rect 512802 373076 512836 373110
rect 512892 373076 512926 373110
rect 512982 373076 513016 373110
rect 513072 373076 513106 373110
rect 513162 373076 513196 373110
rect 513252 373076 513286 373110
rect 513342 373076 513376 373110
rect 512239 372980 512273 373014
rect 512239 372890 512273 372924
rect 512239 372800 512273 372834
rect 512239 372710 512273 372744
rect 512239 372620 512273 372654
rect 512239 372530 512273 372564
rect 512239 372440 512273 372474
rect 512239 372350 512273 372384
rect 512239 372260 512273 372294
rect 512239 372170 512273 372204
rect 512239 372080 512273 372114
rect 512239 371990 512273 372024
rect 513426 372980 513460 373014
rect 513426 372890 513460 372924
rect 513426 372800 513460 372834
rect 513426 372710 513460 372744
rect 513426 372620 513460 372654
rect 513426 372530 513460 372564
rect 513426 372440 513460 372474
rect 513426 372350 513460 372384
rect 516617 373375 516719 373817
rect 520377 373375 520479 373817
rect 513426 372260 513460 372294
rect 513426 372170 513460 372204
rect 513426 372080 513460 372114
rect 513426 371990 513460 372024
rect 512262 371889 512296 371923
rect 512352 371889 512386 371923
rect 512442 371889 512476 371923
rect 512532 371889 512566 371923
rect 512622 371889 512656 371923
rect 512712 371889 512746 371923
rect 512802 371889 512836 371923
rect 512892 371889 512926 371923
rect 512982 371889 513016 371923
rect 513072 371889 513106 371923
rect 513162 371889 513196 371923
rect 513252 371889 513286 371923
rect 513342 371889 513376 371923
rect 512262 371736 512296 371770
rect 512352 371736 512386 371770
rect 512442 371736 512476 371770
rect 512532 371736 512566 371770
rect 512622 371736 512656 371770
rect 512712 371736 512746 371770
rect 512802 371736 512836 371770
rect 512892 371736 512926 371770
rect 512982 371736 513016 371770
rect 513072 371736 513106 371770
rect 513162 371736 513196 371770
rect 513252 371736 513286 371770
rect 513342 371736 513376 371770
rect 512239 371640 512273 371674
rect 512239 371550 512273 371584
rect 512239 371460 512273 371494
rect 512239 371370 512273 371404
rect 512239 371280 512273 371314
rect 512239 371190 512273 371224
rect 512239 371100 512273 371134
rect 512239 371010 512273 371044
rect 512239 370920 512273 370954
rect 512239 370830 512273 370864
rect 512239 370740 512273 370774
rect 512239 370650 512273 370684
rect 513426 371640 513460 371674
rect 513426 371550 513460 371584
rect 513426 371460 513460 371494
rect 513426 371370 513460 371404
rect 513426 371280 513460 371314
rect 513426 371190 513460 371224
rect 513426 371100 513460 371134
rect 513426 371010 513460 371044
rect 513426 370920 513460 370954
rect 513426 370830 513460 370864
rect 513426 370740 513460 370774
rect 513426 370650 513460 370684
rect 512262 370549 512296 370583
rect 512352 370549 512386 370583
rect 512442 370549 512476 370583
rect 512532 370549 512566 370583
rect 512622 370549 512656 370583
rect 512712 370549 512746 370583
rect 512802 370549 512836 370583
rect 512892 370549 512926 370583
rect 512982 370549 513016 370583
rect 513072 370549 513106 370583
rect 513162 370549 513196 370583
rect 513252 370549 513286 370583
rect 513342 370549 513376 370583
rect 512262 370396 512296 370430
rect 512352 370396 512386 370430
rect 512442 370396 512476 370430
rect 512532 370396 512566 370430
rect 512622 370396 512656 370430
rect 512712 370396 512746 370430
rect 512802 370396 512836 370430
rect 512892 370396 512926 370430
rect 512982 370396 513016 370430
rect 513072 370396 513106 370430
rect 513162 370396 513196 370430
rect 513252 370396 513286 370430
rect 513342 370396 513376 370430
rect 512239 370300 512273 370334
rect 512239 370210 512273 370244
rect 512239 370120 512273 370154
rect 512239 370030 512273 370064
rect 512239 369940 512273 369974
rect 512239 369850 512273 369884
rect 512239 369760 512273 369794
rect 512239 369670 512273 369704
rect 512239 369580 512273 369614
rect 512239 369490 512273 369524
rect 512239 369400 512273 369434
rect 512239 369310 512273 369344
rect 513426 370300 513460 370334
rect 513426 370210 513460 370244
rect 513426 370120 513460 370154
rect 513426 370030 513460 370064
rect 513426 369940 513460 369974
rect 513426 369850 513460 369884
rect 513426 369760 513460 369794
rect 513426 369670 513460 369704
rect 516617 370631 516719 371073
rect 513426 369580 513460 369614
rect 513426 369490 513460 369524
rect 513426 369400 513460 369434
rect 513426 369310 513460 369344
rect 512262 369209 512296 369243
rect 512352 369209 512386 369243
rect 512442 369209 512476 369243
rect 512532 369209 512566 369243
rect 512622 369209 512656 369243
rect 512712 369209 512746 369243
rect 512802 369209 512836 369243
rect 512892 369209 512926 369243
rect 512982 369209 513016 369243
rect 513072 369209 513106 369243
rect 513162 369209 513196 369243
rect 513252 369209 513286 369243
rect 513342 369209 513376 369243
rect 512262 369056 512296 369090
rect 512352 369056 512386 369090
rect 512442 369056 512476 369090
rect 512532 369056 512566 369090
rect 512622 369056 512656 369090
rect 512712 369056 512746 369090
rect 512802 369056 512836 369090
rect 512892 369056 512926 369090
rect 512982 369056 513016 369090
rect 513072 369056 513106 369090
rect 513162 369056 513196 369090
rect 513252 369056 513286 369090
rect 513342 369056 513376 369090
rect 512239 368960 512273 368994
rect 512239 368870 512273 368904
rect 512239 368780 512273 368814
rect 512239 368690 512273 368724
rect 512239 368600 512273 368634
rect 512239 368510 512273 368544
rect 512239 368420 512273 368454
rect 512239 368330 512273 368364
rect 512239 368240 512273 368274
rect 512239 368150 512273 368184
rect 512239 368060 512273 368094
rect 512239 367970 512273 368004
rect 513426 368960 513460 368994
rect 513426 368870 513460 368904
rect 513426 368780 513460 368814
rect 513426 368690 513460 368724
rect 513426 368600 513460 368634
rect 513426 368510 513460 368544
rect 513426 368420 513460 368454
rect 513426 368330 513460 368364
rect 513426 368240 513460 368274
rect 513426 368150 513460 368184
rect 513426 368060 513460 368094
rect 513426 367970 513460 368004
rect 512262 367869 512296 367903
rect 512352 367869 512386 367903
rect 512442 367869 512476 367903
rect 512532 367869 512566 367903
rect 512622 367869 512656 367903
rect 512712 367869 512746 367903
rect 512802 367869 512836 367903
rect 512892 367869 512926 367903
rect 512982 367869 513016 367903
rect 513072 367869 513106 367903
rect 513162 367869 513196 367903
rect 513252 367869 513286 367903
rect 513342 367869 513376 367903
rect 512262 367716 512296 367750
rect 512352 367716 512386 367750
rect 512442 367716 512476 367750
rect 512532 367716 512566 367750
rect 512622 367716 512656 367750
rect 512712 367716 512746 367750
rect 512802 367716 512836 367750
rect 512892 367716 512926 367750
rect 512982 367716 513016 367750
rect 513072 367716 513106 367750
rect 513162 367716 513196 367750
rect 513252 367716 513286 367750
rect 513342 367716 513376 367750
rect 512239 367620 512273 367654
rect 512239 367530 512273 367564
rect 512239 367440 512273 367474
rect 512239 367350 512273 367384
rect 512239 367260 512273 367294
rect 512239 367170 512273 367204
rect 512239 367080 512273 367114
rect 512239 366990 512273 367024
rect 512239 366900 512273 366934
rect 512239 366810 512273 366844
rect 512239 366720 512273 366754
rect 512239 366630 512273 366664
rect 513426 367620 513460 367654
rect 513426 367530 513460 367564
rect 513426 367440 513460 367474
rect 513426 367350 513460 367384
rect 513426 367260 513460 367294
rect 513426 367170 513460 367204
rect 513426 367080 513460 367114
rect 513426 366990 513460 367024
rect 513426 366900 513460 366934
rect 516617 367887 516719 368329
rect 527897 369651 527999 370093
rect 531657 369749 531759 370191
rect 513426 366810 513460 366844
rect 513426 366720 513460 366754
rect 513426 366630 513460 366664
rect 512262 366529 512296 366563
rect 512352 366529 512386 366563
rect 512442 366529 512476 366563
rect 512532 366529 512566 366563
rect 512622 366529 512656 366563
rect 512712 366529 512746 366563
rect 512802 366529 512836 366563
rect 512892 366529 512926 366563
rect 512982 366529 513016 366563
rect 513072 366529 513106 366563
rect 513162 366529 513196 366563
rect 513252 366529 513286 366563
rect 513342 366529 513376 366563
rect 512262 366376 512296 366410
rect 512352 366376 512386 366410
rect 512442 366376 512476 366410
rect 512532 366376 512566 366410
rect 512622 366376 512656 366410
rect 512712 366376 512746 366410
rect 512802 366376 512836 366410
rect 512892 366376 512926 366410
rect 512982 366376 513016 366410
rect 513072 366376 513106 366410
rect 513162 366376 513196 366410
rect 513252 366376 513286 366410
rect 513342 366376 513376 366410
rect 512239 366280 512273 366314
rect 512239 366190 512273 366224
rect 512239 366100 512273 366134
rect 512239 366010 512273 366044
rect 512239 365920 512273 365954
rect 512239 365830 512273 365864
rect 512239 365740 512273 365774
rect 512239 365650 512273 365684
rect 512239 365560 512273 365594
rect 512239 365470 512273 365504
rect 512239 365380 512273 365414
rect 512239 365290 512273 365324
rect 513426 366280 513460 366314
rect 513426 366190 513460 366224
rect 513426 366100 513460 366134
rect 513426 366010 513460 366044
rect 513426 365920 513460 365954
rect 513426 365830 513460 365864
rect 513426 365740 513460 365774
rect 513426 365650 513460 365684
rect 513426 365560 513460 365594
rect 513426 365470 513460 365504
rect 513426 365380 513460 365414
rect 513426 365290 513460 365324
rect 512262 365189 512296 365223
rect 512352 365189 512386 365223
rect 512442 365189 512476 365223
rect 512532 365189 512566 365223
rect 512622 365189 512656 365223
rect 512712 365189 512746 365223
rect 512802 365189 512836 365223
rect 512892 365189 512926 365223
rect 512982 365189 513016 365223
rect 513072 365189 513106 365223
rect 513162 365189 513196 365223
rect 513252 365189 513286 365223
rect 513342 365189 513376 365223
rect 512262 365036 512296 365070
rect 512352 365036 512386 365070
rect 512442 365036 512476 365070
rect 512532 365036 512566 365070
rect 512622 365036 512656 365070
rect 512712 365036 512746 365070
rect 512802 365036 512836 365070
rect 512892 365036 512926 365070
rect 512982 365036 513016 365070
rect 513072 365036 513106 365070
rect 513162 365036 513196 365070
rect 513252 365036 513286 365070
rect 513342 365036 513376 365070
rect 512239 364940 512273 364974
rect 512239 364850 512273 364884
rect 512239 364760 512273 364794
rect 512239 364670 512273 364704
rect 512239 364580 512273 364614
rect 512239 364490 512273 364524
rect 512239 364400 512273 364434
rect 512239 364310 512273 364344
rect 512239 364220 512273 364254
rect 512239 364130 512273 364164
rect 512239 364040 512273 364074
rect 512239 363950 512273 363984
rect 513426 364940 513460 364974
rect 513426 364850 513460 364884
rect 513426 364760 513460 364794
rect 513426 364670 513460 364704
rect 513426 364580 513460 364614
rect 513426 364490 513460 364524
rect 513426 364400 513460 364434
rect 513426 364310 513460 364344
rect 513426 364220 513460 364254
rect 513426 364130 513460 364164
rect 516617 365143 516719 365585
rect 520377 365143 520479 365585
rect 527897 366907 527999 367349
rect 531657 367005 531759 367447
rect 535417 368965 535519 369407
rect 513426 364040 513460 364074
rect 513426 363950 513460 363984
rect 512262 363849 512296 363883
rect 512352 363849 512386 363883
rect 512442 363849 512476 363883
rect 512532 363849 512566 363883
rect 512622 363849 512656 363883
rect 512712 363849 512746 363883
rect 512802 363849 512836 363883
rect 512892 363849 512926 363883
rect 512982 363849 513016 363883
rect 513072 363849 513106 363883
rect 513162 363849 513196 363883
rect 513252 363849 513286 363883
rect 513342 363849 513376 363883
rect 512262 363696 512296 363730
rect 512352 363696 512386 363730
rect 512442 363696 512476 363730
rect 512532 363696 512566 363730
rect 512622 363696 512656 363730
rect 512712 363696 512746 363730
rect 512802 363696 512836 363730
rect 512892 363696 512926 363730
rect 512982 363696 513016 363730
rect 513072 363696 513106 363730
rect 513162 363696 513196 363730
rect 513252 363696 513286 363730
rect 513342 363696 513376 363730
rect 512239 363600 512273 363634
rect 512239 363510 512273 363544
rect 512239 363420 512273 363454
rect 512239 363330 512273 363364
rect 512239 363240 512273 363274
rect 512239 363150 512273 363184
rect 512239 363060 512273 363094
rect 512239 362970 512273 363004
rect 512239 362880 512273 362914
rect 512239 362790 512273 362824
rect 512239 362700 512273 362734
rect 512239 362610 512273 362644
rect 513426 363600 513460 363634
rect 513426 363510 513460 363544
rect 513426 363420 513460 363454
rect 513426 363330 513460 363364
rect 513426 363240 513460 363274
rect 513426 363150 513460 363184
rect 513426 363060 513460 363094
rect 527897 364163 527999 364605
rect 531657 364261 531759 364703
rect 535417 366221 535519 366663
rect 513426 362970 513460 363004
rect 513426 362880 513460 362914
rect 513426 362790 513460 362824
rect 513426 362700 513460 362734
rect 513426 362610 513460 362644
rect 512262 362509 512296 362543
rect 512352 362509 512386 362543
rect 512442 362509 512476 362543
rect 512532 362509 512566 362543
rect 512622 362509 512656 362543
rect 512712 362509 512746 362543
rect 512802 362509 512836 362543
rect 512892 362509 512926 362543
rect 512982 362509 513016 362543
rect 513072 362509 513106 362543
rect 513162 362509 513196 362543
rect 513252 362509 513286 362543
rect 513342 362509 513376 362543
rect 535417 363477 535519 363919
rect 562076 357572 562120 357608
rect 563376 357572 563420 357608
rect 564676 357572 564720 357608
rect 565778 357600 565818 357640
rect 561938 311264 561982 311300
rect 563238 311264 563282 311300
rect 564538 311264 564582 311300
rect 565640 311292 565680 311332
<< nsubdiffcont >>
rect 576776 493486 576820 493522
rect 578076 493486 578120 493522
rect 579376 493486 579420 493522
rect 580478 493434 580518 493474
rect 576054 404610 576098 404646
rect 577354 404610 577398 404646
rect 578654 404610 578698 404646
rect 579756 404558 579796 404598
rect 504923 402720 504957 402754
rect 505013 402720 505047 402754
rect 505103 402720 505137 402754
rect 505193 402720 505227 402754
rect 505283 402720 505317 402754
rect 505373 402720 505407 402754
rect 505463 402720 505497 402754
rect 505553 402720 505587 402754
rect 505643 402720 505677 402754
rect 504866 402608 504900 402642
rect 505756 402642 505790 402676
rect 504866 402518 504900 402552
rect 504866 402428 504900 402462
rect 504866 402338 504900 402372
rect 504866 402248 504900 402282
rect 504866 402158 504900 402192
rect 504866 402068 504900 402102
rect 504866 401978 504900 402012
rect 505756 402552 505790 402586
rect 505756 402462 505790 402496
rect 505756 402372 505790 402406
rect 505756 402282 505790 402316
rect 505756 402192 505790 402226
rect 505756 402102 505790 402136
rect 505756 402012 505790 402046
rect 504866 401888 504900 401922
rect 505756 401922 505790 401956
rect 504942 401830 504976 401864
rect 505032 401830 505066 401864
rect 505122 401830 505156 401864
rect 505212 401830 505246 401864
rect 505302 401830 505336 401864
rect 505392 401830 505426 401864
rect 505482 401830 505516 401864
rect 505572 401830 505606 401864
rect 505662 401830 505696 401864
rect 496991 399947 497025 399981
rect 496941 398847 496975 398881
rect 496941 397547 496975 397581
rect 496941 396247 496975 396281
rect 496941 394947 496975 394981
rect 496941 393647 496975 393681
rect 496941 392347 496975 392381
rect 500751 392303 500785 392337
rect 496941 391047 496975 391081
rect 500701 391203 500735 391237
rect 493231 390147 493265 390181
rect 496941 389747 496975 389781
rect 500701 389903 500735 389937
rect 493181 389047 493215 389081
rect 496941 388447 496975 388481
rect 500701 388603 500735 388637
rect 493181 387747 493215 387781
rect 523311 390147 523345 390181
rect 523261 389047 523295 389081
rect 496941 387147 496975 387181
rect 493181 386447 493215 386481
rect 496941 385847 496975 385881
rect 493181 385147 493215 385181
rect 500751 385639 500785 385673
rect 523261 387747 523295 387781
rect 523261 386447 523295 386481
rect 496941 384547 496975 384581
rect 523261 385147 523295 385181
rect 493181 383847 493215 383881
rect 500701 384539 500735 384573
rect 496941 383247 496975 383281
rect 500701 383239 500735 383273
rect 493181 382547 493215 382581
rect 523261 383847 523295 383881
rect 496941 381947 496975 381981
rect 500701 381939 500735 381973
rect 523261 382547 523295 382581
rect 493181 381247 493215 381281
rect 496941 380647 496975 380681
rect 493181 379947 493215 379981
rect 496941 379347 496975 379381
rect 523261 381247 523295 381281
rect 523261 379947 523295 379981
rect 493181 378647 493215 378681
rect 523261 378647 523295 378681
rect 496941 378047 496975 378081
rect 493181 377347 493215 377381
rect 504511 377505 504545 377539
rect 512031 377505 512065 377539
rect 496941 376747 496975 376781
rect 493181 376047 493215 376081
rect 504461 376405 504495 376439
rect 511981 376405 512015 376439
rect 496941 375447 496975 375481
rect 493181 374747 493215 374781
rect 496941 374147 496975 374181
rect 493181 373447 493215 373481
rect 523261 377347 523295 377381
rect 523261 376047 523295 376081
rect 493181 372147 493215 372181
rect 501163 372928 501197 372962
rect 501253 372928 501287 372962
rect 501343 372928 501377 372962
rect 501433 372928 501467 372962
rect 501523 372928 501557 372962
rect 501613 372928 501647 372962
rect 501703 372928 501737 372962
rect 501793 372928 501827 372962
rect 501883 372928 501917 372962
rect 501106 372816 501140 372850
rect 501996 372850 502030 372884
rect 501106 372726 501140 372760
rect 501106 372636 501140 372670
rect 501106 372546 501140 372580
rect 501106 372456 501140 372490
rect 501106 372366 501140 372400
rect 501106 372276 501140 372310
rect 501106 372186 501140 372220
rect 501996 372760 502030 372794
rect 501996 372670 502030 372704
rect 501996 372580 502030 372614
rect 501996 372490 502030 372524
rect 501996 372400 502030 372434
rect 501996 372310 502030 372344
rect 501996 372220 502030 372254
rect 501106 372096 501140 372130
rect 501996 372130 502030 372164
rect 501182 372038 501216 372072
rect 501272 372038 501306 372072
rect 501362 372038 501396 372072
rect 501452 372038 501486 372072
rect 501542 372038 501576 372072
rect 501632 372038 501666 372072
rect 501722 372038 501756 372072
rect 501812 372038 501846 372072
rect 501902 372038 501936 372072
rect 493181 370847 493215 370881
rect 493181 369547 493215 369581
rect 493181 368247 493215 368281
rect 493181 366947 493215 366981
rect 493181 365647 493215 365681
rect 493181 364347 493215 364381
rect 497403 371752 497437 371786
rect 497493 371752 497527 371786
rect 497583 371752 497617 371786
rect 497673 371752 497707 371786
rect 497763 371752 497797 371786
rect 497853 371752 497887 371786
rect 497943 371752 497977 371786
rect 498033 371752 498067 371786
rect 498123 371752 498157 371786
rect 497346 371640 497380 371674
rect 498236 371674 498270 371708
rect 497346 371550 497380 371584
rect 497346 371460 497380 371494
rect 497346 371370 497380 371404
rect 497346 371280 497380 371314
rect 497346 371190 497380 371224
rect 497346 371100 497380 371134
rect 497346 371010 497380 371044
rect 498236 371584 498270 371618
rect 498236 371494 498270 371528
rect 498236 371404 498270 371438
rect 498236 371314 498270 371348
rect 498236 371224 498270 371258
rect 498236 371134 498270 371168
rect 498236 371044 498270 371078
rect 497346 370920 497380 370954
rect 498236 370954 498270 370988
rect 497422 370862 497456 370896
rect 497512 370862 497546 370896
rect 497602 370862 497636 370896
rect 497692 370862 497726 370896
rect 497782 370862 497816 370896
rect 497872 370862 497906 370896
rect 497962 370862 497996 370896
rect 498052 370862 498086 370896
rect 498142 370862 498176 370896
rect 497403 370412 497437 370446
rect 497493 370412 497527 370446
rect 497583 370412 497617 370446
rect 497673 370412 497707 370446
rect 497763 370412 497797 370446
rect 497853 370412 497887 370446
rect 497943 370412 497977 370446
rect 498033 370412 498067 370446
rect 498123 370412 498157 370446
rect 497346 370300 497380 370334
rect 498236 370334 498270 370368
rect 497346 370210 497380 370244
rect 497346 370120 497380 370154
rect 497346 370030 497380 370064
rect 497346 369940 497380 369974
rect 497346 369850 497380 369884
rect 497346 369760 497380 369794
rect 497346 369670 497380 369704
rect 498236 370244 498270 370278
rect 498236 370154 498270 370188
rect 498236 370064 498270 370098
rect 498236 369974 498270 370008
rect 498236 369884 498270 369918
rect 498236 369794 498270 369828
rect 498236 369704 498270 369738
rect 497346 369580 497380 369614
rect 498236 369614 498270 369648
rect 497422 369522 497456 369556
rect 497512 369522 497546 369556
rect 497602 369522 497636 369556
rect 497692 369522 497726 369556
rect 497782 369522 497816 369556
rect 497872 369522 497906 369556
rect 497962 369522 497996 369556
rect 498052 369522 498086 369556
rect 498142 369522 498176 369556
rect 497403 369072 497437 369106
rect 497493 369072 497527 369106
rect 497583 369072 497617 369106
rect 497673 369072 497707 369106
rect 497763 369072 497797 369106
rect 497853 369072 497887 369106
rect 497943 369072 497977 369106
rect 498033 369072 498067 369106
rect 498123 369072 498157 369106
rect 497346 368960 497380 368994
rect 498236 368994 498270 369028
rect 497346 368870 497380 368904
rect 497346 368780 497380 368814
rect 497346 368690 497380 368724
rect 497346 368600 497380 368634
rect 497346 368510 497380 368544
rect 497346 368420 497380 368454
rect 497346 368330 497380 368364
rect 498236 368904 498270 368938
rect 498236 368814 498270 368848
rect 498236 368724 498270 368758
rect 498236 368634 498270 368668
rect 498236 368544 498270 368578
rect 498236 368454 498270 368488
rect 498236 368364 498270 368398
rect 497346 368240 497380 368274
rect 498236 368274 498270 368308
rect 497422 368182 497456 368216
rect 497512 368182 497546 368216
rect 497602 368182 497636 368216
rect 497692 368182 497726 368216
rect 497782 368182 497816 368216
rect 497872 368182 497906 368216
rect 497962 368182 497996 368216
rect 498052 368182 498086 368216
rect 498142 368182 498176 368216
rect 497403 367732 497437 367766
rect 497493 367732 497527 367766
rect 497583 367732 497617 367766
rect 497673 367732 497707 367766
rect 497763 367732 497797 367766
rect 497853 367732 497887 367766
rect 497943 367732 497977 367766
rect 498033 367732 498067 367766
rect 498123 367732 498157 367766
rect 497346 367620 497380 367654
rect 498236 367654 498270 367688
rect 497346 367530 497380 367564
rect 497346 367440 497380 367474
rect 497346 367350 497380 367384
rect 497346 367260 497380 367294
rect 497346 367170 497380 367204
rect 497346 367080 497380 367114
rect 497346 366990 497380 367024
rect 498236 367564 498270 367598
rect 498236 367474 498270 367508
rect 498236 367384 498270 367418
rect 498236 367294 498270 367328
rect 498236 367204 498270 367238
rect 498236 367114 498270 367148
rect 498236 367024 498270 367058
rect 497346 366900 497380 366934
rect 498236 366934 498270 366968
rect 497422 366842 497456 366876
rect 497512 366842 497546 366876
rect 497602 366842 497636 366876
rect 497692 366842 497726 366876
rect 497782 366842 497816 366876
rect 497872 366842 497906 366876
rect 497962 366842 497996 366876
rect 498052 366842 498086 366876
rect 498142 366842 498176 366876
rect 497403 366392 497437 366426
rect 497493 366392 497527 366426
rect 497583 366392 497617 366426
rect 497673 366392 497707 366426
rect 497763 366392 497797 366426
rect 497853 366392 497887 366426
rect 497943 366392 497977 366426
rect 498033 366392 498067 366426
rect 498123 366392 498157 366426
rect 497346 366280 497380 366314
rect 498236 366314 498270 366348
rect 497346 366190 497380 366224
rect 497346 366100 497380 366134
rect 497346 366010 497380 366044
rect 497346 365920 497380 365954
rect 497346 365830 497380 365864
rect 497346 365740 497380 365774
rect 497346 365650 497380 365684
rect 498236 366224 498270 366258
rect 498236 366134 498270 366168
rect 498236 366044 498270 366078
rect 498236 365954 498270 365988
rect 498236 365864 498270 365898
rect 498236 365774 498270 365808
rect 498236 365684 498270 365718
rect 497346 365560 497380 365594
rect 498236 365594 498270 365628
rect 497422 365502 497456 365536
rect 497512 365502 497546 365536
rect 497602 365502 497636 365536
rect 497692 365502 497726 365536
rect 497782 365502 497816 365536
rect 497872 365502 497906 365536
rect 497962 365502 497996 365536
rect 498052 365502 498086 365536
rect 498142 365502 498176 365536
rect 497403 365052 497437 365086
rect 497493 365052 497527 365086
rect 497583 365052 497617 365086
rect 497673 365052 497707 365086
rect 497763 365052 497797 365086
rect 497853 365052 497887 365086
rect 497943 365052 497977 365086
rect 498033 365052 498067 365086
rect 498123 365052 498157 365086
rect 497346 364940 497380 364974
rect 498236 364974 498270 365008
rect 497346 364850 497380 364884
rect 497346 364760 497380 364794
rect 497346 364670 497380 364704
rect 497346 364580 497380 364614
rect 497346 364490 497380 364524
rect 497346 364400 497380 364434
rect 497346 364310 497380 364344
rect 498236 364884 498270 364918
rect 498236 364794 498270 364828
rect 498236 364704 498270 364738
rect 498236 364614 498270 364648
rect 498236 364524 498270 364558
rect 498236 364434 498270 364468
rect 498236 364344 498270 364378
rect 497346 364220 497380 364254
rect 498236 364254 498270 364288
rect 497422 364162 497456 364196
rect 497512 364162 497546 364196
rect 497602 364162 497636 364196
rect 497692 364162 497726 364196
rect 497782 364162 497816 364196
rect 497872 364162 497906 364196
rect 497962 364162 497996 364196
rect 498052 364162 498086 364196
rect 498142 364162 498176 364196
rect 497403 363712 497437 363746
rect 497493 363712 497527 363746
rect 497583 363712 497617 363746
rect 497673 363712 497707 363746
rect 497763 363712 497797 363746
rect 497853 363712 497887 363746
rect 497943 363712 497977 363746
rect 498033 363712 498067 363746
rect 498123 363712 498157 363746
rect 497346 363600 497380 363634
rect 498236 363634 498270 363668
rect 497346 363510 497380 363544
rect 497346 363420 497380 363454
rect 497346 363330 497380 363364
rect 497346 363240 497380 363274
rect 497346 363150 497380 363184
rect 497346 363060 497380 363094
rect 497346 362970 497380 363004
rect 498236 363544 498270 363578
rect 498236 363454 498270 363488
rect 498236 363364 498270 363398
rect 498236 363274 498270 363308
rect 498236 363184 498270 363218
rect 498236 363094 498270 363128
rect 498236 363004 498270 363038
rect 497346 362880 497380 362914
rect 498236 362914 498270 362948
rect 497422 362822 497456 362856
rect 497512 362822 497546 362856
rect 497602 362822 497636 362856
rect 497692 362822 497726 362856
rect 497782 362822 497816 362856
rect 497872 362822 497906 362856
rect 497962 362822 497996 362856
rect 498052 362822 498086 362856
rect 498142 362822 498176 362856
rect 501163 371588 501197 371622
rect 501253 371588 501287 371622
rect 501343 371588 501377 371622
rect 501433 371588 501467 371622
rect 501523 371588 501557 371622
rect 501613 371588 501647 371622
rect 501703 371588 501737 371622
rect 501793 371588 501827 371622
rect 501883 371588 501917 371622
rect 501106 371476 501140 371510
rect 501996 371510 502030 371544
rect 501106 371386 501140 371420
rect 501106 371296 501140 371330
rect 501106 371206 501140 371240
rect 501106 371116 501140 371150
rect 501106 371026 501140 371060
rect 501106 370936 501140 370970
rect 501106 370846 501140 370880
rect 501996 371420 502030 371454
rect 501996 371330 502030 371364
rect 501996 371240 502030 371274
rect 501996 371150 502030 371184
rect 501996 371060 502030 371094
rect 501996 370970 502030 371004
rect 501996 370880 502030 370914
rect 501106 370756 501140 370790
rect 501996 370790 502030 370824
rect 501182 370698 501216 370732
rect 501272 370698 501306 370732
rect 501362 370698 501396 370732
rect 501452 370698 501486 370732
rect 501542 370698 501576 370732
rect 501632 370698 501666 370732
rect 501722 370698 501756 370732
rect 501812 370698 501846 370732
rect 501902 370698 501936 370732
rect 501163 370248 501197 370282
rect 501253 370248 501287 370282
rect 501343 370248 501377 370282
rect 501433 370248 501467 370282
rect 501523 370248 501557 370282
rect 501613 370248 501647 370282
rect 501703 370248 501737 370282
rect 501793 370248 501827 370282
rect 501883 370248 501917 370282
rect 501106 370136 501140 370170
rect 501996 370170 502030 370204
rect 501106 370046 501140 370080
rect 501106 369956 501140 369990
rect 501106 369866 501140 369900
rect 501106 369776 501140 369810
rect 501106 369686 501140 369720
rect 501106 369596 501140 369630
rect 501106 369506 501140 369540
rect 501996 370080 502030 370114
rect 501996 369990 502030 370024
rect 501996 369900 502030 369934
rect 501996 369810 502030 369844
rect 501996 369720 502030 369754
rect 501996 369630 502030 369664
rect 501996 369540 502030 369574
rect 501106 369416 501140 369450
rect 501996 369450 502030 369484
rect 501182 369358 501216 369392
rect 501272 369358 501306 369392
rect 501362 369358 501396 369392
rect 501452 369358 501486 369392
rect 501542 369358 501576 369392
rect 501632 369358 501666 369392
rect 501722 369358 501756 369392
rect 501812 369358 501846 369392
rect 501902 369358 501936 369392
rect 501163 368908 501197 368942
rect 501253 368908 501287 368942
rect 501343 368908 501377 368942
rect 501433 368908 501467 368942
rect 501523 368908 501557 368942
rect 501613 368908 501647 368942
rect 501703 368908 501737 368942
rect 501793 368908 501827 368942
rect 501883 368908 501917 368942
rect 501106 368796 501140 368830
rect 501996 368830 502030 368864
rect 501106 368706 501140 368740
rect 501106 368616 501140 368650
rect 501106 368526 501140 368560
rect 501106 368436 501140 368470
rect 501106 368346 501140 368380
rect 501106 368256 501140 368290
rect 501106 368166 501140 368200
rect 501996 368740 502030 368774
rect 501996 368650 502030 368684
rect 501996 368560 502030 368594
rect 501996 368470 502030 368504
rect 501996 368380 502030 368414
rect 501996 368290 502030 368324
rect 501996 368200 502030 368234
rect 501106 368076 501140 368110
rect 501996 368110 502030 368144
rect 501182 368018 501216 368052
rect 501272 368018 501306 368052
rect 501362 368018 501396 368052
rect 501452 368018 501486 368052
rect 501542 368018 501576 368052
rect 501632 368018 501666 368052
rect 501722 368018 501756 368052
rect 501812 368018 501846 368052
rect 501902 368018 501936 368052
rect 501163 367568 501197 367602
rect 501253 367568 501287 367602
rect 501343 367568 501377 367602
rect 501433 367568 501467 367602
rect 501523 367568 501557 367602
rect 501613 367568 501647 367602
rect 501703 367568 501737 367602
rect 501793 367568 501827 367602
rect 501883 367568 501917 367602
rect 501106 367456 501140 367490
rect 501996 367490 502030 367524
rect 501106 367366 501140 367400
rect 501106 367276 501140 367310
rect 501106 367186 501140 367220
rect 501106 367096 501140 367130
rect 501106 367006 501140 367040
rect 501106 366916 501140 366950
rect 501106 366826 501140 366860
rect 501996 367400 502030 367434
rect 501996 367310 502030 367344
rect 501996 367220 502030 367254
rect 501996 367130 502030 367164
rect 501996 367040 502030 367074
rect 501996 366950 502030 366984
rect 501996 366860 502030 366894
rect 501106 366736 501140 366770
rect 501996 366770 502030 366804
rect 501182 366678 501216 366712
rect 501272 366678 501306 366712
rect 501362 366678 501396 366712
rect 501452 366678 501486 366712
rect 501542 366678 501576 366712
rect 501632 366678 501666 366712
rect 501722 366678 501756 366712
rect 501812 366678 501846 366712
rect 501902 366678 501936 366712
rect 501163 366228 501197 366262
rect 501253 366228 501287 366262
rect 501343 366228 501377 366262
rect 501433 366228 501467 366262
rect 501523 366228 501557 366262
rect 501613 366228 501647 366262
rect 501703 366228 501737 366262
rect 501793 366228 501827 366262
rect 501883 366228 501917 366262
rect 501106 366116 501140 366150
rect 501996 366150 502030 366184
rect 501106 366026 501140 366060
rect 501106 365936 501140 365970
rect 501106 365846 501140 365880
rect 501106 365756 501140 365790
rect 501106 365666 501140 365700
rect 501106 365576 501140 365610
rect 501106 365486 501140 365520
rect 501996 366060 502030 366094
rect 501996 365970 502030 366004
rect 501996 365880 502030 365914
rect 501996 365790 502030 365824
rect 501996 365700 502030 365734
rect 501996 365610 502030 365644
rect 501996 365520 502030 365554
rect 501106 365396 501140 365430
rect 501996 365430 502030 365464
rect 501182 365338 501216 365372
rect 501272 365338 501306 365372
rect 501362 365338 501396 365372
rect 501452 365338 501486 365372
rect 501542 365338 501576 365372
rect 501632 365338 501666 365372
rect 501722 365338 501756 365372
rect 501812 365338 501846 365372
rect 501902 365338 501936 365372
rect 501163 364888 501197 364922
rect 501253 364888 501287 364922
rect 501343 364888 501377 364922
rect 501433 364888 501467 364922
rect 501523 364888 501557 364922
rect 501613 364888 501647 364922
rect 501703 364888 501737 364922
rect 501793 364888 501827 364922
rect 501883 364888 501917 364922
rect 501106 364776 501140 364810
rect 501996 364810 502030 364844
rect 501106 364686 501140 364720
rect 501106 364596 501140 364630
rect 501106 364506 501140 364540
rect 501106 364416 501140 364450
rect 501106 364326 501140 364360
rect 501106 364236 501140 364270
rect 501106 364146 501140 364180
rect 501996 364720 502030 364754
rect 501996 364630 502030 364664
rect 501996 364540 502030 364574
rect 501996 364450 502030 364484
rect 501996 364360 502030 364394
rect 501996 364270 502030 364304
rect 501996 364180 502030 364214
rect 501106 364056 501140 364090
rect 501996 364090 502030 364124
rect 501182 363998 501216 364032
rect 501272 363998 501306 364032
rect 501362 363998 501396 364032
rect 501452 363998 501486 364032
rect 501542 363998 501576 364032
rect 501632 363998 501666 364032
rect 501722 363998 501756 364032
rect 501812 363998 501846 364032
rect 501902 363998 501936 364032
rect 501163 363548 501197 363582
rect 501253 363548 501287 363582
rect 501343 363548 501377 363582
rect 501433 363548 501467 363582
rect 501523 363548 501557 363582
rect 501613 363548 501647 363582
rect 501703 363548 501737 363582
rect 501793 363548 501827 363582
rect 501883 363548 501917 363582
rect 501106 363436 501140 363470
rect 501996 363470 502030 363504
rect 501106 363346 501140 363380
rect 501106 363256 501140 363290
rect 501106 363166 501140 363200
rect 501106 363076 501140 363110
rect 501106 362986 501140 363020
rect 501106 362896 501140 362930
rect 501106 362806 501140 362840
rect 501996 363380 502030 363414
rect 501996 363290 502030 363324
rect 501996 363200 502030 363234
rect 501996 363110 502030 363144
rect 501996 363020 502030 363054
rect 501996 362930 502030 362964
rect 501996 362840 502030 362874
rect 501106 362716 501140 362750
rect 501996 362750 502030 362784
rect 501182 362658 501216 362692
rect 501272 362658 501306 362692
rect 501362 362658 501396 362692
rect 501452 362658 501486 362692
rect 501542 362658 501576 362692
rect 501632 362658 501666 362692
rect 501722 362658 501756 362692
rect 501812 362658 501846 362692
rect 501902 362658 501936 362692
rect 504923 372928 504957 372962
rect 505013 372928 505047 372962
rect 505103 372928 505137 372962
rect 505193 372928 505227 372962
rect 505283 372928 505317 372962
rect 505373 372928 505407 372962
rect 505463 372928 505497 372962
rect 505553 372928 505587 372962
rect 505643 372928 505677 372962
rect 504866 372816 504900 372850
rect 505756 372850 505790 372884
rect 504866 372726 504900 372760
rect 504866 372636 504900 372670
rect 504866 372546 504900 372580
rect 504866 372456 504900 372490
rect 504866 372366 504900 372400
rect 504866 372276 504900 372310
rect 504866 372186 504900 372220
rect 505756 372760 505790 372794
rect 505756 372670 505790 372704
rect 505756 372580 505790 372614
rect 505756 372490 505790 372524
rect 505756 372400 505790 372434
rect 505756 372310 505790 372344
rect 505756 372220 505790 372254
rect 504866 372096 504900 372130
rect 505756 372130 505790 372164
rect 504942 372038 504976 372072
rect 505032 372038 505066 372072
rect 505122 372038 505156 372072
rect 505212 372038 505246 372072
rect 505302 372038 505336 372072
rect 505392 372038 505426 372072
rect 505482 372038 505516 372072
rect 505572 372038 505606 372072
rect 505662 372038 505696 372072
rect 504923 371588 504957 371622
rect 505013 371588 505047 371622
rect 505103 371588 505137 371622
rect 505193 371588 505227 371622
rect 505283 371588 505317 371622
rect 505373 371588 505407 371622
rect 505463 371588 505497 371622
rect 505553 371588 505587 371622
rect 505643 371588 505677 371622
rect 504866 371476 504900 371510
rect 505756 371510 505790 371544
rect 504866 371386 504900 371420
rect 504866 371296 504900 371330
rect 504866 371206 504900 371240
rect 504866 371116 504900 371150
rect 504866 371026 504900 371060
rect 504866 370936 504900 370970
rect 504866 370846 504900 370880
rect 505756 371420 505790 371454
rect 505756 371330 505790 371364
rect 505756 371240 505790 371274
rect 505756 371150 505790 371184
rect 505756 371060 505790 371094
rect 505756 370970 505790 371004
rect 505756 370880 505790 370914
rect 504866 370756 504900 370790
rect 505756 370790 505790 370824
rect 504942 370698 504976 370732
rect 505032 370698 505066 370732
rect 505122 370698 505156 370732
rect 505212 370698 505246 370732
rect 505302 370698 505336 370732
rect 505392 370698 505426 370732
rect 505482 370698 505516 370732
rect 505572 370698 505606 370732
rect 505662 370698 505696 370732
rect 504923 370248 504957 370282
rect 505013 370248 505047 370282
rect 505103 370248 505137 370282
rect 505193 370248 505227 370282
rect 505283 370248 505317 370282
rect 505373 370248 505407 370282
rect 505463 370248 505497 370282
rect 505553 370248 505587 370282
rect 505643 370248 505677 370282
rect 504866 370136 504900 370170
rect 505756 370170 505790 370204
rect 504866 370046 504900 370080
rect 504866 369956 504900 369990
rect 504866 369866 504900 369900
rect 504866 369776 504900 369810
rect 504866 369686 504900 369720
rect 504866 369596 504900 369630
rect 504866 369506 504900 369540
rect 505756 370080 505790 370114
rect 505756 369990 505790 370024
rect 505756 369900 505790 369934
rect 505756 369810 505790 369844
rect 505756 369720 505790 369754
rect 505756 369630 505790 369664
rect 505756 369540 505790 369574
rect 504866 369416 504900 369450
rect 505756 369450 505790 369484
rect 504942 369358 504976 369392
rect 505032 369358 505066 369392
rect 505122 369358 505156 369392
rect 505212 369358 505246 369392
rect 505302 369358 505336 369392
rect 505392 369358 505426 369392
rect 505482 369358 505516 369392
rect 505572 369358 505606 369392
rect 505662 369358 505696 369392
rect 504923 368908 504957 368942
rect 505013 368908 505047 368942
rect 505103 368908 505137 368942
rect 505193 368908 505227 368942
rect 505283 368908 505317 368942
rect 505373 368908 505407 368942
rect 505463 368908 505497 368942
rect 505553 368908 505587 368942
rect 505643 368908 505677 368942
rect 504866 368796 504900 368830
rect 505756 368830 505790 368864
rect 504866 368706 504900 368740
rect 504866 368616 504900 368650
rect 504866 368526 504900 368560
rect 504866 368436 504900 368470
rect 504866 368346 504900 368380
rect 504866 368256 504900 368290
rect 504866 368166 504900 368200
rect 505756 368740 505790 368774
rect 505756 368650 505790 368684
rect 505756 368560 505790 368594
rect 505756 368470 505790 368504
rect 505756 368380 505790 368414
rect 505756 368290 505790 368324
rect 505756 368200 505790 368234
rect 504866 368076 504900 368110
rect 505756 368110 505790 368144
rect 504942 368018 504976 368052
rect 505032 368018 505066 368052
rect 505122 368018 505156 368052
rect 505212 368018 505246 368052
rect 505302 368018 505336 368052
rect 505392 368018 505426 368052
rect 505482 368018 505516 368052
rect 505572 368018 505606 368052
rect 505662 368018 505696 368052
rect 504923 367568 504957 367602
rect 505013 367568 505047 367602
rect 505103 367568 505137 367602
rect 505193 367568 505227 367602
rect 505283 367568 505317 367602
rect 505373 367568 505407 367602
rect 505463 367568 505497 367602
rect 505553 367568 505587 367602
rect 505643 367568 505677 367602
rect 504866 367456 504900 367490
rect 505756 367490 505790 367524
rect 504866 367366 504900 367400
rect 504866 367276 504900 367310
rect 504866 367186 504900 367220
rect 504866 367096 504900 367130
rect 504866 367006 504900 367040
rect 504866 366916 504900 366950
rect 504866 366826 504900 366860
rect 505756 367400 505790 367434
rect 505756 367310 505790 367344
rect 505756 367220 505790 367254
rect 505756 367130 505790 367164
rect 505756 367040 505790 367074
rect 505756 366950 505790 366984
rect 505756 366860 505790 366894
rect 504866 366736 504900 366770
rect 505756 366770 505790 366804
rect 504942 366678 504976 366712
rect 505032 366678 505066 366712
rect 505122 366678 505156 366712
rect 505212 366678 505246 366712
rect 505302 366678 505336 366712
rect 505392 366678 505426 366712
rect 505482 366678 505516 366712
rect 505572 366678 505606 366712
rect 505662 366678 505696 366712
rect 504923 366228 504957 366262
rect 505013 366228 505047 366262
rect 505103 366228 505137 366262
rect 505193 366228 505227 366262
rect 505283 366228 505317 366262
rect 505373 366228 505407 366262
rect 505463 366228 505497 366262
rect 505553 366228 505587 366262
rect 505643 366228 505677 366262
rect 504866 366116 504900 366150
rect 505756 366150 505790 366184
rect 504866 366026 504900 366060
rect 504866 365936 504900 365970
rect 504866 365846 504900 365880
rect 504866 365756 504900 365790
rect 504866 365666 504900 365700
rect 504866 365576 504900 365610
rect 504866 365486 504900 365520
rect 505756 366060 505790 366094
rect 505756 365970 505790 366004
rect 505756 365880 505790 365914
rect 505756 365790 505790 365824
rect 505756 365700 505790 365734
rect 505756 365610 505790 365644
rect 505756 365520 505790 365554
rect 504866 365396 504900 365430
rect 505756 365430 505790 365464
rect 504942 365338 504976 365372
rect 505032 365338 505066 365372
rect 505122 365338 505156 365372
rect 505212 365338 505246 365372
rect 505302 365338 505336 365372
rect 505392 365338 505426 365372
rect 505482 365338 505516 365372
rect 505572 365338 505606 365372
rect 505662 365338 505696 365372
rect 504923 364888 504957 364922
rect 505013 364888 505047 364922
rect 505103 364888 505137 364922
rect 505193 364888 505227 364922
rect 505283 364888 505317 364922
rect 505373 364888 505407 364922
rect 505463 364888 505497 364922
rect 505553 364888 505587 364922
rect 505643 364888 505677 364922
rect 504866 364776 504900 364810
rect 505756 364810 505790 364844
rect 504866 364686 504900 364720
rect 504866 364596 504900 364630
rect 504866 364506 504900 364540
rect 504866 364416 504900 364450
rect 504866 364326 504900 364360
rect 504866 364236 504900 364270
rect 504866 364146 504900 364180
rect 505756 364720 505790 364754
rect 505756 364630 505790 364664
rect 505756 364540 505790 364574
rect 505756 364450 505790 364484
rect 505756 364360 505790 364394
rect 505756 364270 505790 364304
rect 505756 364180 505790 364214
rect 504866 364056 504900 364090
rect 505756 364090 505790 364124
rect 504942 363998 504976 364032
rect 505032 363998 505066 364032
rect 505122 363998 505156 364032
rect 505212 363998 505246 364032
rect 505302 363998 505336 364032
rect 505392 363998 505426 364032
rect 505482 363998 505516 364032
rect 505572 363998 505606 364032
rect 505662 363998 505696 364032
rect 504923 363548 504957 363582
rect 505013 363548 505047 363582
rect 505103 363548 505137 363582
rect 505193 363548 505227 363582
rect 505283 363548 505317 363582
rect 505373 363548 505407 363582
rect 505463 363548 505497 363582
rect 505553 363548 505587 363582
rect 505643 363548 505677 363582
rect 504866 363436 504900 363470
rect 505756 363470 505790 363504
rect 504866 363346 504900 363380
rect 504866 363256 504900 363290
rect 504866 363166 504900 363200
rect 504866 363076 504900 363110
rect 504866 362986 504900 363020
rect 504866 362896 504900 362930
rect 504866 362806 504900 362840
rect 505756 363380 505790 363414
rect 505756 363290 505790 363324
rect 505756 363200 505790 363234
rect 505756 363110 505790 363144
rect 505756 363020 505790 363054
rect 505756 362930 505790 362964
rect 505756 362840 505790 362874
rect 504866 362716 504900 362750
rect 505756 362750 505790 362784
rect 504942 362658 504976 362692
rect 505032 362658 505066 362692
rect 505122 362658 505156 362692
rect 505212 362658 505246 362692
rect 505302 362658 505336 362692
rect 505392 362658 505426 362692
rect 505482 362658 505516 362692
rect 505572 362658 505606 362692
rect 505662 362658 505696 362692
rect 508683 372928 508717 372962
rect 508773 372928 508807 372962
rect 508863 372928 508897 372962
rect 508953 372928 508987 372962
rect 509043 372928 509077 372962
rect 509133 372928 509167 372962
rect 509223 372928 509257 372962
rect 509313 372928 509347 372962
rect 509403 372928 509437 372962
rect 508626 372816 508660 372850
rect 509516 372850 509550 372884
rect 508626 372726 508660 372760
rect 508626 372636 508660 372670
rect 508626 372546 508660 372580
rect 508626 372456 508660 372490
rect 508626 372366 508660 372400
rect 508626 372276 508660 372310
rect 508626 372186 508660 372220
rect 509516 372760 509550 372794
rect 509516 372670 509550 372704
rect 509516 372580 509550 372614
rect 509516 372490 509550 372524
rect 509516 372400 509550 372434
rect 509516 372310 509550 372344
rect 509516 372220 509550 372254
rect 508626 372096 508660 372130
rect 509516 372130 509550 372164
rect 508702 372038 508736 372072
rect 508792 372038 508826 372072
rect 508882 372038 508916 372072
rect 508972 372038 509006 372072
rect 509062 372038 509096 372072
rect 509152 372038 509186 372072
rect 509242 372038 509276 372072
rect 509332 372038 509366 372072
rect 509422 372038 509456 372072
rect 508683 371588 508717 371622
rect 508773 371588 508807 371622
rect 508863 371588 508897 371622
rect 508953 371588 508987 371622
rect 509043 371588 509077 371622
rect 509133 371588 509167 371622
rect 509223 371588 509257 371622
rect 509313 371588 509347 371622
rect 509403 371588 509437 371622
rect 508626 371476 508660 371510
rect 509516 371510 509550 371544
rect 508626 371386 508660 371420
rect 508626 371296 508660 371330
rect 508626 371206 508660 371240
rect 508626 371116 508660 371150
rect 508626 371026 508660 371060
rect 508626 370936 508660 370970
rect 508626 370846 508660 370880
rect 509516 371420 509550 371454
rect 509516 371330 509550 371364
rect 509516 371240 509550 371274
rect 509516 371150 509550 371184
rect 509516 371060 509550 371094
rect 509516 370970 509550 371004
rect 509516 370880 509550 370914
rect 508626 370756 508660 370790
rect 509516 370790 509550 370824
rect 508702 370698 508736 370732
rect 508792 370698 508826 370732
rect 508882 370698 508916 370732
rect 508972 370698 509006 370732
rect 509062 370698 509096 370732
rect 509152 370698 509186 370732
rect 509242 370698 509276 370732
rect 509332 370698 509366 370732
rect 509422 370698 509456 370732
rect 508683 370248 508717 370282
rect 508773 370248 508807 370282
rect 508863 370248 508897 370282
rect 508953 370248 508987 370282
rect 509043 370248 509077 370282
rect 509133 370248 509167 370282
rect 509223 370248 509257 370282
rect 509313 370248 509347 370282
rect 509403 370248 509437 370282
rect 508626 370136 508660 370170
rect 509516 370170 509550 370204
rect 508626 370046 508660 370080
rect 508626 369956 508660 369990
rect 508626 369866 508660 369900
rect 508626 369776 508660 369810
rect 508626 369686 508660 369720
rect 508626 369596 508660 369630
rect 508626 369506 508660 369540
rect 509516 370080 509550 370114
rect 509516 369990 509550 370024
rect 509516 369900 509550 369934
rect 509516 369810 509550 369844
rect 509516 369720 509550 369754
rect 509516 369630 509550 369664
rect 509516 369540 509550 369574
rect 508626 369416 508660 369450
rect 509516 369450 509550 369484
rect 508702 369358 508736 369392
rect 508792 369358 508826 369392
rect 508882 369358 508916 369392
rect 508972 369358 509006 369392
rect 509062 369358 509096 369392
rect 509152 369358 509186 369392
rect 509242 369358 509276 369392
rect 509332 369358 509366 369392
rect 509422 369358 509456 369392
rect 508683 368908 508717 368942
rect 508773 368908 508807 368942
rect 508863 368908 508897 368942
rect 508953 368908 508987 368942
rect 509043 368908 509077 368942
rect 509133 368908 509167 368942
rect 509223 368908 509257 368942
rect 509313 368908 509347 368942
rect 509403 368908 509437 368942
rect 508626 368796 508660 368830
rect 509516 368830 509550 368864
rect 508626 368706 508660 368740
rect 508626 368616 508660 368650
rect 508626 368526 508660 368560
rect 508626 368436 508660 368470
rect 508626 368346 508660 368380
rect 508626 368256 508660 368290
rect 508626 368166 508660 368200
rect 509516 368740 509550 368774
rect 509516 368650 509550 368684
rect 509516 368560 509550 368594
rect 509516 368470 509550 368504
rect 509516 368380 509550 368414
rect 509516 368290 509550 368324
rect 509516 368200 509550 368234
rect 508626 368076 508660 368110
rect 509516 368110 509550 368144
rect 508702 368018 508736 368052
rect 508792 368018 508826 368052
rect 508882 368018 508916 368052
rect 508972 368018 509006 368052
rect 509062 368018 509096 368052
rect 509152 368018 509186 368052
rect 509242 368018 509276 368052
rect 509332 368018 509366 368052
rect 509422 368018 509456 368052
rect 508683 367568 508717 367602
rect 508773 367568 508807 367602
rect 508863 367568 508897 367602
rect 508953 367568 508987 367602
rect 509043 367568 509077 367602
rect 509133 367568 509167 367602
rect 509223 367568 509257 367602
rect 509313 367568 509347 367602
rect 509403 367568 509437 367602
rect 508626 367456 508660 367490
rect 509516 367490 509550 367524
rect 508626 367366 508660 367400
rect 508626 367276 508660 367310
rect 508626 367186 508660 367220
rect 508626 367096 508660 367130
rect 508626 367006 508660 367040
rect 508626 366916 508660 366950
rect 508626 366826 508660 366860
rect 509516 367400 509550 367434
rect 509516 367310 509550 367344
rect 509516 367220 509550 367254
rect 509516 367130 509550 367164
rect 509516 367040 509550 367074
rect 509516 366950 509550 366984
rect 509516 366860 509550 366894
rect 508626 366736 508660 366770
rect 509516 366770 509550 366804
rect 508702 366678 508736 366712
rect 508792 366678 508826 366712
rect 508882 366678 508916 366712
rect 508972 366678 509006 366712
rect 509062 366678 509096 366712
rect 509152 366678 509186 366712
rect 509242 366678 509276 366712
rect 509332 366678 509366 366712
rect 509422 366678 509456 366712
rect 508683 366228 508717 366262
rect 508773 366228 508807 366262
rect 508863 366228 508897 366262
rect 508953 366228 508987 366262
rect 509043 366228 509077 366262
rect 509133 366228 509167 366262
rect 509223 366228 509257 366262
rect 509313 366228 509347 366262
rect 509403 366228 509437 366262
rect 508626 366116 508660 366150
rect 509516 366150 509550 366184
rect 508626 366026 508660 366060
rect 508626 365936 508660 365970
rect 508626 365846 508660 365880
rect 508626 365756 508660 365790
rect 508626 365666 508660 365700
rect 508626 365576 508660 365610
rect 508626 365486 508660 365520
rect 509516 366060 509550 366094
rect 509516 365970 509550 366004
rect 509516 365880 509550 365914
rect 509516 365790 509550 365824
rect 509516 365700 509550 365734
rect 509516 365610 509550 365644
rect 509516 365520 509550 365554
rect 508626 365396 508660 365430
rect 509516 365430 509550 365464
rect 508702 365338 508736 365372
rect 508792 365338 508826 365372
rect 508882 365338 508916 365372
rect 508972 365338 509006 365372
rect 509062 365338 509096 365372
rect 509152 365338 509186 365372
rect 509242 365338 509276 365372
rect 509332 365338 509366 365372
rect 509422 365338 509456 365372
rect 508683 364888 508717 364922
rect 508773 364888 508807 364922
rect 508863 364888 508897 364922
rect 508953 364888 508987 364922
rect 509043 364888 509077 364922
rect 509133 364888 509167 364922
rect 509223 364888 509257 364922
rect 509313 364888 509347 364922
rect 509403 364888 509437 364922
rect 508626 364776 508660 364810
rect 509516 364810 509550 364844
rect 508626 364686 508660 364720
rect 508626 364596 508660 364630
rect 508626 364506 508660 364540
rect 508626 364416 508660 364450
rect 508626 364326 508660 364360
rect 508626 364236 508660 364270
rect 508626 364146 508660 364180
rect 509516 364720 509550 364754
rect 509516 364630 509550 364664
rect 509516 364540 509550 364574
rect 509516 364450 509550 364484
rect 509516 364360 509550 364394
rect 509516 364270 509550 364304
rect 509516 364180 509550 364214
rect 508626 364056 508660 364090
rect 509516 364090 509550 364124
rect 508702 363998 508736 364032
rect 508792 363998 508826 364032
rect 508882 363998 508916 364032
rect 508972 363998 509006 364032
rect 509062 363998 509096 364032
rect 509152 363998 509186 364032
rect 509242 363998 509276 364032
rect 509332 363998 509366 364032
rect 509422 363998 509456 364032
rect 508683 363548 508717 363582
rect 508773 363548 508807 363582
rect 508863 363548 508897 363582
rect 508953 363548 508987 363582
rect 509043 363548 509077 363582
rect 509133 363548 509167 363582
rect 509223 363548 509257 363582
rect 509313 363548 509347 363582
rect 509403 363548 509437 363582
rect 508626 363436 508660 363470
rect 509516 363470 509550 363504
rect 508626 363346 508660 363380
rect 508626 363256 508660 363290
rect 508626 363166 508660 363200
rect 508626 363076 508660 363110
rect 508626 362986 508660 363020
rect 508626 362896 508660 362930
rect 508626 362806 508660 362840
rect 509516 363380 509550 363414
rect 509516 363290 509550 363324
rect 509516 363200 509550 363234
rect 509516 363110 509550 363144
rect 509516 363020 509550 363054
rect 509516 362930 509550 362964
rect 509516 362840 509550 362874
rect 508626 362716 508660 362750
rect 509516 362750 509550 362784
rect 508702 362658 508736 362692
rect 508792 362658 508826 362692
rect 508882 362658 508916 362692
rect 508972 362658 509006 362692
rect 509062 362658 509096 362692
rect 509152 362658 509186 362692
rect 509242 362658 509276 362692
rect 509332 362658 509366 362692
rect 509422 362658 509456 362692
rect 512443 372928 512477 372962
rect 512533 372928 512567 372962
rect 512623 372928 512657 372962
rect 512713 372928 512747 372962
rect 512803 372928 512837 372962
rect 512893 372928 512927 372962
rect 512983 372928 513017 372962
rect 513073 372928 513107 372962
rect 513163 372928 513197 372962
rect 512386 372816 512420 372850
rect 513276 372850 513310 372884
rect 512386 372726 512420 372760
rect 512386 372636 512420 372670
rect 512386 372546 512420 372580
rect 512386 372456 512420 372490
rect 512386 372366 512420 372400
rect 512386 372276 512420 372310
rect 512386 372186 512420 372220
rect 513276 372760 513310 372794
rect 513276 372670 513310 372704
rect 513276 372580 513310 372614
rect 513276 372490 513310 372524
rect 513276 372400 513310 372434
rect 513276 372310 513310 372344
rect 513276 372220 513310 372254
rect 512386 372096 512420 372130
rect 513276 372130 513310 372164
rect 512462 372038 512496 372072
rect 512552 372038 512586 372072
rect 512642 372038 512676 372072
rect 512732 372038 512766 372072
rect 512822 372038 512856 372072
rect 512912 372038 512946 372072
rect 513002 372038 513036 372072
rect 513092 372038 513126 372072
rect 513182 372038 513216 372072
rect 523261 374747 523295 374781
rect 523261 373447 523295 373481
rect 523261 372147 523295 372181
rect 512443 371588 512477 371622
rect 512533 371588 512567 371622
rect 512623 371588 512657 371622
rect 512713 371588 512747 371622
rect 512803 371588 512837 371622
rect 512893 371588 512927 371622
rect 512983 371588 513017 371622
rect 513073 371588 513107 371622
rect 513163 371588 513197 371622
rect 512386 371476 512420 371510
rect 513276 371510 513310 371544
rect 512386 371386 512420 371420
rect 512386 371296 512420 371330
rect 512386 371206 512420 371240
rect 512386 371116 512420 371150
rect 512386 371026 512420 371060
rect 512386 370936 512420 370970
rect 512386 370846 512420 370880
rect 513276 371420 513310 371454
rect 513276 371330 513310 371364
rect 513276 371240 513310 371274
rect 513276 371150 513310 371184
rect 513276 371060 513310 371094
rect 513276 370970 513310 371004
rect 513276 370880 513310 370914
rect 512386 370756 512420 370790
rect 513276 370790 513310 370824
rect 512462 370698 512496 370732
rect 512552 370698 512586 370732
rect 512642 370698 512676 370732
rect 512732 370698 512766 370732
rect 512822 370698 512856 370732
rect 512912 370698 512946 370732
rect 513002 370698 513036 370732
rect 513092 370698 513126 370732
rect 513182 370698 513216 370732
rect 512443 370248 512477 370282
rect 512533 370248 512567 370282
rect 512623 370248 512657 370282
rect 512713 370248 512747 370282
rect 512803 370248 512837 370282
rect 512893 370248 512927 370282
rect 512983 370248 513017 370282
rect 513073 370248 513107 370282
rect 513163 370248 513197 370282
rect 512386 370136 512420 370170
rect 513276 370170 513310 370204
rect 512386 370046 512420 370080
rect 512386 369956 512420 369990
rect 512386 369866 512420 369900
rect 512386 369776 512420 369810
rect 512386 369686 512420 369720
rect 512386 369596 512420 369630
rect 512386 369506 512420 369540
rect 513276 370080 513310 370114
rect 513276 369990 513310 370024
rect 513276 369900 513310 369934
rect 513276 369810 513310 369844
rect 513276 369720 513310 369754
rect 513276 369630 513310 369664
rect 513276 369540 513310 369574
rect 512386 369416 512420 369450
rect 513276 369450 513310 369484
rect 512462 369358 512496 369392
rect 512552 369358 512586 369392
rect 512642 369358 512676 369392
rect 512732 369358 512766 369392
rect 512822 369358 512856 369392
rect 512912 369358 512946 369392
rect 513002 369358 513036 369392
rect 513092 369358 513126 369392
rect 513182 369358 513216 369392
rect 523261 370847 523295 370881
rect 523261 369547 523295 369581
rect 512443 368908 512477 368942
rect 512533 368908 512567 368942
rect 512623 368908 512657 368942
rect 512713 368908 512747 368942
rect 512803 368908 512837 368942
rect 512893 368908 512927 368942
rect 512983 368908 513017 368942
rect 513073 368908 513107 368942
rect 513163 368908 513197 368942
rect 512386 368796 512420 368830
rect 513276 368830 513310 368864
rect 512386 368706 512420 368740
rect 512386 368616 512420 368650
rect 512386 368526 512420 368560
rect 512386 368436 512420 368470
rect 512386 368346 512420 368380
rect 512386 368256 512420 368290
rect 512386 368166 512420 368200
rect 513276 368740 513310 368774
rect 513276 368650 513310 368684
rect 513276 368560 513310 368594
rect 513276 368470 513310 368504
rect 513276 368380 513310 368414
rect 513276 368290 513310 368324
rect 513276 368200 513310 368234
rect 512386 368076 512420 368110
rect 513276 368110 513310 368144
rect 512462 368018 512496 368052
rect 512552 368018 512586 368052
rect 512642 368018 512676 368052
rect 512732 368018 512766 368052
rect 512822 368018 512856 368052
rect 512912 368018 512946 368052
rect 513002 368018 513036 368052
rect 513092 368018 513126 368052
rect 513182 368018 513216 368052
rect 512443 367568 512477 367602
rect 512533 367568 512567 367602
rect 512623 367568 512657 367602
rect 512713 367568 512747 367602
rect 512803 367568 512837 367602
rect 512893 367568 512927 367602
rect 512983 367568 513017 367602
rect 513073 367568 513107 367602
rect 513163 367568 513197 367602
rect 512386 367456 512420 367490
rect 513276 367490 513310 367524
rect 512386 367366 512420 367400
rect 512386 367276 512420 367310
rect 512386 367186 512420 367220
rect 512386 367096 512420 367130
rect 512386 367006 512420 367040
rect 512386 366916 512420 366950
rect 512386 366826 512420 366860
rect 513276 367400 513310 367434
rect 513276 367310 513310 367344
rect 513276 367220 513310 367254
rect 513276 367130 513310 367164
rect 513276 367040 513310 367074
rect 513276 366950 513310 366984
rect 513276 366860 513310 366894
rect 512386 366736 512420 366770
rect 513276 366770 513310 366804
rect 512462 366678 512496 366712
rect 512552 366678 512586 366712
rect 512642 366678 512676 366712
rect 512732 366678 512766 366712
rect 512822 366678 512856 366712
rect 512912 366678 512946 366712
rect 513002 366678 513036 366712
rect 513092 366678 513126 366712
rect 513182 366678 513216 366712
rect 523261 368247 523295 368281
rect 523261 366947 523295 366981
rect 512443 366228 512477 366262
rect 512533 366228 512567 366262
rect 512623 366228 512657 366262
rect 512713 366228 512747 366262
rect 512803 366228 512837 366262
rect 512893 366228 512927 366262
rect 512983 366228 513017 366262
rect 513073 366228 513107 366262
rect 513163 366228 513197 366262
rect 512386 366116 512420 366150
rect 513276 366150 513310 366184
rect 512386 366026 512420 366060
rect 512386 365936 512420 365970
rect 512386 365846 512420 365880
rect 512386 365756 512420 365790
rect 512386 365666 512420 365700
rect 512386 365576 512420 365610
rect 512386 365486 512420 365520
rect 513276 366060 513310 366094
rect 513276 365970 513310 366004
rect 513276 365880 513310 365914
rect 513276 365790 513310 365824
rect 513276 365700 513310 365734
rect 513276 365610 513310 365644
rect 513276 365520 513310 365554
rect 512386 365396 512420 365430
rect 513276 365430 513310 365464
rect 512462 365338 512496 365372
rect 512552 365338 512586 365372
rect 512642 365338 512676 365372
rect 512732 365338 512766 365372
rect 512822 365338 512856 365372
rect 512912 365338 512946 365372
rect 513002 365338 513036 365372
rect 513092 365338 513126 365372
rect 513182 365338 513216 365372
rect 512443 364888 512477 364922
rect 512533 364888 512567 364922
rect 512623 364888 512657 364922
rect 512713 364888 512747 364922
rect 512803 364888 512837 364922
rect 512893 364888 512927 364922
rect 512983 364888 513017 364922
rect 513073 364888 513107 364922
rect 513163 364888 513197 364922
rect 512386 364776 512420 364810
rect 513276 364810 513310 364844
rect 512386 364686 512420 364720
rect 512386 364596 512420 364630
rect 512386 364506 512420 364540
rect 512386 364416 512420 364450
rect 512386 364326 512420 364360
rect 512386 364236 512420 364270
rect 512386 364146 512420 364180
rect 513276 364720 513310 364754
rect 513276 364630 513310 364664
rect 513276 364540 513310 364574
rect 513276 364450 513310 364484
rect 513276 364360 513310 364394
rect 513276 364270 513310 364304
rect 513276 364180 513310 364214
rect 512386 364056 512420 364090
rect 513276 364090 513310 364124
rect 512462 363998 512496 364032
rect 512552 363998 512586 364032
rect 512642 363998 512676 364032
rect 512732 363998 512766 364032
rect 512822 363998 512856 364032
rect 512912 363998 512946 364032
rect 513002 363998 513036 364032
rect 513092 363998 513126 364032
rect 513182 363998 513216 364032
rect 523261 365647 523295 365681
rect 523261 364347 523295 364381
rect 512443 363548 512477 363582
rect 512533 363548 512567 363582
rect 512623 363548 512657 363582
rect 512713 363548 512747 363582
rect 512803 363548 512837 363582
rect 512893 363548 512927 363582
rect 512983 363548 513017 363582
rect 513073 363548 513107 363582
rect 513163 363548 513197 363582
rect 512386 363436 512420 363470
rect 513276 363470 513310 363504
rect 512386 363346 512420 363380
rect 512386 363256 512420 363290
rect 512386 363166 512420 363200
rect 512386 363076 512420 363110
rect 512386 362986 512420 363020
rect 512386 362896 512420 362930
rect 512386 362806 512420 362840
rect 513276 363380 513310 363414
rect 513276 363290 513310 363324
rect 513276 363200 513310 363234
rect 513276 363110 513310 363144
rect 513276 363020 513310 363054
rect 513276 362930 513310 362964
rect 513276 362840 513310 362874
rect 512386 362716 512420 362750
rect 513276 362750 513310 362784
rect 512462 362658 512496 362692
rect 512552 362658 512586 362692
rect 512642 362658 512676 362692
rect 512732 362658 512766 362692
rect 512822 362658 512856 362692
rect 512912 362658 512946 362692
rect 513002 362658 513036 362692
rect 513092 362658 513126 362692
rect 513182 362658 513216 362692
rect 576250 359182 576294 359218
rect 577550 359182 577594 359218
rect 578850 359182 578894 359218
rect 579952 359130 579992 359170
rect 576698 313014 576742 313050
rect 577998 313014 578042 313050
rect 579298 313014 579342 313050
rect 580400 312962 580440 313002
<< poly >>
rect 560707 493440 560907 493466
rect 560965 493440 561165 493466
rect 561223 493440 561423 493466
rect 561481 493440 561681 493466
rect 561739 493440 561939 493466
rect 561997 493440 562197 493466
rect 562255 493440 562455 493466
rect 562513 493440 562713 493466
rect 562771 493440 562971 493466
rect 563029 493440 563229 493466
rect 563287 493440 563487 493466
rect 563545 493440 563745 493466
rect 563803 493440 564003 493466
rect 564061 493440 564261 493466
rect 564319 493440 564519 493466
rect 564577 493440 564777 493466
rect 564835 493440 565035 493466
rect 565093 493440 565293 493466
rect 565351 493440 565551 493466
rect 565609 493440 565809 493466
rect 575263 493214 575463 493240
rect 575521 493214 575721 493240
rect 575779 493214 575979 493240
rect 576037 493214 576237 493240
rect 576295 493214 576495 493240
rect 576553 493214 576753 493240
rect 576811 493214 577011 493240
rect 577069 493214 577269 493240
rect 577327 493214 577527 493240
rect 577585 493214 577785 493240
rect 577843 493214 578043 493240
rect 578101 493214 578301 493240
rect 578359 493214 578559 493240
rect 578617 493214 578817 493240
rect 578875 493214 579075 493240
rect 579133 493214 579333 493240
rect 579391 493214 579591 493240
rect 579649 493214 579849 493240
rect 579907 493214 580107 493240
rect 580165 493214 580365 493240
rect 560707 492414 560907 492440
rect 560965 492414 561165 492440
rect 561223 492414 561423 492440
rect 561481 492414 561681 492440
rect 561739 492414 561939 492440
rect 561997 492414 562197 492440
rect 562255 492414 562455 492440
rect 562513 492414 562713 492440
rect 562771 492414 562971 492440
rect 563029 492414 563229 492440
rect 563287 492414 563487 492440
rect 563545 492414 563745 492440
rect 563803 492414 564003 492440
rect 564061 492414 564261 492440
rect 564319 492414 564519 492440
rect 564577 492414 564777 492440
rect 564835 492414 565035 492440
rect 565093 492414 565293 492440
rect 565351 492414 565551 492440
rect 565609 492414 565809 492440
rect 560762 492224 560882 492414
rect 561018 492224 561138 492414
rect 561274 492224 561394 492414
rect 561530 492224 561650 492414
rect 561786 492224 561906 492414
rect 562042 492224 562162 492414
rect 562298 492224 562418 492414
rect 562554 492224 562674 492414
rect 562810 492224 562930 492414
rect 563066 492224 563186 492414
rect 563322 492224 563442 492414
rect 563578 492224 563698 492414
rect 563834 492224 563954 492414
rect 564090 492224 564210 492414
rect 564346 492224 564466 492414
rect 564602 492224 564722 492414
rect 564858 492224 564978 492414
rect 565114 492224 565234 492414
rect 565370 492224 565490 492414
rect 565626 492224 565746 492414
rect 560650 492204 565786 492224
rect 560650 492144 560836 492204
rect 560896 492144 561036 492204
rect 561096 492144 561236 492204
rect 561296 492144 561436 492204
rect 561496 492144 561636 492204
rect 561696 492144 561836 492204
rect 561896 492144 562036 492204
rect 562096 492144 562236 492204
rect 562296 492144 562436 492204
rect 562496 492144 562636 492204
rect 562696 492144 562836 492204
rect 562896 492144 563036 492204
rect 563096 492144 563236 492204
rect 563296 492144 563436 492204
rect 563496 492144 563636 492204
rect 563696 492144 563836 492204
rect 563896 492144 564036 492204
rect 564096 492144 564236 492204
rect 564296 492144 564436 492204
rect 564496 492144 564636 492204
rect 564696 492144 564836 492204
rect 564896 492144 565036 492204
rect 565096 492144 565236 492204
rect 565296 492144 565436 492204
rect 565496 492144 565636 492204
rect 565696 492144 565786 492204
rect 575263 492188 575463 492214
rect 575521 492188 575721 492214
rect 575779 492188 575979 492214
rect 576037 492188 576237 492214
rect 576295 492188 576495 492214
rect 576553 492188 576753 492214
rect 576811 492188 577011 492214
rect 577069 492188 577269 492214
rect 577327 492188 577527 492214
rect 577585 492188 577785 492214
rect 577843 492188 578043 492214
rect 578101 492188 578301 492214
rect 578359 492188 578559 492214
rect 578617 492188 578817 492214
rect 578875 492188 579075 492214
rect 579133 492188 579333 492214
rect 579391 492188 579591 492214
rect 579649 492188 579849 492214
rect 579907 492188 580107 492214
rect 580165 492188 580365 492214
rect 560650 492124 565786 492144
rect 575334 491942 575454 492188
rect 575590 491942 575710 492188
rect 575846 491942 575966 492188
rect 576102 491942 576222 492188
rect 576358 491942 576478 492188
rect 576614 491942 576734 492188
rect 576870 491942 576990 492188
rect 577126 491942 577246 492188
rect 577382 491942 577502 492188
rect 577638 491942 577758 492188
rect 577894 491942 578014 492188
rect 578150 491942 578270 492188
rect 578406 491942 578526 492188
rect 578662 491942 578782 492188
rect 578918 491942 579038 492188
rect 579174 491942 579294 492188
rect 579430 491942 579550 492188
rect 579686 491942 579806 492188
rect 579942 491942 580062 492188
rect 580198 491942 580318 492188
rect 575170 491922 580458 491942
rect 575170 491862 575228 491922
rect 575288 491862 575428 491922
rect 575488 491862 575628 491922
rect 575688 491862 575828 491922
rect 575888 491862 576028 491922
rect 576088 491862 576228 491922
rect 576288 491862 576428 491922
rect 576488 491862 576628 491922
rect 576688 491862 576828 491922
rect 576888 491862 577028 491922
rect 577088 491862 577228 491922
rect 577288 491862 577428 491922
rect 577488 491862 577628 491922
rect 577688 491862 577828 491922
rect 577888 491862 578028 491922
rect 578088 491862 578228 491922
rect 578288 491862 578428 491922
rect 578488 491862 578628 491922
rect 578688 491862 578828 491922
rect 578888 491862 579028 491922
rect 579088 491862 579228 491922
rect 579288 491862 579428 491922
rect 579488 491862 579628 491922
rect 579688 491862 579828 491922
rect 579888 491862 580028 491922
rect 580088 491862 580228 491922
rect 580288 491862 580458 491922
rect 575170 491842 580458 491862
rect 574541 404338 574741 404364
rect 574799 404338 574999 404364
rect 575057 404338 575257 404364
rect 575315 404338 575515 404364
rect 575573 404338 575773 404364
rect 575831 404338 576031 404364
rect 576089 404338 576289 404364
rect 576347 404338 576547 404364
rect 576605 404338 576805 404364
rect 576863 404338 577063 404364
rect 577121 404338 577321 404364
rect 577379 404338 577579 404364
rect 577637 404338 577837 404364
rect 577895 404338 578095 404364
rect 578153 404338 578353 404364
rect 578411 404338 578611 404364
rect 578669 404338 578869 404364
rect 578927 404338 579127 404364
rect 579185 404338 579385 404364
rect 579443 404338 579643 404364
rect 560747 404298 560947 404324
rect 561005 404298 561205 404324
rect 561263 404298 561463 404324
rect 561521 404298 561721 404324
rect 561779 404298 561979 404324
rect 562037 404298 562237 404324
rect 562295 404298 562495 404324
rect 562553 404298 562753 404324
rect 562811 404298 563011 404324
rect 563069 404298 563269 404324
rect 563327 404298 563527 404324
rect 563585 404298 563785 404324
rect 563843 404298 564043 404324
rect 564101 404298 564301 404324
rect 564359 404298 564559 404324
rect 564617 404298 564817 404324
rect 564875 404298 565075 404324
rect 565133 404298 565333 404324
rect 565391 404298 565591 404324
rect 565649 404298 565849 404324
rect 574541 403312 574741 403338
rect 574799 403312 574999 403338
rect 575057 403312 575257 403338
rect 575315 403312 575515 403338
rect 575573 403312 575773 403338
rect 575831 403312 576031 403338
rect 576089 403312 576289 403338
rect 576347 403312 576547 403338
rect 576605 403312 576805 403338
rect 576863 403312 577063 403338
rect 577121 403312 577321 403338
rect 577379 403312 577579 403338
rect 577637 403312 577837 403338
rect 577895 403312 578095 403338
rect 578153 403312 578353 403338
rect 578411 403312 578611 403338
rect 578669 403312 578869 403338
rect 578927 403312 579127 403338
rect 579185 403312 579385 403338
rect 579443 403312 579643 403338
rect 560747 403272 560947 403298
rect 561005 403272 561205 403298
rect 561263 403272 561463 403298
rect 561521 403272 561721 403298
rect 561779 403272 561979 403298
rect 562037 403272 562237 403298
rect 562295 403272 562495 403298
rect 562553 403272 562753 403298
rect 562811 403272 563011 403298
rect 563069 403272 563269 403298
rect 563327 403272 563527 403298
rect 563585 403272 563785 403298
rect 563843 403272 564043 403298
rect 564101 403272 564301 403298
rect 564359 403272 564559 403298
rect 564617 403272 564817 403298
rect 564875 403272 565075 403298
rect 565133 403272 565333 403298
rect 565391 403272 565591 403298
rect 565649 403272 565849 403298
rect 560810 403082 560930 403272
rect 561066 403082 561186 403272
rect 561322 403082 561442 403272
rect 561578 403082 561698 403272
rect 561834 403082 561954 403272
rect 562090 403082 562210 403272
rect 562346 403082 562466 403272
rect 562602 403082 562722 403272
rect 562858 403082 562978 403272
rect 563114 403082 563234 403272
rect 563370 403082 563490 403272
rect 563626 403082 563746 403272
rect 563882 403082 564002 403272
rect 564138 403082 564258 403272
rect 564394 403082 564514 403272
rect 564650 403082 564770 403272
rect 564906 403082 565026 403272
rect 565162 403082 565282 403272
rect 565418 403082 565538 403272
rect 565674 403082 565794 403272
rect 560770 403062 565906 403082
rect 574612 403066 574732 403312
rect 574868 403066 574988 403312
rect 575124 403066 575244 403312
rect 575380 403066 575500 403312
rect 575636 403066 575756 403312
rect 575892 403066 576012 403312
rect 576148 403066 576268 403312
rect 576404 403066 576524 403312
rect 576660 403066 576780 403312
rect 576916 403066 577036 403312
rect 577172 403066 577292 403312
rect 577428 403066 577548 403312
rect 577684 403066 577804 403312
rect 577940 403066 578060 403312
rect 578196 403066 578316 403312
rect 578452 403066 578572 403312
rect 578708 403066 578828 403312
rect 578964 403066 579084 403312
rect 579220 403066 579340 403312
rect 579476 403066 579596 403312
rect 560770 403002 560860 403062
rect 560920 403002 561060 403062
rect 561120 403002 561260 403062
rect 561320 403002 561460 403062
rect 561520 403002 561660 403062
rect 561720 403002 561860 403062
rect 561920 403002 562060 403062
rect 562120 403002 562260 403062
rect 562320 403002 562460 403062
rect 562520 403002 562660 403062
rect 562720 403002 562860 403062
rect 562920 403002 563060 403062
rect 563120 403002 563260 403062
rect 563320 403002 563460 403062
rect 563520 403002 563660 403062
rect 563720 403002 563860 403062
rect 563920 403002 564060 403062
rect 564120 403002 564260 403062
rect 564320 403002 564460 403062
rect 564520 403002 564660 403062
rect 564720 403002 564860 403062
rect 564920 403002 565060 403062
rect 565120 403002 565260 403062
rect 565320 403002 565460 403062
rect 565520 403002 565660 403062
rect 565720 403002 565906 403062
rect 560770 402982 565906 403002
rect 574448 403046 579736 403066
rect 574448 402986 574506 403046
rect 574566 402986 574706 403046
rect 574766 402986 574906 403046
rect 574966 402986 575106 403046
rect 575166 402986 575306 403046
rect 575366 402986 575506 403046
rect 575566 402986 575706 403046
rect 575766 402986 575906 403046
rect 575966 402986 576106 403046
rect 576166 402986 576306 403046
rect 576366 402986 576506 403046
rect 576566 402986 576706 403046
rect 576766 402986 576906 403046
rect 576966 402986 577106 403046
rect 577166 402986 577306 403046
rect 577366 402986 577506 403046
rect 577566 402986 577706 403046
rect 577766 402986 577906 403046
rect 577966 402986 578106 403046
rect 578166 402986 578306 403046
rect 578366 402986 578506 403046
rect 578566 402986 578706 403046
rect 578766 402986 578906 403046
rect 578966 402986 579106 403046
rect 579166 402986 579306 403046
rect 579366 402986 579506 403046
rect 579566 402986 579736 403046
rect 574448 402966 579736 402986
rect 497322 400378 497348 400778
rect 498148 400630 498174 400778
rect 498524 400653 498624 400756
rect 498524 400630 498557 400653
rect 498148 400619 498557 400630
rect 498591 400619 498624 400653
rect 498148 400510 498624 400619
rect 498148 400378 498174 400510
rect 498524 400320 498624 400510
rect 497077 399431 497103 399831
rect 498393 399684 498419 399831
rect 498564 399741 498664 399924
rect 498564 399707 498597 399741
rect 498631 399707 498664 399741
rect 498564 399684 498664 399707
rect 498393 399564 498664 399684
rect 498393 399431 498419 399564
rect 497077 398973 497103 399373
rect 498393 399228 498419 399373
rect 498564 399341 498664 399564
rect 498564 399307 498597 399341
rect 498631 399307 498664 399341
rect 498564 399228 498664 399307
rect 498393 399108 498664 399228
rect 498393 398973 498419 399108
rect 498564 398941 498664 399108
rect 497077 398515 497103 398915
rect 498393 398772 498419 398915
rect 498564 398907 498597 398941
rect 498631 398907 498664 398941
rect 498564 398772 498664 398907
rect 498393 398652 498664 398772
rect 498393 398515 498419 398652
rect 498564 398541 498664 398652
rect 498564 398507 498597 398541
rect 498631 398507 498664 398541
rect 497077 398057 497103 398457
rect 498393 398316 498419 398457
rect 498564 398316 498664 398507
rect 498393 398196 498664 398316
rect 498393 398057 498419 398196
rect 498564 398141 498664 398196
rect 498564 398107 498597 398141
rect 498631 398107 498664 398141
rect 497077 397599 497103 397999
rect 498393 397860 498419 397999
rect 498564 397860 498664 398107
rect 498393 397741 498664 397860
rect 498393 397740 498597 397741
rect 498393 397599 498419 397740
rect 498564 397707 498597 397740
rect 498631 397707 498664 397741
rect 497077 397141 497103 397541
rect 498393 397404 498419 397541
rect 498564 397404 498664 397707
rect 498393 397341 498664 397404
rect 498393 397307 498597 397341
rect 498631 397307 498664 397341
rect 498393 397284 498664 397307
rect 498393 397141 498419 397284
rect 497077 396683 497103 397083
rect 498393 396948 498419 397083
rect 498564 396948 498664 397284
rect 498393 396941 498664 396948
rect 498393 396907 498597 396941
rect 498631 396907 498664 396941
rect 498393 396828 498664 396907
rect 498393 396683 498419 396828
rect 497077 396225 497103 396625
rect 498393 396492 498419 396625
rect 498564 396541 498664 396828
rect 498564 396507 498597 396541
rect 498631 396507 498664 396541
rect 498564 396492 498664 396507
rect 498393 396372 498664 396492
rect 498393 396225 498419 396372
rect 497077 395767 497103 396167
rect 498393 396036 498419 396167
rect 498564 396141 498664 396372
rect 498564 396107 498597 396141
rect 498631 396107 498664 396141
rect 498564 396036 498664 396107
rect 498393 395916 498664 396036
rect 498393 395767 498419 395916
rect 498564 395741 498664 395916
rect 497077 395309 497103 395709
rect 498393 395580 498419 395709
rect 498564 395707 498597 395741
rect 498631 395707 498664 395741
rect 498564 395580 498664 395707
rect 498393 395460 498664 395580
rect 498393 395309 498419 395460
rect 498564 395341 498664 395460
rect 498564 395307 498597 395341
rect 498631 395307 498664 395341
rect 497077 394851 497103 395251
rect 498393 395124 498419 395251
rect 498564 395124 498664 395307
rect 498393 395004 498664 395124
rect 498393 394851 498419 395004
rect 498564 394941 498664 395004
rect 498564 394907 498597 394941
rect 498631 394907 498664 394941
rect 497077 394393 497103 394793
rect 498393 394668 498419 394793
rect 498564 394668 498664 394907
rect 498393 394548 498664 394668
rect 498393 394393 498419 394548
rect 498564 394541 498664 394548
rect 498564 394507 498597 394541
rect 498631 394507 498664 394541
rect 497077 393935 497103 394335
rect 498393 394212 498419 394335
rect 498564 394212 498664 394507
rect 498393 394141 498664 394212
rect 498393 394107 498597 394141
rect 498631 394107 498664 394141
rect 498393 394092 498664 394107
rect 498393 393935 498419 394092
rect 497077 393477 497103 393877
rect 498393 393756 498419 393877
rect 498564 393756 498664 394092
rect 498393 393741 498664 393756
rect 498393 393707 498597 393741
rect 498631 393707 498664 393741
rect 498393 393636 498664 393707
rect 498393 393477 498419 393636
rect 497077 393019 497103 393419
rect 498393 393300 498419 393419
rect 498564 393341 498664 393636
rect 498564 393307 498597 393341
rect 498631 393307 498664 393341
rect 498564 393300 498664 393307
rect 498393 393180 498664 393300
rect 498393 393019 498419 393180
rect 497077 392561 497103 392961
rect 498393 392844 498419 392961
rect 498564 392941 498664 393180
rect 498564 392907 498597 392941
rect 498631 392907 498664 392941
rect 498564 392844 498664 392907
rect 498393 392724 498664 392844
rect 498393 392561 498419 392724
rect 498564 392541 498664 392724
rect 498564 392507 498597 392541
rect 498631 392507 498664 392541
rect 497077 392103 497103 392503
rect 498393 392388 498419 392503
rect 498564 392388 498664 392507
rect 498393 392268 498664 392388
rect 498393 392103 498419 392268
rect 498564 392141 498664 392268
rect 498564 392107 498597 392141
rect 498631 392107 498664 392141
rect 497077 391645 497103 392045
rect 498393 391932 498419 392045
rect 498564 391932 498664 392107
rect 498393 391812 498664 391932
rect 498393 391645 498419 391812
rect 498564 391741 498664 391812
rect 500837 391787 500863 392187
rect 502153 392040 502179 392187
rect 502324 392097 502424 392280
rect 502324 392063 502357 392097
rect 502391 392063 502424 392097
rect 502324 392040 502424 392063
rect 502153 391920 502424 392040
rect 502153 391787 502179 391920
rect 498564 391707 498597 391741
rect 498631 391707 498664 391741
rect 497077 391187 497103 391587
rect 498393 391476 498419 391587
rect 498564 391476 498664 391707
rect 498393 391356 498664 391476
rect 498393 391187 498419 391356
rect 498564 391341 498664 391356
rect 498564 391307 498597 391341
rect 498631 391307 498664 391341
rect 500837 391329 500863 391729
rect 502153 391584 502179 391729
rect 502324 391697 502424 391920
rect 502324 391663 502357 391697
rect 502391 391663 502424 391697
rect 502324 391584 502424 391663
rect 502153 391464 502424 391584
rect 502153 391329 502179 391464
rect 493562 390578 493588 390978
rect 494388 390830 494414 390978
rect 494764 390853 494864 390956
rect 494764 390830 494797 390853
rect 494388 390819 494797 390830
rect 494831 390819 494864 390853
rect 494388 390710 494864 390819
rect 497077 390729 497103 391129
rect 498393 391020 498419 391129
rect 498564 391020 498664 391307
rect 502324 391297 502424 391464
rect 498393 390941 498664 391020
rect 498393 390907 498597 390941
rect 498631 390907 498664 390941
rect 498393 390900 498664 390907
rect 498393 390729 498419 390900
rect 494388 390578 494414 390710
rect 494764 390520 494864 390710
rect 497077 390271 497103 390671
rect 498393 390564 498419 390671
rect 498564 390564 498664 390900
rect 500837 390871 500863 391271
rect 502153 391128 502179 391271
rect 502324 391263 502357 391297
rect 502391 391263 502424 391297
rect 502324 391128 502424 391263
rect 502153 391008 502424 391128
rect 502153 390871 502179 391008
rect 502324 390897 502424 391008
rect 502324 390863 502357 390897
rect 502391 390863 502424 390897
rect 498393 390541 498664 390564
rect 498393 390507 498597 390541
rect 498631 390507 498664 390541
rect 498393 390444 498664 390507
rect 498393 390271 498419 390444
rect 493317 389631 493343 390031
rect 494633 389884 494659 390031
rect 494804 389941 494904 390124
rect 494804 389907 494837 389941
rect 494871 389907 494904 389941
rect 494804 389884 494904 389907
rect 494633 389764 494904 389884
rect 494633 389631 494659 389764
rect 493317 389173 493343 389573
rect 494633 389428 494659 389573
rect 494804 389541 494904 389764
rect 497077 389813 497103 390213
rect 498393 390108 498419 390213
rect 498564 390141 498664 390444
rect 500837 390413 500863 390813
rect 502153 390672 502179 390813
rect 502324 390672 502424 390863
rect 502153 390552 502424 390672
rect 502153 390413 502179 390552
rect 502324 390497 502424 390552
rect 502324 390463 502357 390497
rect 502391 390463 502424 390497
rect 498564 390108 498597 390141
rect 498393 390107 498597 390108
rect 498631 390107 498664 390141
rect 498393 389988 498664 390107
rect 498393 389813 498419 389988
rect 494804 389507 494837 389541
rect 494871 389507 494904 389541
rect 494804 389428 494904 389507
rect 494633 389308 494904 389428
rect 497077 389355 497103 389755
rect 498393 389652 498419 389755
rect 498564 389741 498664 389988
rect 500837 389955 500863 390355
rect 502153 390216 502179 390355
rect 502324 390216 502424 390463
rect 502153 390097 502424 390216
rect 502153 390096 502357 390097
rect 502153 389955 502179 390096
rect 502324 390063 502357 390096
rect 502391 390063 502424 390097
rect 498564 389707 498597 389741
rect 498631 389707 498664 389741
rect 498564 389652 498664 389707
rect 498393 389532 498664 389652
rect 498393 389355 498419 389532
rect 494633 389173 494659 389308
rect 494804 389141 494904 389308
rect 498564 389341 498664 389532
rect 500837 389497 500863 389897
rect 502153 389760 502179 389897
rect 502324 389760 502424 390063
rect 502153 389697 502424 389760
rect 502153 389663 502357 389697
rect 502391 389663 502424 389697
rect 502153 389640 502424 389663
rect 502153 389497 502179 389640
rect 498564 389307 498597 389341
rect 498631 389307 498664 389341
rect 493317 388715 493343 389115
rect 494633 388972 494659 389115
rect 494804 389107 494837 389141
rect 494871 389107 494904 389141
rect 494804 388972 494904 389107
rect 494633 388852 494904 388972
rect 497077 388897 497103 389297
rect 498393 389196 498419 389297
rect 498564 389196 498664 389307
rect 498393 389076 498664 389196
rect 498393 388897 498419 389076
rect 498564 388941 498664 389076
rect 500837 389039 500863 389439
rect 502153 389304 502179 389439
rect 502324 389304 502424 389640
rect 502153 389297 502424 389304
rect 502153 389263 502357 389297
rect 502391 389263 502424 389297
rect 502153 389184 502424 389263
rect 502153 389039 502179 389184
rect 498564 388907 498597 388941
rect 498631 388907 498664 388941
rect 494633 388715 494659 388852
rect 494804 388741 494904 388852
rect 494804 388707 494837 388741
rect 494871 388707 494904 388741
rect 493317 388257 493343 388657
rect 494633 388516 494659 388657
rect 494804 388516 494904 388707
rect 494633 388396 494904 388516
rect 497077 388439 497103 388839
rect 498393 388740 498419 388839
rect 498564 388740 498664 388907
rect 498393 388620 498664 388740
rect 498393 388439 498419 388620
rect 498564 388541 498664 388620
rect 500837 388581 500863 388981
rect 502153 388848 502179 388981
rect 502324 388897 502424 389184
rect 504842 389078 504868 389478
rect 505668 389330 505694 389478
rect 505884 389353 505984 389456
rect 505884 389330 505917 389353
rect 505668 389319 505917 389330
rect 505951 389319 505984 389353
rect 505668 389210 505984 389319
rect 505668 389078 505694 389210
rect 502324 388863 502357 388897
rect 502391 388863 502424 388897
rect 502324 388848 502424 388863
rect 502153 388728 502424 388848
rect 502153 388581 502179 388728
rect 498564 388507 498597 388541
rect 498631 388507 498664 388541
rect 494633 388257 494659 388396
rect 494804 388341 494904 388396
rect 494804 388307 494837 388341
rect 494871 388307 494904 388341
rect 493317 387799 493343 388199
rect 494633 388060 494659 388199
rect 494804 388060 494904 388307
rect 494633 387941 494904 388060
rect 497077 387981 497103 388381
rect 498393 388284 498419 388381
rect 498564 388284 498664 388507
rect 498393 388164 498664 388284
rect 498393 387981 498419 388164
rect 498564 388141 498664 388164
rect 498564 388107 498597 388141
rect 498631 388107 498664 388141
rect 500837 388123 500863 388523
rect 502153 388392 502179 388523
rect 502324 388497 502424 388728
rect 504842 388620 504868 389020
rect 505668 388874 505694 389020
rect 505884 388953 505984 389210
rect 516122 389078 516148 389478
rect 516948 389330 516974 389478
rect 517164 389353 517264 389456
rect 517164 389330 517197 389353
rect 516948 389319 517197 389330
rect 517231 389319 517264 389353
rect 516948 389210 517264 389319
rect 516948 389078 516974 389210
rect 505884 388919 505917 388953
rect 505951 388919 505984 388953
rect 505884 388874 505984 388919
rect 505668 388754 505984 388874
rect 505668 388620 505694 388754
rect 502324 388463 502357 388497
rect 502391 388463 502424 388497
rect 502324 388392 502424 388463
rect 502153 388272 502424 388392
rect 502153 388123 502179 388272
rect 494633 387940 494837 387941
rect 494633 387799 494659 387940
rect 494804 387907 494837 387940
rect 494871 387907 494904 387941
rect 493317 387341 493343 387741
rect 494633 387604 494659 387741
rect 494804 387604 494904 387907
rect 494633 387541 494904 387604
rect 494633 387507 494837 387541
rect 494871 387507 494904 387541
rect 497077 387523 497103 387923
rect 498393 387828 498419 387923
rect 498564 387828 498664 388107
rect 502324 388097 502424 388272
rect 504842 388162 504868 388562
rect 505668 388418 505694 388562
rect 505884 388553 505984 388754
rect 516122 388620 516148 389020
rect 516948 388874 516974 389020
rect 517164 388953 517264 389210
rect 517164 388919 517197 388953
rect 517231 388919 517264 388953
rect 517164 388874 517264 388919
rect 516948 388754 517264 388874
rect 516948 388620 516974 388754
rect 505884 388519 505917 388553
rect 505951 388519 505984 388553
rect 505884 388418 505984 388519
rect 505668 388298 505984 388418
rect 505668 388162 505694 388298
rect 505884 388153 505984 388298
rect 516122 388162 516148 388562
rect 516948 388418 516974 388562
rect 517164 388553 517264 388754
rect 523397 389631 523423 390031
rect 524713 389884 524739 390031
rect 524884 389941 524984 390124
rect 524884 389907 524917 389941
rect 524951 389907 524984 389941
rect 524884 389884 524984 389907
rect 524713 389764 524984 389884
rect 524713 389631 524739 389764
rect 523397 389173 523423 389573
rect 524713 389428 524739 389573
rect 524884 389541 524984 389764
rect 524884 389507 524917 389541
rect 524951 389507 524984 389541
rect 524884 389428 524984 389507
rect 524713 389308 524984 389428
rect 524713 389173 524739 389308
rect 524884 389141 524984 389308
rect 523397 388715 523423 389115
rect 524713 388972 524739 389115
rect 524884 389107 524917 389141
rect 524951 389107 524984 389141
rect 524884 388972 524984 389107
rect 524713 388852 524984 388972
rect 524713 388715 524739 388852
rect 524884 388741 524984 388852
rect 524884 388707 524917 388741
rect 524951 388707 524984 388741
rect 517164 388519 517197 388553
rect 517231 388519 517264 388553
rect 517164 388418 517264 388519
rect 516948 388298 517264 388418
rect 516948 388162 516974 388298
rect 505884 388119 505917 388153
rect 505951 388119 505984 388153
rect 498393 387741 498664 387828
rect 498393 387708 498597 387741
rect 498393 387523 498419 387708
rect 498564 387707 498597 387708
rect 498631 387707 498664 387741
rect 494633 387484 494904 387507
rect 494633 387341 494659 387484
rect 493317 386883 493343 387283
rect 494633 387148 494659 387283
rect 494804 387148 494904 387484
rect 494633 387141 494904 387148
rect 494633 387107 494837 387141
rect 494871 387107 494904 387141
rect 494633 387028 494904 387107
rect 497077 387065 497103 387465
rect 498393 387372 498419 387465
rect 498564 387372 498664 387707
rect 500837 387665 500863 388065
rect 502153 387936 502179 388065
rect 502324 388063 502357 388097
rect 502391 388063 502424 388097
rect 502324 387936 502424 388063
rect 502153 387816 502424 387936
rect 502153 387665 502179 387816
rect 502324 387697 502424 387816
rect 504842 387704 504868 388104
rect 505668 387962 505694 388104
rect 505884 387962 505984 388119
rect 517164 388153 517264 388298
rect 523397 388257 523423 388657
rect 524713 388516 524739 388657
rect 524884 388516 524984 388707
rect 524713 388396 524984 388516
rect 524713 388257 524739 388396
rect 524884 388341 524984 388396
rect 524884 388307 524917 388341
rect 524951 388307 524984 388341
rect 517164 388119 517197 388153
rect 517231 388119 517264 388153
rect 505668 387842 505984 387962
rect 505668 387704 505694 387842
rect 505884 387753 505984 387842
rect 505884 387719 505917 387753
rect 505951 387719 505984 387753
rect 502324 387663 502357 387697
rect 502391 387663 502424 387697
rect 498393 387341 498664 387372
rect 498393 387307 498597 387341
rect 498631 387307 498664 387341
rect 498393 387252 498664 387307
rect 498393 387065 498419 387252
rect 494633 386883 494659 387028
rect 493317 386425 493343 386825
rect 494633 386692 494659 386825
rect 494804 386741 494904 387028
rect 494804 386707 494837 386741
rect 494871 386707 494904 386741
rect 494804 386692 494904 386707
rect 494633 386572 494904 386692
rect 497077 386607 497103 387007
rect 498393 386916 498419 387007
rect 498564 386941 498664 387252
rect 500837 387207 500863 387607
rect 502153 387480 502179 387607
rect 502324 387480 502424 387663
rect 502153 387360 502424 387480
rect 502153 387207 502179 387360
rect 502324 387297 502424 387360
rect 502324 387263 502357 387297
rect 502391 387263 502424 387297
rect 498564 386916 498597 386941
rect 498393 386907 498597 386916
rect 498631 386907 498664 386941
rect 498393 386796 498664 386907
rect 498393 386607 498419 386796
rect 494633 386425 494659 386572
rect 493317 385967 493343 386367
rect 494633 386236 494659 386367
rect 494804 386341 494904 386572
rect 494804 386307 494837 386341
rect 494871 386307 494904 386341
rect 494804 386236 494904 386307
rect 494633 386116 494904 386236
rect 497077 386149 497103 386549
rect 498393 386460 498419 386549
rect 498564 386541 498664 386796
rect 500837 386749 500863 387149
rect 502153 387024 502179 387149
rect 502324 387024 502424 387263
rect 504842 387246 504868 387646
rect 505668 387506 505694 387646
rect 505884 387506 505984 387719
rect 505668 387386 505984 387506
rect 505668 387246 505694 387386
rect 505884 387353 505984 387386
rect 505884 387319 505917 387353
rect 505951 387319 505984 387353
rect 502153 386904 502424 387024
rect 502153 386749 502179 386904
rect 502324 386897 502424 386904
rect 502324 386863 502357 386897
rect 502391 386863 502424 386897
rect 502324 386656 502424 386863
rect 504842 386788 504868 387188
rect 505668 387050 505694 387188
rect 505884 387050 505984 387319
rect 505668 386953 505984 387050
rect 505668 386930 505917 386953
rect 505668 386788 505694 386930
rect 505884 386919 505917 386930
rect 505951 386919 505984 386953
rect 498564 386507 498597 386541
rect 498631 386507 498664 386541
rect 498564 386460 498664 386507
rect 498393 386340 498664 386460
rect 498393 386149 498419 386340
rect 494633 385967 494659 386116
rect 494804 385941 494904 386116
rect 498564 386141 498664 386340
rect 504842 386330 504868 386730
rect 505668 386594 505694 386730
rect 505884 386594 505984 386919
rect 505668 386553 505984 386594
rect 505668 386519 505917 386553
rect 505951 386519 505984 386553
rect 505668 386474 505984 386519
rect 505668 386330 505694 386474
rect 498564 386107 498597 386141
rect 498631 386107 498664 386141
rect 493317 385509 493343 385909
rect 494633 385780 494659 385909
rect 494804 385907 494837 385941
rect 494871 385907 494904 385941
rect 494804 385780 494904 385907
rect 494633 385660 494904 385780
rect 497077 385691 497103 386091
rect 498393 386004 498419 386091
rect 498564 386004 498664 386107
rect 498393 385884 498664 386004
rect 498393 385691 498419 385884
rect 498564 385741 498664 385884
rect 504842 385872 504868 386272
rect 505668 386138 505694 386272
rect 505884 386153 505984 386474
rect 505884 386138 505917 386153
rect 505668 386119 505917 386138
rect 505951 386119 505984 386153
rect 505668 386018 505984 386119
rect 505668 385872 505694 386018
rect 498564 385707 498597 385741
rect 498631 385707 498664 385741
rect 494633 385509 494659 385660
rect 494804 385541 494904 385660
rect 494804 385507 494837 385541
rect 494871 385507 494904 385541
rect 493317 385051 493343 385451
rect 494633 385324 494659 385451
rect 494804 385324 494904 385507
rect 494633 385204 494904 385324
rect 497077 385233 497103 385633
rect 498393 385548 498419 385633
rect 498564 385548 498664 385707
rect 498393 385428 498664 385548
rect 498393 385233 498419 385428
rect 498564 385341 498664 385428
rect 498564 385307 498597 385341
rect 498631 385307 498664 385341
rect 494633 385051 494659 385204
rect 494804 385141 494904 385204
rect 494804 385107 494837 385141
rect 494871 385107 494904 385141
rect 493317 384593 493343 384993
rect 494633 384868 494659 384993
rect 494804 384868 494904 385107
rect 494633 384748 494904 384868
rect 497077 384775 497103 385175
rect 498393 385092 498419 385175
rect 498564 385092 498664 385307
rect 500837 385123 500863 385523
rect 502153 385376 502179 385523
rect 502324 385433 502424 385616
rect 502324 385399 502357 385433
rect 502391 385399 502424 385433
rect 504842 385414 504868 385814
rect 505668 385682 505694 385814
rect 505884 385753 505984 386018
rect 505884 385719 505917 385753
rect 505951 385719 505984 385753
rect 505884 385682 505984 385719
rect 505668 385562 505984 385682
rect 505668 385414 505694 385562
rect 502324 385376 502424 385399
rect 502153 385256 502424 385376
rect 505884 385356 505984 385562
rect 516122 387704 516148 388104
rect 516948 387962 516974 388104
rect 517164 387962 517264 388119
rect 516948 387842 517264 387962
rect 516948 387704 516974 387842
rect 517164 387753 517264 387842
rect 517164 387719 517197 387753
rect 517231 387719 517264 387753
rect 523397 387799 523423 388199
rect 524713 388060 524739 388199
rect 524884 388060 524984 388307
rect 524713 387941 524984 388060
rect 524713 387940 524917 387941
rect 524713 387799 524739 387940
rect 524884 387907 524917 387940
rect 524951 387907 524984 387941
rect 516122 387246 516148 387646
rect 516948 387506 516974 387646
rect 517164 387506 517264 387719
rect 516948 387386 517264 387506
rect 516948 387246 516974 387386
rect 517164 387353 517264 387386
rect 517164 387319 517197 387353
rect 517231 387319 517264 387353
rect 516122 386788 516148 387188
rect 516948 387050 516974 387188
rect 517164 387050 517264 387319
rect 516948 386953 517264 387050
rect 516948 386930 517197 386953
rect 516948 386788 516974 386930
rect 517164 386919 517197 386930
rect 517231 386919 517264 386953
rect 516122 386330 516148 386730
rect 516948 386594 516974 386730
rect 517164 386594 517264 386919
rect 516948 386553 517264 386594
rect 516948 386519 517197 386553
rect 517231 386519 517264 386553
rect 516948 386474 517264 386519
rect 516948 386330 516974 386474
rect 516122 385872 516148 386272
rect 516948 386138 516974 386272
rect 517164 386153 517264 386474
rect 517164 386138 517197 386153
rect 516948 386119 517197 386138
rect 517231 386119 517264 386153
rect 516948 386018 517264 386119
rect 516948 385872 516974 386018
rect 516122 385414 516148 385814
rect 516948 385682 516974 385814
rect 517164 385753 517264 386018
rect 517164 385719 517197 385753
rect 517231 385719 517264 385753
rect 517164 385682 517264 385719
rect 516948 385562 517264 385682
rect 516948 385414 516974 385562
rect 517164 385356 517264 385562
rect 523397 387341 523423 387741
rect 524713 387604 524739 387741
rect 524884 387604 524984 387907
rect 524713 387541 524984 387604
rect 524713 387507 524917 387541
rect 524951 387507 524984 387541
rect 524713 387484 524984 387507
rect 524713 387341 524739 387484
rect 523397 386883 523423 387283
rect 524713 387148 524739 387283
rect 524884 387148 524984 387484
rect 524713 387141 524984 387148
rect 524713 387107 524917 387141
rect 524951 387107 524984 387141
rect 524713 387028 524984 387107
rect 524713 386883 524739 387028
rect 523397 386425 523423 386825
rect 524713 386692 524739 386825
rect 524884 386741 524984 387028
rect 524884 386707 524917 386741
rect 524951 386707 524984 386741
rect 524884 386692 524984 386707
rect 524713 386572 524984 386692
rect 524713 386425 524739 386572
rect 523397 385967 523423 386367
rect 524713 386236 524739 386367
rect 524884 386341 524984 386572
rect 524884 386307 524917 386341
rect 524951 386307 524984 386341
rect 524884 386236 524984 386307
rect 524713 386116 524984 386236
rect 524713 385967 524739 386116
rect 524884 385941 524984 386116
rect 523397 385509 523423 385909
rect 524713 385780 524739 385909
rect 524884 385907 524917 385941
rect 524951 385907 524984 385941
rect 524884 385780 524984 385907
rect 524713 385660 524984 385780
rect 524713 385509 524739 385660
rect 524884 385541 524984 385660
rect 524884 385507 524917 385541
rect 524951 385507 524984 385541
rect 502153 385123 502179 385256
rect 498393 384972 498664 385092
rect 498393 384775 498419 384972
rect 498564 384941 498664 384972
rect 498564 384907 498597 384941
rect 498631 384907 498664 384941
rect 494633 384593 494659 384748
rect 494804 384741 494904 384748
rect 494804 384707 494837 384741
rect 494871 384707 494904 384741
rect 493317 384135 493343 384535
rect 494633 384412 494659 384535
rect 494804 384412 494904 384707
rect 494633 384341 494904 384412
rect 494633 384307 494837 384341
rect 494871 384307 494904 384341
rect 497077 384317 497103 384717
rect 498393 384636 498419 384717
rect 498564 384636 498664 384907
rect 500837 384665 500863 385065
rect 502153 384920 502179 385065
rect 502324 385033 502424 385256
rect 523397 385051 523423 385451
rect 524713 385324 524739 385451
rect 524884 385324 524984 385507
rect 524713 385204 524984 385324
rect 524713 385051 524739 385204
rect 524884 385141 524984 385204
rect 524884 385107 524917 385141
rect 524951 385107 524984 385141
rect 502324 384999 502357 385033
rect 502391 384999 502424 385033
rect 502324 384920 502424 384999
rect 502153 384800 502424 384920
rect 502153 384665 502179 384800
rect 498393 384541 498664 384636
rect 498393 384516 498597 384541
rect 498393 384317 498419 384516
rect 498564 384507 498597 384516
rect 498631 384507 498664 384541
rect 494633 384292 494904 384307
rect 494633 384135 494659 384292
rect 493317 383677 493343 384077
rect 494633 383956 494659 384077
rect 494804 383956 494904 384292
rect 494633 383941 494904 383956
rect 494633 383907 494837 383941
rect 494871 383907 494904 383941
rect 494633 383836 494904 383907
rect 497077 383859 497103 384259
rect 498393 384180 498419 384259
rect 498564 384180 498664 384507
rect 502324 384633 502424 384800
rect 500837 384207 500863 384607
rect 502153 384464 502179 384607
rect 502324 384599 502357 384633
rect 502391 384599 502424 384633
rect 502324 384464 502424 384599
rect 502153 384344 502424 384464
rect 502153 384207 502179 384344
rect 502324 384233 502424 384344
rect 498393 384141 498664 384180
rect 502324 384199 502357 384233
rect 502391 384199 502424 384233
rect 498393 384107 498597 384141
rect 498631 384107 498664 384141
rect 498393 384060 498664 384107
rect 498393 383859 498419 384060
rect 494633 383677 494659 383836
rect 493317 383219 493343 383619
rect 494633 383500 494659 383619
rect 494804 383541 494904 383836
rect 494804 383507 494837 383541
rect 494871 383507 494904 383541
rect 494804 383500 494904 383507
rect 494633 383380 494904 383500
rect 497077 383401 497103 383801
rect 498393 383724 498419 383801
rect 498564 383741 498664 384060
rect 500837 383749 500863 384149
rect 502153 384008 502179 384149
rect 502324 384008 502424 384199
rect 502153 383888 502424 384008
rect 502153 383749 502179 383888
rect 502324 383833 502424 383888
rect 502324 383799 502357 383833
rect 502391 383799 502424 383833
rect 498564 383724 498597 383741
rect 498393 383707 498597 383724
rect 498631 383707 498664 383741
rect 498393 383604 498664 383707
rect 498393 383401 498419 383604
rect 494633 383219 494659 383380
rect 493317 382761 493343 383161
rect 494633 383044 494659 383161
rect 494804 383141 494904 383380
rect 494804 383107 494837 383141
rect 494871 383107 494904 383141
rect 494804 383044 494904 383107
rect 494633 382924 494904 383044
rect 497077 382943 497103 383343
rect 498393 383268 498419 383343
rect 498564 383341 498664 383604
rect 498564 383307 498597 383341
rect 498631 383307 498664 383341
rect 498564 383268 498664 383307
rect 498393 383148 498664 383268
rect 500837 383291 500863 383691
rect 502153 383552 502179 383691
rect 502324 383552 502424 383799
rect 502153 383433 502424 383552
rect 502153 383432 502357 383433
rect 502153 383291 502179 383432
rect 502324 383399 502357 383432
rect 502391 383399 502424 383433
rect 498393 382943 498419 383148
rect 494633 382761 494659 382924
rect 494804 382741 494904 382924
rect 498564 382941 498664 383148
rect 498564 382907 498597 382941
rect 498631 382907 498664 382941
rect 494804 382707 494837 382741
rect 494871 382707 494904 382741
rect 493317 382303 493343 382703
rect 494633 382588 494659 382703
rect 494804 382588 494904 382707
rect 494633 382468 494904 382588
rect 497077 382485 497103 382885
rect 498393 382812 498419 382885
rect 498564 382812 498664 382907
rect 500837 382833 500863 383233
rect 502153 383096 502179 383233
rect 502324 383096 502424 383399
rect 502153 383033 502424 383096
rect 502153 382999 502357 383033
rect 502391 382999 502424 383033
rect 502153 382976 502424 382999
rect 502153 382833 502179 382976
rect 498393 382692 498664 382812
rect 498393 382485 498419 382692
rect 498564 382541 498664 382692
rect 498564 382507 498597 382541
rect 498631 382507 498664 382541
rect 494633 382303 494659 382468
rect 494804 382341 494904 382468
rect 494804 382307 494837 382341
rect 494871 382307 494904 382341
rect 493317 381845 493343 382245
rect 494633 382132 494659 382245
rect 494804 382132 494904 382307
rect 494633 382012 494904 382132
rect 497077 382027 497103 382427
rect 498393 382356 498419 382427
rect 498564 382356 498664 382507
rect 500837 382375 500863 382775
rect 502153 382640 502179 382775
rect 502324 382640 502424 382976
rect 502153 382633 502424 382640
rect 502153 382599 502357 382633
rect 502391 382599 502424 382633
rect 502153 382520 502424 382599
rect 523397 384593 523423 384993
rect 524713 384868 524739 384993
rect 524884 384868 524984 385107
rect 524713 384748 524984 384868
rect 524713 384593 524739 384748
rect 524884 384741 524984 384748
rect 524884 384707 524917 384741
rect 524951 384707 524984 384741
rect 523397 384135 523423 384535
rect 524713 384412 524739 384535
rect 524884 384412 524984 384707
rect 524713 384341 524984 384412
rect 524713 384307 524917 384341
rect 524951 384307 524984 384341
rect 524713 384292 524984 384307
rect 524713 384135 524739 384292
rect 523397 383677 523423 384077
rect 524713 383956 524739 384077
rect 524884 383956 524984 384292
rect 524713 383941 524984 383956
rect 524713 383907 524917 383941
rect 524951 383907 524984 383941
rect 524713 383836 524984 383907
rect 524713 383677 524739 383836
rect 523397 383219 523423 383619
rect 524713 383500 524739 383619
rect 524884 383541 524984 383836
rect 524884 383507 524917 383541
rect 524951 383507 524984 383541
rect 524884 383500 524984 383507
rect 524713 383380 524984 383500
rect 524713 383219 524739 383380
rect 523397 382761 523423 383161
rect 524713 383044 524739 383161
rect 524884 383141 524984 383380
rect 524884 383107 524917 383141
rect 524951 383107 524984 383141
rect 524884 383044 524984 383107
rect 524713 382924 524984 383044
rect 524713 382761 524739 382924
rect 524884 382741 524984 382924
rect 524884 382707 524917 382741
rect 524951 382707 524984 382741
rect 502153 382375 502179 382520
rect 498393 382236 498664 382356
rect 498393 382027 498419 382236
rect 498564 382141 498664 382236
rect 498564 382107 498597 382141
rect 498631 382107 498664 382141
rect 494633 381845 494659 382012
rect 494804 381941 494904 382012
rect 494804 381907 494837 381941
rect 494871 381907 494904 381941
rect 493317 381387 493343 381787
rect 494633 381676 494659 381787
rect 494804 381676 494904 381907
rect 494633 381556 494904 381676
rect 497077 381569 497103 381969
rect 498393 381900 498419 381969
rect 498564 381900 498664 382107
rect 498393 381780 498664 381900
rect 500837 381917 500863 382317
rect 502153 382184 502179 382317
rect 502324 382233 502424 382520
rect 523397 382303 523423 382703
rect 524713 382588 524739 382703
rect 524884 382588 524984 382707
rect 524713 382468 524984 382588
rect 524713 382303 524739 382468
rect 524884 382341 524984 382468
rect 524884 382307 524917 382341
rect 524951 382307 524984 382341
rect 502324 382199 502357 382233
rect 502391 382199 502424 382233
rect 502324 382184 502424 382199
rect 502153 382064 502424 382184
rect 502153 381917 502179 382064
rect 498393 381569 498419 381780
rect 498564 381741 498664 381780
rect 498564 381707 498597 381741
rect 498631 381707 498664 381741
rect 494633 381387 494659 381556
rect 494804 381541 494904 381556
rect 494804 381507 494837 381541
rect 494871 381507 494904 381541
rect 493317 380929 493343 381329
rect 494633 381220 494659 381329
rect 494804 381220 494904 381507
rect 494633 381141 494904 381220
rect 494633 381107 494837 381141
rect 494871 381107 494904 381141
rect 497077 381111 497103 381511
rect 498393 381444 498419 381511
rect 498564 381444 498664 381707
rect 500837 381459 500863 381859
rect 502153 381728 502179 381859
rect 502324 381833 502424 382064
rect 523397 381845 523423 382245
rect 524713 382132 524739 382245
rect 524884 382132 524984 382307
rect 524713 382012 524984 382132
rect 524713 381845 524739 382012
rect 524884 381941 524984 382012
rect 524884 381907 524917 381941
rect 524951 381907 524984 381941
rect 502324 381799 502357 381833
rect 502391 381799 502424 381833
rect 502324 381728 502424 381799
rect 502153 381608 502424 381728
rect 502153 381459 502179 381608
rect 498393 381341 498664 381444
rect 502324 381433 502424 381608
rect 498393 381324 498597 381341
rect 498393 381111 498419 381324
rect 498564 381307 498597 381324
rect 498631 381307 498664 381341
rect 494633 381100 494904 381107
rect 494633 380929 494659 381100
rect 493317 380471 493343 380871
rect 494633 380764 494659 380871
rect 494804 380764 494904 381100
rect 494633 380741 494904 380764
rect 494633 380707 494837 380741
rect 494871 380707 494904 380741
rect 494633 380644 494904 380707
rect 494633 380471 494659 380644
rect 493317 380013 493343 380413
rect 494633 380308 494659 380413
rect 494804 380341 494904 380644
rect 497077 380653 497103 381053
rect 498393 380988 498419 381053
rect 498564 380988 498664 381307
rect 500837 381001 500863 381401
rect 502153 381272 502179 381401
rect 502324 381399 502357 381433
rect 502391 381399 502424 381433
rect 502324 381272 502424 381399
rect 502153 381152 502424 381272
rect 502153 381001 502179 381152
rect 502324 381033 502424 381152
rect 498393 380941 498664 380988
rect 502324 380999 502357 381033
rect 502391 380999 502424 381033
rect 498393 380907 498597 380941
rect 498631 380907 498664 380941
rect 498393 380868 498664 380907
rect 498393 380653 498419 380868
rect 494804 380308 494837 380341
rect 494633 380307 494837 380308
rect 494871 380307 494904 380341
rect 494633 380188 494904 380307
rect 497077 380195 497103 380595
rect 498393 380532 498419 380595
rect 498564 380541 498664 380868
rect 500837 380543 500863 380943
rect 502153 380816 502179 380943
rect 502324 380816 502424 380999
rect 502153 380696 502424 380816
rect 502153 380543 502179 380696
rect 502324 380633 502424 380696
rect 502324 380599 502357 380633
rect 502391 380599 502424 380633
rect 498564 380532 498597 380541
rect 498393 380507 498597 380532
rect 498631 380507 498664 380541
rect 498393 380412 498664 380507
rect 498393 380195 498419 380412
rect 494633 380013 494659 380188
rect 493317 379555 493343 379955
rect 494633 379852 494659 379955
rect 494804 379941 494904 380188
rect 498564 380141 498664 380412
rect 494804 379907 494837 379941
rect 494871 379907 494904 379941
rect 494804 379852 494904 379907
rect 494633 379732 494904 379852
rect 497077 379737 497103 380137
rect 498393 380076 498419 380137
rect 498564 380107 498597 380141
rect 498631 380107 498664 380141
rect 498564 380076 498664 380107
rect 500837 380085 500863 380485
rect 502153 380360 502179 380485
rect 502324 380360 502424 380599
rect 502153 380240 502424 380360
rect 502153 380085 502179 380240
rect 502324 380233 502424 380240
rect 502324 380199 502357 380233
rect 502391 380199 502424 380233
rect 498393 379956 498664 380076
rect 502324 379992 502424 380199
rect 498393 379737 498419 379956
rect 498564 379741 498664 379956
rect 494633 379555 494659 379732
rect 494804 379541 494904 379732
rect 498564 379707 498597 379741
rect 498631 379707 498664 379741
rect 494804 379507 494837 379541
rect 494871 379507 494904 379541
rect 493317 379097 493343 379497
rect 494633 379396 494659 379497
rect 494804 379396 494904 379507
rect 494633 379276 494904 379396
rect 497077 379279 497103 379679
rect 498393 379620 498419 379679
rect 498564 379620 498664 379707
rect 498393 379500 498664 379620
rect 498393 379279 498419 379500
rect 498564 379341 498664 379500
rect 498564 379307 498597 379341
rect 498631 379307 498664 379341
rect 523397 381387 523423 381787
rect 524713 381676 524739 381787
rect 524884 381676 524984 381907
rect 524713 381556 524984 381676
rect 524713 381387 524739 381556
rect 524884 381541 524984 381556
rect 524884 381507 524917 381541
rect 524951 381507 524984 381541
rect 523397 380929 523423 381329
rect 524713 381220 524739 381329
rect 524884 381220 524984 381507
rect 524713 381141 524984 381220
rect 524713 381107 524917 381141
rect 524951 381107 524984 381141
rect 524713 381100 524984 381107
rect 524713 380929 524739 381100
rect 523397 380471 523423 380871
rect 524713 380764 524739 380871
rect 524884 380764 524984 381100
rect 524713 380741 524984 380764
rect 524713 380707 524917 380741
rect 524951 380707 524984 380741
rect 524713 380644 524984 380707
rect 524713 380471 524739 380644
rect 523397 380013 523423 380413
rect 524713 380308 524739 380413
rect 524884 380341 524984 380644
rect 524884 380308 524917 380341
rect 524713 380307 524917 380308
rect 524951 380307 524984 380341
rect 524713 380188 524984 380307
rect 524713 380013 524739 380188
rect 523397 379555 523423 379955
rect 524713 379852 524739 379955
rect 524884 379941 524984 380188
rect 524884 379907 524917 379941
rect 524951 379907 524984 379941
rect 524884 379852 524984 379907
rect 524713 379732 524984 379852
rect 524713 379555 524739 379732
rect 524884 379541 524984 379732
rect 524884 379507 524917 379541
rect 524951 379507 524984 379541
rect 494633 379097 494659 379276
rect 494804 379141 494904 379276
rect 494804 379107 494837 379141
rect 494871 379107 494904 379141
rect 493317 378639 493343 379039
rect 494633 378940 494659 379039
rect 494804 378940 494904 379107
rect 494633 378820 494904 378940
rect 497077 378821 497103 379221
rect 498393 379164 498419 379221
rect 498564 379164 498664 379307
rect 498393 379044 498664 379164
rect 523397 379097 523423 379497
rect 524713 379396 524739 379497
rect 524884 379396 524984 379507
rect 524713 379276 524984 379396
rect 524713 379097 524739 379276
rect 524884 379141 524984 379276
rect 524884 379107 524917 379141
rect 524951 379107 524984 379141
rect 498393 378821 498419 379044
rect 498564 378941 498664 379044
rect 498564 378907 498597 378941
rect 498631 378907 498664 378941
rect 494633 378639 494659 378820
rect 494804 378741 494904 378820
rect 494804 378707 494837 378741
rect 494871 378707 494904 378741
rect 493317 378181 493343 378581
rect 494633 378484 494659 378581
rect 494804 378484 494904 378707
rect 494633 378364 494904 378484
rect 494633 378181 494659 378364
rect 494804 378341 494904 378364
rect 497077 378363 497103 378763
rect 498393 378708 498419 378763
rect 498564 378708 498664 378907
rect 498393 378588 498664 378708
rect 523397 378639 523423 379039
rect 524713 378940 524739 379039
rect 524884 378940 524984 379107
rect 524713 378820 524984 378940
rect 524713 378639 524739 378820
rect 524884 378741 524984 378820
rect 524884 378707 524917 378741
rect 524951 378707 524984 378741
rect 498393 378363 498419 378588
rect 498564 378541 498664 378588
rect 498564 378507 498597 378541
rect 498631 378507 498664 378541
rect 494804 378307 494837 378341
rect 494871 378307 494904 378341
rect 493317 377723 493343 378123
rect 494633 378028 494659 378123
rect 494804 378028 494904 378307
rect 494633 377941 494904 378028
rect 494633 377908 494837 377941
rect 494633 377723 494659 377908
rect 494804 377907 494837 377908
rect 494871 377907 494904 377941
rect 493317 377265 493343 377665
rect 494633 377572 494659 377665
rect 494804 377572 494904 377907
rect 497077 377905 497103 378305
rect 498393 378252 498419 378305
rect 498564 378252 498664 378507
rect 498393 378141 498664 378252
rect 523397 378181 523423 378581
rect 524713 378484 524739 378581
rect 524884 378484 524984 378707
rect 524713 378364 524984 378484
rect 524713 378181 524739 378364
rect 524884 378341 524984 378364
rect 524884 378307 524917 378341
rect 524951 378307 524984 378341
rect 498393 378132 498597 378141
rect 498393 377905 498419 378132
rect 498564 378107 498597 378132
rect 498631 378107 498664 378141
rect 494633 377541 494904 377572
rect 494633 377507 494837 377541
rect 494871 377507 494904 377541
rect 494633 377452 494904 377507
rect 494633 377265 494659 377452
rect 493317 376807 493343 377207
rect 494633 377116 494659 377207
rect 494804 377141 494904 377452
rect 497077 377447 497103 377847
rect 498393 377796 498419 377847
rect 498564 377796 498664 378107
rect 498393 377741 498664 377796
rect 498393 377707 498597 377741
rect 498631 377707 498664 377741
rect 498393 377676 498664 377707
rect 523397 377723 523423 378123
rect 524713 378028 524739 378123
rect 524884 378028 524984 378307
rect 524713 377941 524984 378028
rect 524713 377908 524917 377941
rect 524713 377723 524739 377908
rect 524884 377907 524917 377908
rect 524951 377907 524984 377941
rect 498393 377447 498419 377676
rect 494804 377116 494837 377141
rect 494633 377107 494837 377116
rect 494871 377107 494904 377141
rect 494633 376996 494904 377107
rect 494633 376807 494659 376996
rect 493317 376349 493343 376749
rect 494633 376660 494659 376749
rect 494804 376741 494904 376996
rect 497077 376989 497103 377389
rect 498393 377340 498419 377389
rect 498564 377341 498664 377676
rect 498564 377340 498597 377341
rect 498393 377307 498597 377340
rect 498631 377307 498664 377341
rect 498393 377220 498664 377307
rect 501082 377220 501108 377620
rect 501908 377472 501934 377620
rect 502124 377495 502224 377598
rect 502124 377472 502157 377495
rect 501908 377461 502157 377472
rect 502191 377461 502224 377495
rect 501908 377352 502224 377461
rect 501908 377220 501934 377352
rect 498393 376989 498419 377220
rect 498564 376941 498664 377220
rect 494804 376707 494837 376741
rect 494871 376707 494904 376741
rect 494804 376660 494904 376707
rect 494633 376540 494904 376660
rect 494633 376349 494659 376540
rect 494804 376341 494904 376540
rect 497077 376531 497103 376931
rect 498393 376884 498419 376931
rect 498564 376907 498597 376941
rect 498631 376907 498664 376941
rect 498564 376884 498664 376907
rect 498393 376764 498664 376884
rect 498393 376531 498419 376764
rect 498564 376541 498664 376764
rect 501082 376762 501108 377162
rect 501908 377016 501934 377162
rect 502124 377095 502224 377352
rect 502124 377061 502157 377095
rect 502191 377061 502224 377095
rect 502124 377016 502224 377061
rect 501908 376896 502224 377016
rect 504597 376989 504623 377389
rect 505913 377242 505939 377389
rect 506084 377299 506184 377482
rect 506084 377265 506117 377299
rect 506151 377265 506184 377299
rect 506084 377242 506184 377265
rect 505913 377122 506184 377242
rect 505913 376989 505939 377122
rect 501908 376762 501934 376896
rect 498564 376507 498597 376541
rect 498631 376507 498664 376541
rect 494804 376307 494837 376341
rect 494871 376307 494904 376341
rect 493317 375891 493343 376291
rect 494633 376204 494659 376291
rect 494804 376204 494904 376307
rect 494633 376084 494904 376204
rect 494633 375891 494659 376084
rect 494804 375941 494904 376084
rect 497077 376073 497103 376473
rect 498393 376428 498419 376473
rect 498564 376428 498664 376507
rect 498393 376308 498664 376428
rect 498393 376073 498419 376308
rect 498564 376141 498664 376308
rect 501082 376304 501108 376704
rect 501908 376560 501934 376704
rect 502124 376695 502224 376896
rect 502124 376661 502157 376695
rect 502191 376661 502224 376695
rect 502124 376560 502224 376661
rect 501908 376440 502224 376560
rect 504597 376531 504623 376931
rect 505913 376786 505939 376931
rect 506084 376899 506184 377122
rect 512117 376989 512143 377389
rect 513433 377242 513459 377389
rect 513604 377299 513704 377482
rect 513604 377265 513637 377299
rect 513671 377265 513704 377299
rect 513604 377242 513704 377265
rect 513433 377122 513704 377242
rect 513433 376989 513459 377122
rect 506084 376865 506117 376899
rect 506151 376865 506184 376899
rect 506084 376786 506184 376865
rect 505913 376666 506184 376786
rect 505913 376531 505939 376666
rect 501908 376304 501934 376440
rect 502124 376295 502224 376440
rect 506084 376499 506184 376666
rect 512117 376531 512143 376931
rect 513433 376786 513459 376931
rect 513604 376899 513704 377122
rect 513604 376865 513637 376899
rect 513671 376865 513704 376899
rect 513604 376786 513704 376865
rect 513433 376666 513704 376786
rect 513433 376531 513459 376666
rect 502124 376261 502157 376295
rect 502191 376261 502224 376295
rect 498564 376107 498597 376141
rect 498631 376107 498664 376141
rect 494804 375907 494837 375941
rect 494871 375907 494904 375941
rect 493317 375433 493343 375833
rect 494633 375748 494659 375833
rect 494804 375748 494904 375907
rect 494633 375628 494904 375748
rect 494633 375433 494659 375628
rect 494804 375541 494904 375628
rect 497077 375615 497103 376015
rect 498393 375972 498419 376015
rect 498564 375972 498664 376107
rect 498393 375852 498664 375972
rect 498393 375615 498419 375852
rect 498564 375741 498664 375852
rect 501082 375846 501108 376246
rect 501908 376104 501934 376246
rect 502124 376104 502224 376261
rect 501908 375984 502224 376104
rect 504597 376073 504623 376473
rect 505913 376330 505939 376473
rect 506084 376465 506117 376499
rect 506151 376465 506184 376499
rect 506084 376330 506184 376465
rect 513604 376499 513704 376666
rect 505913 376210 506184 376330
rect 505913 376073 505939 376210
rect 506084 376099 506184 376210
rect 506084 376065 506117 376099
rect 506151 376065 506184 376099
rect 512117 376073 512143 376473
rect 513433 376330 513459 376473
rect 513604 376465 513637 376499
rect 513671 376465 513704 376499
rect 513604 376330 513704 376465
rect 513433 376210 513704 376330
rect 513433 376073 513459 376210
rect 513604 376099 513704 376210
rect 501908 375846 501934 375984
rect 502124 375895 502224 375984
rect 502124 375861 502157 375895
rect 502191 375861 502224 375895
rect 498564 375707 498597 375741
rect 498631 375707 498664 375741
rect 494804 375507 494837 375541
rect 494871 375507 494904 375541
rect 493317 374975 493343 375375
rect 494633 375292 494659 375375
rect 494804 375292 494904 375507
rect 494633 375172 494904 375292
rect 494633 374975 494659 375172
rect 494804 375141 494904 375172
rect 497077 375157 497103 375557
rect 498393 375516 498419 375557
rect 498564 375516 498664 375707
rect 498393 375396 498664 375516
rect 498393 375157 498419 375396
rect 498564 375341 498664 375396
rect 501082 375388 501108 375788
rect 501908 375648 501934 375788
rect 502124 375648 502224 375861
rect 501908 375528 502224 375648
rect 504597 375615 504623 376015
rect 505913 375874 505939 376015
rect 506084 375874 506184 376065
rect 513604 376065 513637 376099
rect 513671 376065 513704 376099
rect 505913 375754 506184 375874
rect 505913 375615 505939 375754
rect 506084 375699 506184 375754
rect 506084 375665 506117 375699
rect 506151 375665 506184 375699
rect 501908 375388 501934 375528
rect 502124 375495 502224 375528
rect 502124 375461 502157 375495
rect 502191 375461 502224 375495
rect 498564 375307 498597 375341
rect 498631 375307 498664 375341
rect 494804 375107 494837 375141
rect 494871 375107 494904 375141
rect 493317 374517 493343 374917
rect 494633 374836 494659 374917
rect 494804 374836 494904 375107
rect 494633 374741 494904 374836
rect 494633 374716 494837 374741
rect 494633 374517 494659 374716
rect 494804 374707 494837 374716
rect 494871 374707 494904 374741
rect 493317 374059 493343 374459
rect 494633 374380 494659 374459
rect 494804 374380 494904 374707
rect 497077 374699 497103 375099
rect 498393 375060 498419 375099
rect 498564 375060 498664 375307
rect 498393 374941 498664 375060
rect 498393 374940 498597 374941
rect 498393 374699 498419 374940
rect 498564 374907 498597 374940
rect 498631 374907 498664 374941
rect 501082 374930 501108 375330
rect 501908 375192 501934 375330
rect 502124 375192 502224 375461
rect 501908 375095 502224 375192
rect 504597 375157 504623 375557
rect 505913 375418 505939 375557
rect 506084 375418 506184 375665
rect 512117 375615 512143 376015
rect 513433 375874 513459 376015
rect 513604 375874 513704 376065
rect 513433 375754 513704 375874
rect 513433 375615 513459 375754
rect 513604 375699 513704 375754
rect 513604 375665 513637 375699
rect 513671 375665 513704 375699
rect 505913 375299 506184 375418
rect 505913 375298 506117 375299
rect 505913 375157 505939 375298
rect 506084 375265 506117 375298
rect 506151 375265 506184 375299
rect 501908 375072 502157 375095
rect 501908 374930 501934 375072
rect 502124 375061 502157 375072
rect 502191 375061 502224 375095
rect 494633 374341 494904 374380
rect 494633 374307 494837 374341
rect 494871 374307 494904 374341
rect 494633 374260 494904 374307
rect 494633 374059 494659 374260
rect 493317 373601 493343 374001
rect 494633 373924 494659 374001
rect 494804 373941 494904 374260
rect 497077 374241 497103 374641
rect 498393 374604 498419 374641
rect 498564 374604 498664 374907
rect 498393 374541 498664 374604
rect 498393 374507 498597 374541
rect 498631 374507 498664 374541
rect 498393 374484 498664 374507
rect 498393 374241 498419 374484
rect 494804 373924 494837 373941
rect 494633 373907 494837 373924
rect 494871 373907 494904 373941
rect 494633 373804 494904 373907
rect 494633 373601 494659 373804
rect 493317 373143 493343 373543
rect 494633 373468 494659 373543
rect 494804 373541 494904 373804
rect 497077 373783 497103 374183
rect 498393 374148 498419 374183
rect 498564 374148 498664 374484
rect 501082 374472 501108 374872
rect 501908 374736 501934 374872
rect 502124 374736 502224 375061
rect 501908 374695 502224 374736
rect 504597 374699 504623 375099
rect 505913 374962 505939 375099
rect 506084 374962 506184 375265
rect 512117 375157 512143 375557
rect 513433 375418 513459 375557
rect 513604 375418 513704 375665
rect 513433 375299 513704 375418
rect 513433 375298 513637 375299
rect 513433 375157 513459 375298
rect 513604 375265 513637 375298
rect 513671 375265 513704 375299
rect 505913 374899 506184 374962
rect 505913 374865 506117 374899
rect 506151 374865 506184 374899
rect 505913 374842 506184 374865
rect 505913 374699 505939 374842
rect 501908 374661 502157 374695
rect 502191 374661 502224 374695
rect 501908 374616 502224 374661
rect 501908 374472 501934 374616
rect 498393 374141 498664 374148
rect 498393 374107 498597 374141
rect 498631 374107 498664 374141
rect 498393 374028 498664 374107
rect 498393 373783 498419 374028
rect 498564 373741 498664 374028
rect 501082 374014 501108 374414
rect 501908 374280 501934 374414
rect 502124 374295 502224 374616
rect 506084 374606 506184 374842
rect 512117 374699 512143 375099
rect 513433 374962 513459 375099
rect 513604 374962 513704 375265
rect 523397 377265 523423 377665
rect 524713 377572 524739 377665
rect 524884 377572 524984 377907
rect 524713 377541 524984 377572
rect 524713 377507 524917 377541
rect 524951 377507 524984 377541
rect 524713 377452 524984 377507
rect 524713 377265 524739 377452
rect 523397 376807 523423 377207
rect 524713 377116 524739 377207
rect 524884 377141 524984 377452
rect 524884 377116 524917 377141
rect 524713 377107 524917 377116
rect 524951 377107 524984 377141
rect 524713 376996 524984 377107
rect 524713 376807 524739 376996
rect 523397 376349 523423 376749
rect 524713 376660 524739 376749
rect 524884 376741 524984 376996
rect 524884 376707 524917 376741
rect 524951 376707 524984 376741
rect 524884 376660 524984 376707
rect 524713 376540 524984 376660
rect 524713 376349 524739 376540
rect 524884 376341 524984 376540
rect 524884 376307 524917 376341
rect 524951 376307 524984 376341
rect 523397 375891 523423 376291
rect 524713 376204 524739 376291
rect 524884 376204 524984 376307
rect 524713 376084 524984 376204
rect 524713 375891 524739 376084
rect 524884 375941 524984 376084
rect 524884 375907 524917 375941
rect 524951 375907 524984 375941
rect 523397 375433 523423 375833
rect 524713 375748 524739 375833
rect 524884 375748 524984 375907
rect 524713 375628 524984 375748
rect 524713 375433 524739 375628
rect 524884 375541 524984 375628
rect 524884 375507 524917 375541
rect 524951 375507 524984 375541
rect 523397 374975 523423 375375
rect 524713 375292 524739 375375
rect 524884 375292 524984 375507
rect 524713 375172 524984 375292
rect 524713 374975 524739 375172
rect 524884 375141 524984 375172
rect 524884 375107 524917 375141
rect 524951 375107 524984 375141
rect 513433 374899 513704 374962
rect 513433 374865 513637 374899
rect 513671 374865 513704 374899
rect 513433 374842 513704 374865
rect 513433 374699 513459 374842
rect 513604 374606 513704 374842
rect 502124 374280 502157 374295
rect 501908 374261 502157 374280
rect 502191 374261 502224 374295
rect 501908 374160 502224 374261
rect 501908 374014 501934 374160
rect 494804 373507 494837 373541
rect 494871 373507 494904 373541
rect 494804 373468 494904 373507
rect 494633 373348 494904 373468
rect 494633 373143 494659 373348
rect 494804 373141 494904 373348
rect 497077 373325 497103 373725
rect 498393 373692 498419 373725
rect 498564 373707 498597 373741
rect 498631 373707 498664 373741
rect 498564 373692 498664 373707
rect 498393 373572 498664 373692
rect 498393 373325 498419 373572
rect 498564 373341 498664 373572
rect 501082 373556 501108 373956
rect 501908 373824 501934 373956
rect 502124 373895 502224 374160
rect 502124 373861 502157 373895
rect 502191 373861 502224 373895
rect 502124 373824 502224 373861
rect 501908 373704 502224 373824
rect 501908 373556 501934 373704
rect 502124 373498 502224 373704
rect 498564 373307 498597 373341
rect 498631 373307 498664 373341
rect 494804 373107 494837 373141
rect 494871 373107 494904 373141
rect 493317 372685 493343 373085
rect 494633 373012 494659 373085
rect 494804 373012 494904 373107
rect 494633 372892 494904 373012
rect 494633 372685 494659 372892
rect 494804 372741 494904 372892
rect 497077 372867 497103 373267
rect 498393 373236 498419 373267
rect 498564 373236 498664 373307
rect 498393 373116 498664 373236
rect 498393 372867 498419 373116
rect 498564 372941 498664 373116
rect 498564 372907 498597 372941
rect 498631 372907 498664 372941
rect 494804 372707 494837 372741
rect 494871 372707 494904 372741
rect 493317 372227 493343 372627
rect 494633 372556 494659 372627
rect 494804 372556 494904 372707
rect 494633 372436 494904 372556
rect 494633 372227 494659 372436
rect 494804 372341 494904 372436
rect 497077 372409 497103 372809
rect 498393 372780 498419 372809
rect 498564 372780 498664 372907
rect 498393 372660 498664 372780
rect 498393 372409 498419 372660
rect 498564 372541 498664 372660
rect 498564 372507 498597 372541
rect 498631 372507 498664 372541
rect 494804 372307 494837 372341
rect 494871 372307 494904 372341
rect 498564 372316 498664 372507
rect 493317 371769 493343 372169
rect 494633 372100 494659 372169
rect 494804 372100 494904 372307
rect 494633 371980 494904 372100
rect 494633 371769 494659 371980
rect 494804 371941 494904 371980
rect 494804 371907 494837 371941
rect 494871 371907 494904 371941
rect 493317 371311 493343 371711
rect 494633 371644 494659 371711
rect 494804 371644 494904 371907
rect 494633 371541 494904 371644
rect 494633 371524 494837 371541
rect 494633 371311 494659 371524
rect 494804 371507 494837 371524
rect 494871 371507 494904 371541
rect 493317 370853 493343 371253
rect 494633 371188 494659 371253
rect 494804 371188 494904 371507
rect 494633 371141 494904 371188
rect 494633 371107 494837 371141
rect 494871 371107 494904 371141
rect 494633 371068 494904 371107
rect 494633 370853 494659 371068
rect 493317 370395 493343 370795
rect 494633 370732 494659 370795
rect 494804 370741 494904 371068
rect 494804 370732 494837 370741
rect 494633 370707 494837 370732
rect 494871 370707 494904 370741
rect 494633 370612 494904 370707
rect 494633 370395 494659 370612
rect 494804 370341 494904 370612
rect 493317 369937 493343 370337
rect 494633 370276 494659 370337
rect 494804 370307 494837 370341
rect 494871 370307 494904 370341
rect 494804 370276 494904 370307
rect 494633 370156 494904 370276
rect 494633 369937 494659 370156
rect 494804 369941 494904 370156
rect 494804 369907 494837 369941
rect 494871 369907 494904 369941
rect 493317 369479 493343 369879
rect 494633 369820 494659 369879
rect 494804 369820 494904 369907
rect 494633 369700 494904 369820
rect 494633 369479 494659 369700
rect 494804 369541 494904 369700
rect 494804 369507 494837 369541
rect 494871 369507 494904 369541
rect 493317 369021 493343 369421
rect 494633 369364 494659 369421
rect 494804 369364 494904 369507
rect 494633 369244 494904 369364
rect 494633 369021 494659 369244
rect 494804 369141 494904 369244
rect 494804 369107 494837 369141
rect 494871 369107 494904 369141
rect 493317 368563 493343 368963
rect 494633 368908 494659 368963
rect 494804 368908 494904 369107
rect 494633 368788 494904 368908
rect 494633 368563 494659 368788
rect 494804 368741 494904 368788
rect 494804 368707 494837 368741
rect 494871 368707 494904 368741
rect 493317 368105 493343 368505
rect 494633 368452 494659 368505
rect 494804 368452 494904 368707
rect 494633 368341 494904 368452
rect 494633 368332 494837 368341
rect 494633 368105 494659 368332
rect 494804 368307 494837 368332
rect 494871 368307 494904 368341
rect 493317 367647 493343 368047
rect 494633 367996 494659 368047
rect 494804 367996 494904 368307
rect 494633 367941 494904 367996
rect 494633 367907 494837 367941
rect 494871 367907 494904 367941
rect 494633 367876 494904 367907
rect 494633 367647 494659 367876
rect 493317 367189 493343 367589
rect 494633 367540 494659 367589
rect 494804 367541 494904 367876
rect 494804 367540 494837 367541
rect 494633 367507 494837 367540
rect 494871 367507 494904 367541
rect 494633 367420 494904 367507
rect 494633 367189 494659 367420
rect 494804 367141 494904 367420
rect 493317 366731 493343 367131
rect 494633 367084 494659 367131
rect 494804 367107 494837 367141
rect 494871 367107 494904 367141
rect 494804 367084 494904 367107
rect 494633 366964 494904 367084
rect 494633 366731 494659 366964
rect 494804 366741 494904 366964
rect 494804 366707 494837 366741
rect 494871 366707 494904 366741
rect 493317 366273 493343 366673
rect 494633 366628 494659 366673
rect 494804 366628 494904 366707
rect 494633 366508 494904 366628
rect 494633 366273 494659 366508
rect 494804 366341 494904 366508
rect 494804 366307 494837 366341
rect 494871 366307 494904 366341
rect 493317 365815 493343 366215
rect 494633 366172 494659 366215
rect 494804 366172 494904 366307
rect 494633 366052 494904 366172
rect 494633 365815 494659 366052
rect 494804 365941 494904 366052
rect 494804 365907 494837 365941
rect 494871 365907 494904 365941
rect 493317 365357 493343 365757
rect 494633 365716 494659 365757
rect 494804 365716 494904 365907
rect 494633 365596 494904 365716
rect 494633 365357 494659 365596
rect 494804 365541 494904 365596
rect 494804 365507 494837 365541
rect 494871 365507 494904 365541
rect 493317 364899 493343 365299
rect 494633 365260 494659 365299
rect 494804 365260 494904 365507
rect 494633 365141 494904 365260
rect 494633 365140 494837 365141
rect 494633 364899 494659 365140
rect 494804 365107 494837 365140
rect 494871 365107 494904 365141
rect 493317 364441 493343 364841
rect 494633 364804 494659 364841
rect 494804 364804 494904 365107
rect 494633 364741 494904 364804
rect 494633 364707 494837 364741
rect 494871 364707 494904 364741
rect 494633 364684 494904 364707
rect 494633 364441 494659 364684
rect 493317 363983 493343 364383
rect 494633 364348 494659 364383
rect 494804 364348 494904 364684
rect 494633 364341 494904 364348
rect 494633 364307 494837 364341
rect 494871 364307 494904 364341
rect 494633 364228 494904 364307
rect 494633 363983 494659 364228
rect 494804 363941 494904 364228
rect 493317 363525 493343 363925
rect 494633 363892 494659 363925
rect 494804 363907 494837 363941
rect 494871 363907 494904 363941
rect 494804 363892 494904 363907
rect 494633 363772 494904 363892
rect 494633 363525 494659 363772
rect 494804 363541 494904 363772
rect 494804 363507 494837 363541
rect 494871 363507 494904 363541
rect 493317 363067 493343 363467
rect 494633 363436 494659 363467
rect 494804 363436 494904 363507
rect 494633 363316 494904 363436
rect 494633 363067 494659 363316
rect 494804 363141 494904 363316
rect 494804 363107 494837 363141
rect 494871 363107 494904 363141
rect 493317 362609 493343 363009
rect 494633 362980 494659 363009
rect 494804 362980 494904 363107
rect 494633 362860 494904 362980
rect 494633 362609 494659 362860
rect 494804 362741 494904 362860
rect 494804 362707 494837 362741
rect 494871 362707 494904 362741
rect 494804 362516 494904 362707
rect 523397 374517 523423 374917
rect 524713 374836 524739 374917
rect 524884 374836 524984 375107
rect 524713 374741 524984 374836
rect 524713 374716 524917 374741
rect 524713 374517 524739 374716
rect 524884 374707 524917 374716
rect 524951 374707 524984 374741
rect 523397 374059 523423 374459
rect 524713 374380 524739 374459
rect 524884 374380 524984 374707
rect 524713 374341 524984 374380
rect 524713 374307 524917 374341
rect 524951 374307 524984 374341
rect 524713 374260 524984 374307
rect 524713 374059 524739 374260
rect 523397 373601 523423 374001
rect 524713 373924 524739 374001
rect 524884 373941 524984 374260
rect 524884 373924 524917 373941
rect 524713 373907 524917 373924
rect 524951 373907 524984 373941
rect 524713 373804 524984 373907
rect 524713 373601 524739 373804
rect 523397 373143 523423 373543
rect 524713 373468 524739 373543
rect 524884 373541 524984 373804
rect 524884 373507 524917 373541
rect 524951 373507 524984 373541
rect 524884 373468 524984 373507
rect 524713 373348 524984 373468
rect 524713 373143 524739 373348
rect 524884 373141 524984 373348
rect 524884 373107 524917 373141
rect 524951 373107 524984 373141
rect 523397 372685 523423 373085
rect 524713 373012 524739 373085
rect 524884 373012 524984 373107
rect 524713 372892 524984 373012
rect 524713 372685 524739 372892
rect 524884 372741 524984 372892
rect 524884 372707 524917 372741
rect 524951 372707 524984 372741
rect 523397 372227 523423 372627
rect 524713 372556 524739 372627
rect 524884 372556 524984 372707
rect 524713 372436 524984 372556
rect 524713 372227 524739 372436
rect 524884 372341 524984 372436
rect 524884 372307 524917 372341
rect 524951 372307 524984 372341
rect 523397 371769 523423 372169
rect 524713 372100 524739 372169
rect 524884 372100 524984 372307
rect 524713 371980 524984 372100
rect 524713 371769 524739 371980
rect 524884 371941 524984 371980
rect 524884 371907 524917 371941
rect 524951 371907 524984 371941
rect 523397 371311 523423 371711
rect 524713 371644 524739 371711
rect 524884 371644 524984 371907
rect 524713 371541 524984 371644
rect 524713 371524 524917 371541
rect 524713 371311 524739 371524
rect 524884 371507 524917 371524
rect 524951 371507 524984 371541
rect 523397 370853 523423 371253
rect 524713 371188 524739 371253
rect 524884 371188 524984 371507
rect 524713 371141 524984 371188
rect 524713 371107 524917 371141
rect 524951 371107 524984 371141
rect 524713 371068 524984 371107
rect 524713 370853 524739 371068
rect 523397 370395 523423 370795
rect 524713 370732 524739 370795
rect 524884 370741 524984 371068
rect 524884 370732 524917 370741
rect 524713 370707 524917 370732
rect 524951 370707 524984 370741
rect 524713 370612 524984 370707
rect 524713 370395 524739 370612
rect 524884 370341 524984 370612
rect 523397 369937 523423 370337
rect 524713 370276 524739 370337
rect 524884 370307 524917 370341
rect 524951 370307 524984 370341
rect 524884 370276 524984 370307
rect 524713 370156 524984 370276
rect 524713 369937 524739 370156
rect 524884 369941 524984 370156
rect 524884 369907 524917 369941
rect 524951 369907 524984 369941
rect 523397 369479 523423 369879
rect 524713 369820 524739 369879
rect 524884 369820 524984 369907
rect 524713 369700 524984 369820
rect 524713 369479 524739 369700
rect 524884 369541 524984 369700
rect 524884 369507 524917 369541
rect 524951 369507 524984 369541
rect 523397 369021 523423 369421
rect 524713 369364 524739 369421
rect 524884 369364 524984 369507
rect 524713 369244 524984 369364
rect 524713 369021 524739 369244
rect 524884 369141 524984 369244
rect 524884 369107 524917 369141
rect 524951 369107 524984 369141
rect 523397 368563 523423 368963
rect 524713 368908 524739 368963
rect 524884 368908 524984 369107
rect 524713 368788 524984 368908
rect 524713 368563 524739 368788
rect 524884 368741 524984 368788
rect 524884 368707 524917 368741
rect 524951 368707 524984 368741
rect 523397 368105 523423 368505
rect 524713 368452 524739 368505
rect 524884 368452 524984 368707
rect 524713 368341 524984 368452
rect 524713 368332 524917 368341
rect 524713 368105 524739 368332
rect 524884 368307 524917 368332
rect 524951 368307 524984 368341
rect 523397 367647 523423 368047
rect 524713 367996 524739 368047
rect 524884 367996 524984 368307
rect 524713 367941 524984 367996
rect 524713 367907 524917 367941
rect 524951 367907 524984 367941
rect 524713 367876 524984 367907
rect 524713 367647 524739 367876
rect 523397 367189 523423 367589
rect 524713 367540 524739 367589
rect 524884 367541 524984 367876
rect 524884 367540 524917 367541
rect 524713 367507 524917 367540
rect 524951 367507 524984 367541
rect 524713 367420 524984 367507
rect 524713 367189 524739 367420
rect 524884 367141 524984 367420
rect 523397 366731 523423 367131
rect 524713 367084 524739 367131
rect 524884 367107 524917 367141
rect 524951 367107 524984 367141
rect 524884 367084 524984 367107
rect 524713 366964 524984 367084
rect 524713 366731 524739 366964
rect 524884 366741 524984 366964
rect 524884 366707 524917 366741
rect 524951 366707 524984 366741
rect 523397 366273 523423 366673
rect 524713 366628 524739 366673
rect 524884 366628 524984 366707
rect 524713 366508 524984 366628
rect 524713 366273 524739 366508
rect 524884 366341 524984 366508
rect 524884 366307 524917 366341
rect 524951 366307 524984 366341
rect 523397 365815 523423 366215
rect 524713 366172 524739 366215
rect 524884 366172 524984 366307
rect 524713 366052 524984 366172
rect 524713 365815 524739 366052
rect 524884 365941 524984 366052
rect 524884 365907 524917 365941
rect 524951 365907 524984 365941
rect 523397 365357 523423 365757
rect 524713 365716 524739 365757
rect 524884 365716 524984 365907
rect 524713 365596 524984 365716
rect 524713 365357 524739 365596
rect 524884 365541 524984 365596
rect 524884 365507 524917 365541
rect 524951 365507 524984 365541
rect 523397 364899 523423 365299
rect 524713 365260 524739 365299
rect 524884 365260 524984 365507
rect 524713 365141 524984 365260
rect 524713 365140 524917 365141
rect 524713 364899 524739 365140
rect 524884 365107 524917 365140
rect 524951 365107 524984 365141
rect 523397 364441 523423 364841
rect 524713 364804 524739 364841
rect 524884 364804 524984 365107
rect 524713 364741 524984 364804
rect 524713 364707 524917 364741
rect 524951 364707 524984 364741
rect 524713 364684 524984 364707
rect 524713 364441 524739 364684
rect 523397 363983 523423 364383
rect 524713 364348 524739 364383
rect 524884 364348 524984 364684
rect 524713 364341 524984 364348
rect 524713 364307 524917 364341
rect 524951 364307 524984 364341
rect 524713 364228 524984 364307
rect 524713 363983 524739 364228
rect 524884 363941 524984 364228
rect 523397 363525 523423 363925
rect 524713 363892 524739 363925
rect 524884 363907 524917 363941
rect 524951 363907 524984 363941
rect 524884 363892 524984 363907
rect 524713 363772 524984 363892
rect 524713 363525 524739 363772
rect 524884 363541 524984 363772
rect 524884 363507 524917 363541
rect 524951 363507 524984 363541
rect 523397 363067 523423 363467
rect 524713 363436 524739 363467
rect 524884 363436 524984 363507
rect 524713 363316 524984 363436
rect 524713 363067 524739 363316
rect 524884 363141 524984 363316
rect 524884 363107 524917 363141
rect 524951 363107 524984 363141
rect 523397 362609 523423 363009
rect 524713 362980 524739 363009
rect 524884 362980 524984 363107
rect 524713 362860 524984 362980
rect 524713 362609 524739 362860
rect 524884 362741 524984 362860
rect 524884 362707 524917 362741
rect 524951 362707 524984 362741
rect 524884 362516 524984 362707
rect 560599 358980 560799 359006
rect 560857 358980 561057 359006
rect 561115 358980 561315 359006
rect 561373 358980 561573 359006
rect 561631 358980 561831 359006
rect 561889 358980 562089 359006
rect 562147 358980 562347 359006
rect 562405 358980 562605 359006
rect 562663 358980 562863 359006
rect 562921 358980 563121 359006
rect 563179 358980 563379 359006
rect 563437 358980 563637 359006
rect 563695 358980 563895 359006
rect 563953 358980 564153 359006
rect 564211 358980 564411 359006
rect 564469 358980 564669 359006
rect 564727 358980 564927 359006
rect 564985 358980 565185 359006
rect 565243 358980 565443 359006
rect 565501 358980 565701 359006
rect 574737 358910 574937 358936
rect 574995 358910 575195 358936
rect 575253 358910 575453 358936
rect 575511 358910 575711 358936
rect 575769 358910 575969 358936
rect 576027 358910 576227 358936
rect 576285 358910 576485 358936
rect 576543 358910 576743 358936
rect 576801 358910 577001 358936
rect 577059 358910 577259 358936
rect 577317 358910 577517 358936
rect 577575 358910 577775 358936
rect 577833 358910 578033 358936
rect 578091 358910 578291 358936
rect 578349 358910 578549 358936
rect 578607 358910 578807 358936
rect 578865 358910 579065 358936
rect 579123 358910 579323 358936
rect 579381 358910 579581 358936
rect 579639 358910 579839 358936
rect 560599 357954 560799 357980
rect 560857 357954 561057 357980
rect 561115 357954 561315 357980
rect 561373 357954 561573 357980
rect 561631 357954 561831 357980
rect 561889 357954 562089 357980
rect 562147 357954 562347 357980
rect 562405 357954 562605 357980
rect 562663 357954 562863 357980
rect 562921 357954 563121 357980
rect 563179 357954 563379 357980
rect 563437 357954 563637 357980
rect 563695 357954 563895 357980
rect 563953 357954 564153 357980
rect 564211 357954 564411 357980
rect 564469 357954 564669 357980
rect 564727 357954 564927 357980
rect 564985 357954 565185 357980
rect 565243 357954 565443 357980
rect 565501 357954 565701 357980
rect 560654 357764 560774 357954
rect 560910 357764 561030 357954
rect 561166 357764 561286 357954
rect 561422 357764 561542 357954
rect 561678 357764 561798 357954
rect 561934 357764 562054 357954
rect 562190 357764 562310 357954
rect 562446 357764 562566 357954
rect 562702 357764 562822 357954
rect 562958 357764 563078 357954
rect 563214 357764 563334 357954
rect 563470 357764 563590 357954
rect 563726 357764 563846 357954
rect 563982 357764 564102 357954
rect 564238 357764 564358 357954
rect 564494 357764 564614 357954
rect 564750 357764 564870 357954
rect 565006 357764 565126 357954
rect 565262 357764 565382 357954
rect 565518 357764 565638 357954
rect 574737 357884 574937 357910
rect 574995 357884 575195 357910
rect 575253 357884 575453 357910
rect 575511 357884 575711 357910
rect 575769 357884 575969 357910
rect 576027 357884 576227 357910
rect 576285 357884 576485 357910
rect 576543 357884 576743 357910
rect 576801 357884 577001 357910
rect 577059 357884 577259 357910
rect 577317 357884 577517 357910
rect 577575 357884 577775 357910
rect 577833 357884 578033 357910
rect 578091 357884 578291 357910
rect 578349 357884 578549 357910
rect 578607 357884 578807 357910
rect 578865 357884 579065 357910
rect 579123 357884 579323 357910
rect 579381 357884 579581 357910
rect 579639 357884 579839 357910
rect 560542 357744 565678 357764
rect 560542 357684 560728 357744
rect 560788 357684 560928 357744
rect 560988 357684 561128 357744
rect 561188 357684 561328 357744
rect 561388 357684 561528 357744
rect 561588 357684 561728 357744
rect 561788 357684 561928 357744
rect 561988 357684 562128 357744
rect 562188 357684 562328 357744
rect 562388 357684 562528 357744
rect 562588 357684 562728 357744
rect 562788 357684 562928 357744
rect 562988 357684 563128 357744
rect 563188 357684 563328 357744
rect 563388 357684 563528 357744
rect 563588 357684 563728 357744
rect 563788 357684 563928 357744
rect 563988 357684 564128 357744
rect 564188 357684 564328 357744
rect 564388 357684 564528 357744
rect 564588 357684 564728 357744
rect 564788 357684 564928 357744
rect 564988 357684 565128 357744
rect 565188 357684 565328 357744
rect 565388 357684 565528 357744
rect 565588 357684 565678 357744
rect 560542 357664 565678 357684
rect 574808 357638 574928 357884
rect 575064 357638 575184 357884
rect 575320 357638 575440 357884
rect 575576 357638 575696 357884
rect 575832 357638 575952 357884
rect 576088 357638 576208 357884
rect 576344 357638 576464 357884
rect 576600 357638 576720 357884
rect 576856 357638 576976 357884
rect 577112 357638 577232 357884
rect 577368 357638 577488 357884
rect 577624 357638 577744 357884
rect 577880 357638 578000 357884
rect 578136 357638 578256 357884
rect 578392 357638 578512 357884
rect 578648 357638 578768 357884
rect 578904 357638 579024 357884
rect 579160 357638 579280 357884
rect 579416 357638 579536 357884
rect 579672 357638 579792 357884
rect 574644 357618 579932 357638
rect 574644 357558 574702 357618
rect 574762 357558 574902 357618
rect 574962 357558 575102 357618
rect 575162 357558 575302 357618
rect 575362 357558 575502 357618
rect 575562 357558 575702 357618
rect 575762 357558 575902 357618
rect 575962 357558 576102 357618
rect 576162 357558 576302 357618
rect 576362 357558 576502 357618
rect 576562 357558 576702 357618
rect 576762 357558 576902 357618
rect 576962 357558 577102 357618
rect 577162 357558 577302 357618
rect 577362 357558 577502 357618
rect 577562 357558 577702 357618
rect 577762 357558 577902 357618
rect 577962 357558 578102 357618
rect 578162 357558 578302 357618
rect 578362 357558 578502 357618
rect 578562 357558 578702 357618
rect 578762 357558 578902 357618
rect 578962 357558 579102 357618
rect 579162 357558 579302 357618
rect 579362 357558 579502 357618
rect 579562 357558 579702 357618
rect 579762 357558 579932 357618
rect 574644 357538 579932 357558
rect 575185 312742 575385 312768
rect 575443 312742 575643 312768
rect 575701 312742 575901 312768
rect 575959 312742 576159 312768
rect 576217 312742 576417 312768
rect 576475 312742 576675 312768
rect 576733 312742 576933 312768
rect 576991 312742 577191 312768
rect 577249 312742 577449 312768
rect 577507 312742 577707 312768
rect 577765 312742 577965 312768
rect 578023 312742 578223 312768
rect 578281 312742 578481 312768
rect 578539 312742 578739 312768
rect 578797 312742 578997 312768
rect 579055 312742 579255 312768
rect 579313 312742 579513 312768
rect 579571 312742 579771 312768
rect 579829 312742 580029 312768
rect 580087 312742 580287 312768
rect 560461 312672 560661 312698
rect 560719 312672 560919 312698
rect 560977 312672 561177 312698
rect 561235 312672 561435 312698
rect 561493 312672 561693 312698
rect 561751 312672 561951 312698
rect 562009 312672 562209 312698
rect 562267 312672 562467 312698
rect 562525 312672 562725 312698
rect 562783 312672 562983 312698
rect 563041 312672 563241 312698
rect 563299 312672 563499 312698
rect 563557 312672 563757 312698
rect 563815 312672 564015 312698
rect 564073 312672 564273 312698
rect 564331 312672 564531 312698
rect 564589 312672 564789 312698
rect 564847 312672 565047 312698
rect 565105 312672 565305 312698
rect 565363 312672 565563 312698
rect 575185 311716 575385 311742
rect 575443 311716 575643 311742
rect 575701 311716 575901 311742
rect 575959 311716 576159 311742
rect 576217 311716 576417 311742
rect 576475 311716 576675 311742
rect 576733 311716 576933 311742
rect 576991 311716 577191 311742
rect 577249 311716 577449 311742
rect 577507 311716 577707 311742
rect 577765 311716 577965 311742
rect 578023 311716 578223 311742
rect 578281 311716 578481 311742
rect 578539 311716 578739 311742
rect 578797 311716 578997 311742
rect 579055 311716 579255 311742
rect 579313 311716 579513 311742
rect 579571 311716 579771 311742
rect 579829 311716 580029 311742
rect 580087 311716 580287 311742
rect 560461 311646 560661 311672
rect 560719 311646 560919 311672
rect 560977 311646 561177 311672
rect 561235 311646 561435 311672
rect 561493 311646 561693 311672
rect 561751 311646 561951 311672
rect 562009 311646 562209 311672
rect 562267 311646 562467 311672
rect 562525 311646 562725 311672
rect 562783 311646 562983 311672
rect 563041 311646 563241 311672
rect 563299 311646 563499 311672
rect 563557 311646 563757 311672
rect 563815 311646 564015 311672
rect 564073 311646 564273 311672
rect 564331 311646 564531 311672
rect 564589 311646 564789 311672
rect 564847 311646 565047 311672
rect 565105 311646 565305 311672
rect 565363 311646 565563 311672
rect 560516 311456 560636 311646
rect 560772 311456 560892 311646
rect 561028 311456 561148 311646
rect 561284 311456 561404 311646
rect 561540 311456 561660 311646
rect 561796 311456 561916 311646
rect 562052 311456 562172 311646
rect 562308 311456 562428 311646
rect 562564 311456 562684 311646
rect 562820 311456 562940 311646
rect 563076 311456 563196 311646
rect 563332 311456 563452 311646
rect 563588 311456 563708 311646
rect 563844 311456 563964 311646
rect 564100 311456 564220 311646
rect 564356 311456 564476 311646
rect 564612 311456 564732 311646
rect 564868 311456 564988 311646
rect 565124 311456 565244 311646
rect 565380 311456 565500 311646
rect 575256 311470 575376 311716
rect 575512 311470 575632 311716
rect 575768 311470 575888 311716
rect 576024 311470 576144 311716
rect 576280 311470 576400 311716
rect 576536 311470 576656 311716
rect 576792 311470 576912 311716
rect 577048 311470 577168 311716
rect 577304 311470 577424 311716
rect 577560 311470 577680 311716
rect 577816 311470 577936 311716
rect 578072 311470 578192 311716
rect 578328 311470 578448 311716
rect 578584 311470 578704 311716
rect 578840 311470 578960 311716
rect 579096 311470 579216 311716
rect 579352 311470 579472 311716
rect 579608 311470 579728 311716
rect 579864 311470 579984 311716
rect 580120 311470 580240 311716
rect 560404 311436 565540 311456
rect 560404 311376 560590 311436
rect 560650 311376 560790 311436
rect 560850 311376 560990 311436
rect 561050 311376 561190 311436
rect 561250 311376 561390 311436
rect 561450 311376 561590 311436
rect 561650 311376 561790 311436
rect 561850 311376 561990 311436
rect 562050 311376 562190 311436
rect 562250 311376 562390 311436
rect 562450 311376 562590 311436
rect 562650 311376 562790 311436
rect 562850 311376 562990 311436
rect 563050 311376 563190 311436
rect 563250 311376 563390 311436
rect 563450 311376 563590 311436
rect 563650 311376 563790 311436
rect 563850 311376 563990 311436
rect 564050 311376 564190 311436
rect 564250 311376 564390 311436
rect 564450 311376 564590 311436
rect 564650 311376 564790 311436
rect 564850 311376 564990 311436
rect 565050 311376 565190 311436
rect 565250 311376 565390 311436
rect 565450 311376 565540 311436
rect 560404 311356 565540 311376
rect 575092 311450 580380 311470
rect 575092 311390 575150 311450
rect 575210 311390 575350 311450
rect 575410 311390 575550 311450
rect 575610 311390 575750 311450
rect 575810 311390 575950 311450
rect 576010 311390 576150 311450
rect 576210 311390 576350 311450
rect 576410 311390 576550 311450
rect 576610 311390 576750 311450
rect 576810 311390 576950 311450
rect 577010 311390 577150 311450
rect 577210 311390 577350 311450
rect 577410 311390 577550 311450
rect 577610 311390 577750 311450
rect 577810 311390 577950 311450
rect 578010 311390 578150 311450
rect 578210 311390 578350 311450
rect 578410 311390 578550 311450
rect 578610 311390 578750 311450
rect 578810 311390 578950 311450
rect 579010 311390 579150 311450
rect 579210 311390 579350 311450
rect 579410 311390 579550 311450
rect 579610 311390 579750 311450
rect 579810 311390 579950 311450
rect 580010 311390 580150 311450
rect 580210 311390 580380 311450
rect 575092 311370 580380 311390
<< polycont >>
rect 560836 492144 560896 492204
rect 561036 492144 561096 492204
rect 561236 492144 561296 492204
rect 561436 492144 561496 492204
rect 561636 492144 561696 492204
rect 561836 492144 561896 492204
rect 562036 492144 562096 492204
rect 562236 492144 562296 492204
rect 562436 492144 562496 492204
rect 562636 492144 562696 492204
rect 562836 492144 562896 492204
rect 563036 492144 563096 492204
rect 563236 492144 563296 492204
rect 563436 492144 563496 492204
rect 563636 492144 563696 492204
rect 563836 492144 563896 492204
rect 564036 492144 564096 492204
rect 564236 492144 564296 492204
rect 564436 492144 564496 492204
rect 564636 492144 564696 492204
rect 564836 492144 564896 492204
rect 565036 492144 565096 492204
rect 565236 492144 565296 492204
rect 565436 492144 565496 492204
rect 565636 492144 565696 492204
rect 575228 491862 575288 491922
rect 575428 491862 575488 491922
rect 575628 491862 575688 491922
rect 575828 491862 575888 491922
rect 576028 491862 576088 491922
rect 576228 491862 576288 491922
rect 576428 491862 576488 491922
rect 576628 491862 576688 491922
rect 576828 491862 576888 491922
rect 577028 491862 577088 491922
rect 577228 491862 577288 491922
rect 577428 491862 577488 491922
rect 577628 491862 577688 491922
rect 577828 491862 577888 491922
rect 578028 491862 578088 491922
rect 578228 491862 578288 491922
rect 578428 491862 578488 491922
rect 578628 491862 578688 491922
rect 578828 491862 578888 491922
rect 579028 491862 579088 491922
rect 579228 491862 579288 491922
rect 579428 491862 579488 491922
rect 579628 491862 579688 491922
rect 579828 491862 579888 491922
rect 580028 491862 580088 491922
rect 580228 491862 580288 491922
rect 560860 403002 560920 403062
rect 561060 403002 561120 403062
rect 561260 403002 561320 403062
rect 561460 403002 561520 403062
rect 561660 403002 561720 403062
rect 561860 403002 561920 403062
rect 562060 403002 562120 403062
rect 562260 403002 562320 403062
rect 562460 403002 562520 403062
rect 562660 403002 562720 403062
rect 562860 403002 562920 403062
rect 563060 403002 563120 403062
rect 563260 403002 563320 403062
rect 563460 403002 563520 403062
rect 563660 403002 563720 403062
rect 563860 403002 563920 403062
rect 564060 403002 564120 403062
rect 564260 403002 564320 403062
rect 564460 403002 564520 403062
rect 564660 403002 564720 403062
rect 564860 403002 564920 403062
rect 565060 403002 565120 403062
rect 565260 403002 565320 403062
rect 565460 403002 565520 403062
rect 565660 403002 565720 403062
rect 574506 402986 574566 403046
rect 574706 402986 574766 403046
rect 574906 402986 574966 403046
rect 575106 402986 575166 403046
rect 575306 402986 575366 403046
rect 575506 402986 575566 403046
rect 575706 402986 575766 403046
rect 575906 402986 575966 403046
rect 576106 402986 576166 403046
rect 576306 402986 576366 403046
rect 576506 402986 576566 403046
rect 576706 402986 576766 403046
rect 576906 402986 576966 403046
rect 577106 402986 577166 403046
rect 577306 402986 577366 403046
rect 577506 402986 577566 403046
rect 577706 402986 577766 403046
rect 577906 402986 577966 403046
rect 578106 402986 578166 403046
rect 578306 402986 578366 403046
rect 578506 402986 578566 403046
rect 578706 402986 578766 403046
rect 578906 402986 578966 403046
rect 579106 402986 579166 403046
rect 579306 402986 579366 403046
rect 579506 402986 579566 403046
rect 498557 400619 498591 400653
rect 498597 399707 498631 399741
rect 498597 399307 498631 399341
rect 498597 398907 498631 398941
rect 498597 398507 498631 398541
rect 498597 398107 498631 398141
rect 498597 397707 498631 397741
rect 498597 397307 498631 397341
rect 498597 396907 498631 396941
rect 498597 396507 498631 396541
rect 498597 396107 498631 396141
rect 498597 395707 498631 395741
rect 498597 395307 498631 395341
rect 498597 394907 498631 394941
rect 498597 394507 498631 394541
rect 498597 394107 498631 394141
rect 498597 393707 498631 393741
rect 498597 393307 498631 393341
rect 498597 392907 498631 392941
rect 498597 392507 498631 392541
rect 498597 392107 498631 392141
rect 502357 392063 502391 392097
rect 498597 391707 498631 391741
rect 498597 391307 498631 391341
rect 502357 391663 502391 391697
rect 494797 390819 494831 390853
rect 498597 390907 498631 390941
rect 502357 391263 502391 391297
rect 502357 390863 502391 390897
rect 498597 390507 498631 390541
rect 494837 389907 494871 389941
rect 502357 390463 502391 390497
rect 498597 390107 498631 390141
rect 494837 389507 494871 389541
rect 502357 390063 502391 390097
rect 498597 389707 498631 389741
rect 502357 389663 502391 389697
rect 498597 389307 498631 389341
rect 494837 389107 494871 389141
rect 502357 389263 502391 389297
rect 498597 388907 498631 388941
rect 494837 388707 494871 388741
rect 505917 389319 505951 389353
rect 502357 388863 502391 388897
rect 498597 388507 498631 388541
rect 494837 388307 494871 388341
rect 498597 388107 498631 388141
rect 517197 389319 517231 389353
rect 505917 388919 505951 388953
rect 502357 388463 502391 388497
rect 494837 387907 494871 387941
rect 494837 387507 494871 387541
rect 517197 388919 517231 388953
rect 505917 388519 505951 388553
rect 524917 389907 524951 389941
rect 524917 389507 524951 389541
rect 524917 389107 524951 389141
rect 524917 388707 524951 388741
rect 517197 388519 517231 388553
rect 505917 388119 505951 388153
rect 498597 387707 498631 387741
rect 494837 387107 494871 387141
rect 502357 388063 502391 388097
rect 524917 388307 524951 388341
rect 517197 388119 517231 388153
rect 505917 387719 505951 387753
rect 502357 387663 502391 387697
rect 498597 387307 498631 387341
rect 494837 386707 494871 386741
rect 502357 387263 502391 387297
rect 498597 386907 498631 386941
rect 494837 386307 494871 386341
rect 505917 387319 505951 387353
rect 502357 386863 502391 386897
rect 505917 386919 505951 386953
rect 498597 386507 498631 386541
rect 505917 386519 505951 386553
rect 498597 386107 498631 386141
rect 494837 385907 494871 385941
rect 505917 386119 505951 386153
rect 498597 385707 498631 385741
rect 494837 385507 494871 385541
rect 498597 385307 498631 385341
rect 494837 385107 494871 385141
rect 502357 385399 502391 385433
rect 505917 385719 505951 385753
rect 517197 387719 517231 387753
rect 524917 387907 524951 387941
rect 517197 387319 517231 387353
rect 517197 386919 517231 386953
rect 517197 386519 517231 386553
rect 517197 386119 517231 386153
rect 517197 385719 517231 385753
rect 524917 387507 524951 387541
rect 524917 387107 524951 387141
rect 524917 386707 524951 386741
rect 524917 386307 524951 386341
rect 524917 385907 524951 385941
rect 524917 385507 524951 385541
rect 498597 384907 498631 384941
rect 494837 384707 494871 384741
rect 494837 384307 494871 384341
rect 524917 385107 524951 385141
rect 502357 384999 502391 385033
rect 498597 384507 498631 384541
rect 494837 383907 494871 383941
rect 502357 384599 502391 384633
rect 502357 384199 502391 384233
rect 498597 384107 498631 384141
rect 494837 383507 494871 383541
rect 502357 383799 502391 383833
rect 498597 383707 498631 383741
rect 494837 383107 494871 383141
rect 498597 383307 498631 383341
rect 502357 383399 502391 383433
rect 498597 382907 498631 382941
rect 494837 382707 494871 382741
rect 502357 382999 502391 383033
rect 498597 382507 498631 382541
rect 494837 382307 494871 382341
rect 502357 382599 502391 382633
rect 524917 384707 524951 384741
rect 524917 384307 524951 384341
rect 524917 383907 524951 383941
rect 524917 383507 524951 383541
rect 524917 383107 524951 383141
rect 524917 382707 524951 382741
rect 498597 382107 498631 382141
rect 494837 381907 494871 381941
rect 524917 382307 524951 382341
rect 502357 382199 502391 382233
rect 498597 381707 498631 381741
rect 494837 381507 494871 381541
rect 494837 381107 494871 381141
rect 524917 381907 524951 381941
rect 502357 381799 502391 381833
rect 498597 381307 498631 381341
rect 494837 380707 494871 380741
rect 502357 381399 502391 381433
rect 502357 380999 502391 381033
rect 498597 380907 498631 380941
rect 494837 380307 494871 380341
rect 502357 380599 502391 380633
rect 498597 380507 498631 380541
rect 494837 379907 494871 379941
rect 498597 380107 498631 380141
rect 502357 380199 502391 380233
rect 498597 379707 498631 379741
rect 494837 379507 494871 379541
rect 498597 379307 498631 379341
rect 524917 381507 524951 381541
rect 524917 381107 524951 381141
rect 524917 380707 524951 380741
rect 524917 380307 524951 380341
rect 524917 379907 524951 379941
rect 524917 379507 524951 379541
rect 494837 379107 494871 379141
rect 524917 379107 524951 379141
rect 498597 378907 498631 378941
rect 494837 378707 494871 378741
rect 524917 378707 524951 378741
rect 498597 378507 498631 378541
rect 494837 378307 494871 378341
rect 494837 377907 494871 377941
rect 524917 378307 524951 378341
rect 498597 378107 498631 378141
rect 494837 377507 494871 377541
rect 498597 377707 498631 377741
rect 524917 377907 524951 377941
rect 494837 377107 494871 377141
rect 498597 377307 498631 377341
rect 502157 377461 502191 377495
rect 494837 376707 494871 376741
rect 498597 376907 498631 376941
rect 502157 377061 502191 377095
rect 506117 377265 506151 377299
rect 498597 376507 498631 376541
rect 494837 376307 494871 376341
rect 502157 376661 502191 376695
rect 513637 377265 513671 377299
rect 506117 376865 506151 376899
rect 513637 376865 513671 376899
rect 502157 376261 502191 376295
rect 498597 376107 498631 376141
rect 494837 375907 494871 375941
rect 506117 376465 506151 376499
rect 506117 376065 506151 376099
rect 513637 376465 513671 376499
rect 502157 375861 502191 375895
rect 498597 375707 498631 375741
rect 494837 375507 494871 375541
rect 513637 376065 513671 376099
rect 506117 375665 506151 375699
rect 502157 375461 502191 375495
rect 498597 375307 498631 375341
rect 494837 375107 494871 375141
rect 494837 374707 494871 374741
rect 498597 374907 498631 374941
rect 513637 375665 513671 375699
rect 506117 375265 506151 375299
rect 502157 375061 502191 375095
rect 494837 374307 494871 374341
rect 498597 374507 498631 374541
rect 494837 373907 494871 373941
rect 513637 375265 513671 375299
rect 506117 374865 506151 374899
rect 502157 374661 502191 374695
rect 498597 374107 498631 374141
rect 524917 377507 524951 377541
rect 524917 377107 524951 377141
rect 524917 376707 524951 376741
rect 524917 376307 524951 376341
rect 524917 375907 524951 375941
rect 524917 375507 524951 375541
rect 524917 375107 524951 375141
rect 513637 374865 513671 374899
rect 502157 374261 502191 374295
rect 494837 373507 494871 373541
rect 498597 373707 498631 373741
rect 502157 373861 502191 373895
rect 498597 373307 498631 373341
rect 494837 373107 494871 373141
rect 498597 372907 498631 372941
rect 494837 372707 494871 372741
rect 498597 372507 498631 372541
rect 494837 372307 494871 372341
rect 494837 371907 494871 371941
rect 494837 371507 494871 371541
rect 494837 371107 494871 371141
rect 494837 370707 494871 370741
rect 494837 370307 494871 370341
rect 494837 369907 494871 369941
rect 494837 369507 494871 369541
rect 494837 369107 494871 369141
rect 494837 368707 494871 368741
rect 494837 368307 494871 368341
rect 494837 367907 494871 367941
rect 494837 367507 494871 367541
rect 494837 367107 494871 367141
rect 494837 366707 494871 366741
rect 494837 366307 494871 366341
rect 494837 365907 494871 365941
rect 494837 365507 494871 365541
rect 494837 365107 494871 365141
rect 494837 364707 494871 364741
rect 494837 364307 494871 364341
rect 494837 363907 494871 363941
rect 494837 363507 494871 363541
rect 494837 363107 494871 363141
rect 494837 362707 494871 362741
rect 524917 374707 524951 374741
rect 524917 374307 524951 374341
rect 524917 373907 524951 373941
rect 524917 373507 524951 373541
rect 524917 373107 524951 373141
rect 524917 372707 524951 372741
rect 524917 372307 524951 372341
rect 524917 371907 524951 371941
rect 524917 371507 524951 371541
rect 524917 371107 524951 371141
rect 524917 370707 524951 370741
rect 524917 370307 524951 370341
rect 524917 369907 524951 369941
rect 524917 369507 524951 369541
rect 524917 369107 524951 369141
rect 524917 368707 524951 368741
rect 524917 368307 524951 368341
rect 524917 367907 524951 367941
rect 524917 367507 524951 367541
rect 524917 367107 524951 367141
rect 524917 366707 524951 366741
rect 524917 366307 524951 366341
rect 524917 365907 524951 365941
rect 524917 365507 524951 365541
rect 524917 365107 524951 365141
rect 524917 364707 524951 364741
rect 524917 364307 524951 364341
rect 524917 363907 524951 363941
rect 524917 363507 524951 363541
rect 524917 363107 524951 363141
rect 524917 362707 524951 362741
rect 560728 357684 560788 357744
rect 560928 357684 560988 357744
rect 561128 357684 561188 357744
rect 561328 357684 561388 357744
rect 561528 357684 561588 357744
rect 561728 357684 561788 357744
rect 561928 357684 561988 357744
rect 562128 357684 562188 357744
rect 562328 357684 562388 357744
rect 562528 357684 562588 357744
rect 562728 357684 562788 357744
rect 562928 357684 562988 357744
rect 563128 357684 563188 357744
rect 563328 357684 563388 357744
rect 563528 357684 563588 357744
rect 563728 357684 563788 357744
rect 563928 357684 563988 357744
rect 564128 357684 564188 357744
rect 564328 357684 564388 357744
rect 564528 357684 564588 357744
rect 564728 357684 564788 357744
rect 564928 357684 564988 357744
rect 565128 357684 565188 357744
rect 565328 357684 565388 357744
rect 565528 357684 565588 357744
rect 574702 357558 574762 357618
rect 574902 357558 574962 357618
rect 575102 357558 575162 357618
rect 575302 357558 575362 357618
rect 575502 357558 575562 357618
rect 575702 357558 575762 357618
rect 575902 357558 575962 357618
rect 576102 357558 576162 357618
rect 576302 357558 576362 357618
rect 576502 357558 576562 357618
rect 576702 357558 576762 357618
rect 576902 357558 576962 357618
rect 577102 357558 577162 357618
rect 577302 357558 577362 357618
rect 577502 357558 577562 357618
rect 577702 357558 577762 357618
rect 577902 357558 577962 357618
rect 578102 357558 578162 357618
rect 578302 357558 578362 357618
rect 578502 357558 578562 357618
rect 578702 357558 578762 357618
rect 578902 357558 578962 357618
rect 579102 357558 579162 357618
rect 579302 357558 579362 357618
rect 579502 357558 579562 357618
rect 579702 357558 579762 357618
rect 560590 311376 560650 311436
rect 560790 311376 560850 311436
rect 560990 311376 561050 311436
rect 561190 311376 561250 311436
rect 561390 311376 561450 311436
rect 561590 311376 561650 311436
rect 561790 311376 561850 311436
rect 561990 311376 562050 311436
rect 562190 311376 562250 311436
rect 562390 311376 562450 311436
rect 562590 311376 562650 311436
rect 562790 311376 562850 311436
rect 562990 311376 563050 311436
rect 563190 311376 563250 311436
rect 563390 311376 563450 311436
rect 563590 311376 563650 311436
rect 563790 311376 563850 311436
rect 563990 311376 564050 311436
rect 564190 311376 564250 311436
rect 564390 311376 564450 311436
rect 564590 311376 564650 311436
rect 564790 311376 564850 311436
rect 564990 311376 565050 311436
rect 565190 311376 565250 311436
rect 565390 311376 565450 311436
rect 575150 311390 575210 311450
rect 575350 311390 575410 311450
rect 575550 311390 575610 311450
rect 575750 311390 575810 311450
rect 575950 311390 576010 311450
rect 576150 311390 576210 311450
rect 576350 311390 576410 311450
rect 576550 311390 576610 311450
rect 576750 311390 576810 311450
rect 576950 311390 577010 311450
rect 577150 311390 577210 311450
rect 577350 311390 577410 311450
rect 577550 311390 577610 311450
rect 577750 311390 577810 311450
rect 577950 311390 578010 311450
rect 578150 311390 578210 311450
rect 578350 311390 578410 311450
rect 578550 311390 578610 311450
rect 578750 311390 578810 311450
rect 578950 311390 579010 311450
rect 579150 311390 579210 311450
rect 579350 311390 579410 311450
rect 579550 311390 579610 311450
rect 579750 311390 579810 311450
rect 579950 311390 580010 311450
rect 580150 311390 580210 311450
<< xpolycontact >>
rect 504623 400844 505193 401276
rect 505583 400844 506153 401276
rect 504623 398836 505193 399268
rect 505583 398836 506153 399268
rect 504623 398100 505193 398532
rect 505583 398100 506153 398532
rect 504623 396092 505193 396524
rect 505583 396092 506153 396524
rect 512143 398002 512713 398434
rect 513103 398002 513673 398434
rect 512143 395994 512713 396426
rect 513103 395994 513673 396426
rect 493343 393690 493913 394122
rect 494303 393690 494873 394122
rect 493343 391682 493913 392114
rect 504623 395355 505193 395787
rect 505583 395355 506153 395787
rect 504623 392773 505193 393205
rect 508383 395258 508953 395690
rect 509343 395258 509913 395690
rect 508383 393250 508953 393682
rect 509343 393250 509913 393682
rect 512143 395258 512713 395690
rect 513103 395258 513673 395690
rect 512143 393250 512713 393682
rect 513103 393250 513673 393682
rect 505583 392773 506153 393205
rect 494303 391682 494873 392114
rect 508383 392513 508953 392945
rect 504623 392024 505193 392456
rect 505583 392024 506153 392456
rect 504623 390016 505193 390448
rect 505583 390016 506153 390448
rect 509343 392513 509913 392945
rect 508383 389931 508953 390363
rect 512143 392514 512713 392946
rect 513103 392514 513673 392946
rect 512143 390506 512713 390938
rect 513103 390506 513673 390938
rect 515903 392122 516473 392554
rect 516863 392122 517433 392554
rect 509343 389931 509913 390363
rect 515903 390114 516473 390546
rect 516863 390114 517433 390546
rect 519663 390652 520233 391084
rect 520623 390652 521193 391084
rect 519663 388644 520233 389076
rect 520623 388644 521193 389076
rect 512143 387320 512713 387752
rect 513103 387320 513673 387752
rect 512143 385312 512713 385744
rect 519663 387320 520233 387752
rect 513103 385312 513673 385744
rect 520623 387320 521193 387752
rect 519663 385312 520233 385744
rect 520623 385312 521193 385744
rect 519663 384576 520233 385008
rect 520623 384576 521193 385008
rect 519663 382568 520233 383000
rect 520623 382568 521193 383000
rect 519663 381342 520233 381774
rect 520623 381342 521193 381774
rect 519663 379334 520233 379766
rect 520623 379334 521193 379766
rect 515903 377128 516473 377560
rect 516863 377128 517433 377560
rect 515903 375120 516473 375552
rect 516863 375120 517433 375552
rect 519663 377128 520233 377560
rect 520623 377128 521193 377560
rect 519663 375120 520233 375552
rect 520623 375120 521193 375552
rect 515903 374384 516473 374816
rect 516863 374384 517433 374816
rect 515903 372376 516473 372808
rect 516863 372376 517433 372808
rect 519663 374384 520233 374816
rect 520623 374384 521193 374816
rect 519663 372376 520233 372808
rect 520623 372376 521193 372808
rect 515903 371640 516473 372072
rect 516863 371640 517433 372072
rect 515903 369632 516473 370064
rect 516863 369632 517433 370064
rect 515903 368896 516473 369328
rect 516863 368896 517433 369328
rect 515903 366888 516473 367320
rect 527183 370660 527753 371092
rect 528143 370660 528713 371092
rect 527183 368652 527753 369084
rect 528143 368652 528713 369084
rect 530943 370758 531513 371190
rect 531903 370758 532473 371190
rect 530943 368750 531513 369182
rect 531903 368750 532473 369182
rect 534703 369974 535273 370406
rect 516863 366888 517433 367320
rect 515903 366152 516473 366584
rect 516863 366152 517433 366584
rect 515903 364144 516473 364576
rect 516863 364144 517433 364576
rect 519663 366152 520233 366584
rect 520623 366152 521193 366584
rect 519663 364144 520233 364576
rect 527183 367916 527753 368348
rect 528143 367916 528713 368348
rect 527183 365908 527753 366340
rect 528143 365908 528713 366340
rect 530943 368014 531513 368446
rect 531903 368014 532473 368446
rect 530943 366006 531513 366438
rect 535663 369974 536233 370406
rect 534703 367966 535273 368398
rect 535663 367966 536233 368398
rect 531903 366006 532473 366438
rect 534703 367230 535273 367662
rect 520623 364144 521193 364576
rect 527183 365172 527753 365604
rect 528143 365172 528713 365604
rect 527183 363164 527753 363596
rect 528143 363164 528713 363596
rect 530943 365270 531513 365702
rect 531903 365270 532473 365702
rect 530943 363262 531513 363694
rect 535663 367230 536233 367662
rect 534703 365222 535273 365654
rect 535663 365222 536233 365654
rect 531903 363262 532473 363694
rect 534703 364486 535273 364918
rect 535663 364486 536233 364918
rect 534703 362478 535273 362910
rect 535663 362478 536233 362910
<< xpolyres >>
rect 504623 399268 505193 400844
rect 505583 399268 506153 400844
rect 504623 396524 505193 398100
rect 505583 396524 506153 398100
rect 512143 396426 512713 398002
rect 513103 396426 513673 398002
rect 493343 392114 493913 393690
rect 494303 392114 494873 393690
rect 504623 393205 505193 395355
rect 505583 393205 506153 395355
rect 508383 393682 508953 395258
rect 509343 393682 509913 395258
rect 512143 393682 512713 395258
rect 513103 393682 513673 395258
rect 504623 390448 505193 392024
rect 505583 390448 506153 392024
rect 508383 390363 508953 392513
rect 509343 390363 509913 392513
rect 512143 390938 512713 392514
rect 513103 390938 513673 392514
rect 515903 390546 516473 392122
rect 516863 390546 517433 392122
rect 519663 389076 520233 390652
rect 520623 389076 521193 390652
rect 512143 385744 512713 387320
rect 513103 385744 513673 387320
rect 519663 385744 520233 387320
rect 520623 385744 521193 387320
rect 519663 383000 520233 384576
rect 520623 383000 521193 384576
rect 519663 379766 520233 381342
rect 520623 379766 521193 381342
rect 515903 375552 516473 377128
rect 516863 375552 517433 377128
rect 519663 375552 520233 377128
rect 520623 375552 521193 377128
rect 515903 372808 516473 374384
rect 516863 372808 517433 374384
rect 519663 372808 520233 374384
rect 520623 372808 521193 374384
rect 515903 370064 516473 371640
rect 516863 370064 517433 371640
rect 515903 367320 516473 368896
rect 516863 367320 517433 368896
rect 527183 369084 527753 370660
rect 528143 369084 528713 370660
rect 530943 369182 531513 370758
rect 531903 369182 532473 370758
rect 515903 364576 516473 366152
rect 516863 364576 517433 366152
rect 519663 364576 520233 366152
rect 520623 364576 521193 366152
rect 527183 366340 527753 367916
rect 528143 366340 528713 367916
rect 530943 366438 531513 368014
rect 531903 366438 532473 368014
rect 534703 368398 535273 369974
rect 535663 368398 536233 369974
rect 527183 363596 527753 365172
rect 528143 363596 528713 365172
rect 530943 363694 531513 365270
rect 531903 363694 532473 365270
rect 534703 365654 535273 367230
rect 535663 365654 536233 367230
rect 534703 362910 535273 364486
rect 535663 362910 536233 364486
<< locali >>
rect 560650 493790 560836 493850
rect 560896 493790 561036 493850
rect 561096 493790 561236 493850
rect 561296 493790 561436 493850
rect 561496 493790 561636 493850
rect 561696 493790 561836 493850
rect 561896 493790 562036 493850
rect 562096 493790 562236 493850
rect 562296 493790 562436 493850
rect 562496 493790 562636 493850
rect 562696 493790 562836 493850
rect 562896 493790 563036 493850
rect 563096 493790 563236 493850
rect 563296 493790 563436 493850
rect 563496 493790 563636 493850
rect 563696 493790 563836 493850
rect 563896 493790 564036 493850
rect 564096 493790 564236 493850
rect 564296 493790 564436 493850
rect 564496 493790 564636 493850
rect 564696 493790 564836 493850
rect 564896 493790 565036 493850
rect 565096 493790 565236 493850
rect 565296 493790 565436 493850
rect 565496 493790 565636 493850
rect 565696 493790 565964 493850
rect 560388 493690 560448 493692
rect 560388 493630 565866 493690
rect 560388 492522 560482 493630
rect 560342 492504 560482 492522
rect 560330 492482 560482 492504
rect 560330 492332 560340 492482
rect 560472 492332 560482 492482
rect 560661 493428 560695 493444
rect 560661 492436 560695 492452
rect 560919 493428 560953 493630
rect 560919 492436 560953 492452
rect 561177 493428 561211 493444
rect 561177 492370 561211 492452
rect 561435 493428 561469 493630
rect 561435 492436 561469 492452
rect 561693 493428 561727 493444
rect 561693 492370 561727 492452
rect 561951 493428 561985 493630
rect 561951 492436 561985 492452
rect 562209 493428 562243 493444
rect 562209 492370 562243 492452
rect 562467 493428 562501 493630
rect 562467 492436 562501 492452
rect 562725 493428 562759 493444
rect 562725 492370 562759 492452
rect 562983 493428 563017 493630
rect 562983 492436 563017 492452
rect 563241 493428 563275 493444
rect 563241 492370 563275 492452
rect 563499 493428 563533 493630
rect 563499 492436 563533 492452
rect 563757 493428 563791 493444
rect 563757 492370 563791 492452
rect 564015 493428 564049 493630
rect 564015 492436 564049 492452
rect 564273 493428 564307 493444
rect 564273 492370 564307 492452
rect 564531 493428 564565 493630
rect 564531 492436 564565 492452
rect 564789 493428 564823 493444
rect 564789 492370 564823 492452
rect 565047 493428 565081 493630
rect 565047 492436 565081 492452
rect 565305 493428 565339 493444
rect 565305 492370 565339 492452
rect 565563 493428 565597 493630
rect 575170 493564 575228 493624
rect 575288 493564 575428 493624
rect 575488 493564 575628 493624
rect 575688 493564 575828 493624
rect 575888 493564 576028 493624
rect 576088 493564 576228 493624
rect 576288 493564 576428 493624
rect 576488 493564 576628 493624
rect 576688 493564 576828 493624
rect 576888 493564 577028 493624
rect 577088 493564 577228 493624
rect 577288 493564 577428 493624
rect 577488 493564 577628 493624
rect 577688 493564 577828 493624
rect 577888 493564 578028 493624
rect 578088 493564 578228 493624
rect 578288 493564 578428 493624
rect 578488 493564 578628 493624
rect 578688 493564 578828 493624
rect 578888 493564 579028 493624
rect 579088 493564 579228 493624
rect 579288 493564 579428 493624
rect 579488 493564 579628 493624
rect 579688 493564 579828 493624
rect 579888 493564 580028 493624
rect 580088 493564 580228 493624
rect 580288 493564 580556 493624
rect 576720 493522 576880 493564
rect 576720 493486 576776 493522
rect 576820 493486 576880 493522
rect 576720 493484 576880 493486
rect 578020 493522 578180 493564
rect 578020 493486 578076 493522
rect 578120 493486 578180 493522
rect 578020 493484 578180 493486
rect 579320 493522 579480 493564
rect 579320 493486 579376 493522
rect 579420 493486 579480 493522
rect 579320 493484 579480 493486
rect 580468 493474 580528 493564
rect 574980 493444 575040 493446
rect 565563 492436 565597 492452
rect 565821 493428 565855 493444
rect 565821 492444 565855 492452
rect 574980 493404 580398 493444
rect 580468 493434 580478 493474
rect 580518 493434 580528 493474
rect 574980 493384 580396 493404
rect 565821 492424 565880 492444
rect 565821 492370 566074 492424
rect 560330 492312 560482 492332
rect 560388 492204 560482 492312
rect 560648 492320 566074 492370
rect 566234 492320 566240 492424
rect 560648 492310 566240 492320
rect 560388 492144 560836 492204
rect 560896 492144 561036 492204
rect 561096 492144 561236 492204
rect 561296 492144 561436 492204
rect 561496 492144 561636 492204
rect 561696 492144 561836 492204
rect 561896 492144 562036 492204
rect 562096 492144 562236 492204
rect 562296 492144 562436 492204
rect 562496 492144 562636 492204
rect 562696 492144 562836 492204
rect 562896 492144 563036 492204
rect 563096 492144 563236 492204
rect 563296 492144 563436 492204
rect 563496 492144 563636 492204
rect 563696 492144 563836 492204
rect 563896 492144 564036 492204
rect 564096 492144 564236 492204
rect 564296 492144 564436 492204
rect 564496 492144 564636 492204
rect 564696 492144 564836 492204
rect 564896 492144 565036 492204
rect 565096 492144 565236 492204
rect 565296 492144 565436 492204
rect 565496 492144 565636 492204
rect 565696 492144 565786 492204
rect 565876 492100 565936 492180
rect 562128 492068 562288 492090
rect 562128 492032 562184 492068
rect 562228 492032 562288 492068
rect 562128 491970 562288 492032
rect 563428 492068 563588 492090
rect 563428 492032 563484 492068
rect 563528 492032 563588 492068
rect 563428 491970 563588 492032
rect 564728 492068 564888 492090
rect 564728 492032 564784 492068
rect 564828 492032 564888 492068
rect 564728 491970 564888 492032
rect 565876 492060 565886 492100
rect 565926 492060 565936 492100
rect 565876 491970 565936 492060
rect 574980 492038 575040 493384
rect 575217 493202 575251 493218
rect 575217 492084 575251 492226
rect 575475 493202 575509 493384
rect 575475 492210 575509 492226
rect 575733 493202 575767 493218
rect 575733 492084 575767 492226
rect 575991 493202 576025 493384
rect 575991 492210 576025 492226
rect 576249 493202 576283 493218
rect 576249 492084 576283 492226
rect 576507 493202 576541 493384
rect 576507 492210 576541 492226
rect 576765 493202 576799 493218
rect 576765 492084 576799 492226
rect 577023 493202 577057 493384
rect 577023 492210 577057 492226
rect 577281 493202 577315 493218
rect 577281 492084 577315 492226
rect 577539 493202 577573 493384
rect 577539 492210 577573 492226
rect 577797 493202 577831 493218
rect 577797 492084 577831 492226
rect 578055 493202 578089 493384
rect 578055 492210 578089 492226
rect 578313 493202 578347 493218
rect 578313 492084 578347 492226
rect 578571 493202 578605 493384
rect 578571 492210 578605 492226
rect 578829 493202 578863 493218
rect 578829 492084 578863 492226
rect 579087 493202 579121 493384
rect 579087 492210 579121 492226
rect 579345 493202 579379 493218
rect 579345 492084 579379 492226
rect 579603 493202 579637 493384
rect 579603 492210 579637 492226
rect 579861 493202 579895 493218
rect 579861 492084 579895 492226
rect 580119 493202 580153 493384
rect 580468 493354 580528 493434
rect 580119 492210 580153 492226
rect 580377 493202 580411 493218
rect 580377 492128 580411 492226
rect 580377 492118 580642 492128
rect 580377 492084 580542 492118
rect 574924 491984 575040 492038
rect 575164 492030 580542 492084
rect 580632 492030 580642 492118
rect 575164 492024 580642 492030
rect 560650 491910 560836 491970
rect 560896 491910 561036 491970
rect 561096 491910 561236 491970
rect 561296 491910 561436 491970
rect 561496 491910 561636 491970
rect 561696 491910 561836 491970
rect 561896 491910 562036 491970
rect 562096 491910 562236 491970
rect 562296 491910 562436 491970
rect 562496 491910 562636 491970
rect 562696 491910 562836 491970
rect 562896 491910 563036 491970
rect 563096 491910 563236 491970
rect 563296 491910 563436 491970
rect 563496 491910 563636 491970
rect 563696 491910 563836 491970
rect 563896 491910 564036 491970
rect 564096 491910 564236 491970
rect 564296 491910 564436 491970
rect 564496 491910 564636 491970
rect 564696 491910 564836 491970
rect 564896 491910 565036 491970
rect 565096 491910 565236 491970
rect 565296 491910 565436 491970
rect 565496 491910 565636 491970
rect 565696 491910 565964 491970
rect 574924 491880 574934 491984
rect 575026 491922 575040 491984
rect 575026 491880 575228 491922
rect 574924 491864 575228 491880
rect 574962 491862 575228 491864
rect 575288 491862 575428 491922
rect 575488 491862 575628 491922
rect 575688 491862 575828 491922
rect 575888 491862 576028 491922
rect 576088 491862 576228 491922
rect 576288 491862 576428 491922
rect 576488 491862 576628 491922
rect 576688 491862 576828 491922
rect 576888 491862 577028 491922
rect 577088 491862 577228 491922
rect 577288 491862 577428 491922
rect 577488 491862 577628 491922
rect 577688 491862 577828 491922
rect 577888 491862 578028 491922
rect 578088 491862 578228 491922
rect 578288 491862 578428 491922
rect 578488 491862 578628 491922
rect 578688 491862 578828 491922
rect 578888 491862 579028 491922
rect 579088 491862 579228 491922
rect 579288 491862 579428 491922
rect 579488 491862 579628 491922
rect 579688 491862 579828 491922
rect 579888 491862 580028 491922
rect 580088 491862 580228 491922
rect 580288 491862 580458 491922
rect 575170 491684 575228 491744
rect 575288 491684 575428 491744
rect 575488 491684 575628 491744
rect 575688 491684 575828 491744
rect 575888 491684 576028 491744
rect 576088 491684 576228 491744
rect 576288 491684 576428 491744
rect 576488 491684 576628 491744
rect 576688 491684 576828 491744
rect 576888 491684 577028 491744
rect 577088 491684 577228 491744
rect 577288 491684 577428 491744
rect 577488 491684 577628 491744
rect 577688 491684 577828 491744
rect 577888 491684 578028 491744
rect 578088 491684 578228 491744
rect 578288 491684 578428 491744
rect 578488 491684 578628 491744
rect 578688 491684 578828 491744
rect 578888 491684 579028 491744
rect 579088 491684 579228 491744
rect 579288 491684 579428 491744
rect 579488 491684 579628 491744
rect 579688 491684 579828 491744
rect 579888 491684 580028 491744
rect 580088 491684 580228 491744
rect 580288 491684 580556 491744
rect 493078 408853 493138 409036
rect 493078 408819 493091 408853
rect 493125 408819 493138 408853
rect 493078 408453 493138 408819
rect 493078 408419 493091 408453
rect 493125 408419 493138 408453
rect 493078 408053 493138 408419
rect 493078 408019 493091 408053
rect 493125 408019 493138 408053
rect 493078 407653 493138 408019
rect 493078 407619 493091 407653
rect 493125 407619 493138 407653
rect 493078 407253 493138 407619
rect 493078 407219 493091 407253
rect 493125 407219 493138 407253
rect 493078 406853 493138 407219
rect 493078 406819 493091 406853
rect 493125 406819 493138 406853
rect 493078 406453 493138 406819
rect 493078 406419 493091 406453
rect 493125 406419 493138 406453
rect 493078 406053 493138 406419
rect 493078 406019 493091 406053
rect 493125 406019 493138 406053
rect 493078 405653 493138 406019
rect 493078 405619 493091 405653
rect 493125 405619 493138 405653
rect 493078 405253 493138 405619
rect 493078 405219 493091 405253
rect 493125 405219 493138 405253
rect 493078 404853 493138 405219
rect 493078 404819 493091 404853
rect 493125 404819 493138 404853
rect 493078 404453 493138 404819
rect 493078 404419 493091 404453
rect 493125 404419 493138 404453
rect 493078 404053 493138 404419
rect 493078 404019 493091 404053
rect 493125 404019 493138 404053
rect 493078 403653 493138 404019
rect 493078 403619 493091 403653
rect 493125 403619 493138 403653
rect 493078 403253 493138 403619
rect 493078 403219 493091 403253
rect 493125 403219 493138 403253
rect 493078 402853 493138 403219
rect 493078 402819 493091 402853
rect 493125 402819 493138 402853
rect 493078 402453 493138 402819
rect 493078 402419 493091 402453
rect 493125 402419 493138 402453
rect 493078 402053 493138 402419
rect 493078 402019 493091 402053
rect 493125 402019 493138 402053
rect 493078 401868 493138 402019
rect 494958 408853 495018 409036
rect 494958 408819 494971 408853
rect 495005 408819 495018 408853
rect 494958 408453 495018 408819
rect 494958 408419 494971 408453
rect 495005 408419 495018 408453
rect 494958 408053 495018 408419
rect 494958 408019 494971 408053
rect 495005 408019 495018 408053
rect 494958 407653 495018 408019
rect 494958 407619 494971 407653
rect 495005 407619 495018 407653
rect 494958 407253 495018 407619
rect 494958 407219 494971 407253
rect 495005 407219 495018 407253
rect 494958 406853 495018 407219
rect 494958 406819 494971 406853
rect 495005 406819 495018 406853
rect 494958 406453 495018 406819
rect 494958 406419 494971 406453
rect 495005 406419 495018 406453
rect 494958 406053 495018 406419
rect 494958 406019 494971 406053
rect 495005 406019 495018 406053
rect 494958 405653 495018 406019
rect 494958 405619 494971 405653
rect 495005 405619 495018 405653
rect 494958 405253 495018 405619
rect 494958 405219 494971 405253
rect 495005 405219 495018 405253
rect 494958 404853 495018 405219
rect 494958 404819 494971 404853
rect 495005 404819 495018 404853
rect 494958 404453 495018 404819
rect 494958 404419 494971 404453
rect 495005 404419 495018 404453
rect 494958 404053 495018 404419
rect 494958 404019 494971 404053
rect 495005 404019 495018 404053
rect 494958 403653 495018 404019
rect 494958 403619 494971 403653
rect 495005 403619 495018 403653
rect 494958 403253 495018 403619
rect 494958 403219 494971 403253
rect 495005 403219 495018 403253
rect 494958 402853 495018 403219
rect 494958 402819 494971 402853
rect 495005 402819 495018 402853
rect 494958 402453 495018 402819
rect 494958 402419 494971 402453
rect 495005 402419 495018 402453
rect 494958 402053 495018 402419
rect 494958 402019 494971 402053
rect 495005 402019 495018 402053
rect 494958 401868 495018 402019
rect 496838 408853 496898 409036
rect 496838 408819 496851 408853
rect 496885 408819 496898 408853
rect 496838 408453 496898 408819
rect 496838 408419 496851 408453
rect 496885 408419 496898 408453
rect 496838 408053 496898 408419
rect 496838 408019 496851 408053
rect 496885 408019 496898 408053
rect 496838 407653 496898 408019
rect 496838 407619 496851 407653
rect 496885 407619 496898 407653
rect 496838 407253 496898 407619
rect 496838 407219 496851 407253
rect 496885 407219 496898 407253
rect 496838 406853 496898 407219
rect 496838 406819 496851 406853
rect 496885 406819 496898 406853
rect 496838 406453 496898 406819
rect 496838 406419 496851 406453
rect 496885 406419 496898 406453
rect 496838 406053 496898 406419
rect 496838 406019 496851 406053
rect 496885 406019 496898 406053
rect 496838 405653 496898 406019
rect 496838 405619 496851 405653
rect 496885 405619 496898 405653
rect 496838 405253 496898 405619
rect 496838 405219 496851 405253
rect 496885 405219 496898 405253
rect 496838 404853 496898 405219
rect 496838 404819 496851 404853
rect 496885 404819 496898 404853
rect 496838 404453 496898 404819
rect 496838 404419 496851 404453
rect 496885 404419 496898 404453
rect 496838 404053 496898 404419
rect 496838 404019 496851 404053
rect 496885 404019 496898 404053
rect 496838 403653 496898 404019
rect 496838 403619 496851 403653
rect 496885 403619 496898 403653
rect 496838 403253 496898 403619
rect 496838 403219 496851 403253
rect 496885 403219 496898 403253
rect 496838 402853 496898 403219
rect 496838 402819 496851 402853
rect 496885 402819 496898 402853
rect 496838 402453 496898 402819
rect 496838 402419 496851 402453
rect 496885 402419 496898 402453
rect 496838 402053 496898 402419
rect 496838 402019 496851 402053
rect 496885 402019 496898 402053
rect 496838 401868 496898 402019
rect 498718 408853 498778 409036
rect 498718 408819 498731 408853
rect 498765 408819 498778 408853
rect 498718 408453 498778 408819
rect 498718 408419 498731 408453
rect 498765 408419 498778 408453
rect 498718 408053 498778 408419
rect 498718 408019 498731 408053
rect 498765 408019 498778 408053
rect 498718 407653 498778 408019
rect 498718 407619 498731 407653
rect 498765 407619 498778 407653
rect 498718 407253 498778 407619
rect 498718 407219 498731 407253
rect 498765 407219 498778 407253
rect 498718 406853 498778 407219
rect 498718 406819 498731 406853
rect 498765 406819 498778 406853
rect 498718 406453 498778 406819
rect 498718 406419 498731 406453
rect 498765 406419 498778 406453
rect 498718 406053 498778 406419
rect 498718 406019 498731 406053
rect 498765 406019 498778 406053
rect 498718 405653 498778 406019
rect 498718 405619 498731 405653
rect 498765 405619 498778 405653
rect 498718 405253 498778 405619
rect 498718 405219 498731 405253
rect 498765 405219 498778 405253
rect 498718 404853 498778 405219
rect 498718 404819 498731 404853
rect 498765 404819 498778 404853
rect 498718 404453 498778 404819
rect 498718 404419 498731 404453
rect 498765 404419 498778 404453
rect 498718 404053 498778 404419
rect 498718 404019 498731 404053
rect 498765 404019 498778 404053
rect 498718 403653 498778 404019
rect 498718 403619 498731 403653
rect 498765 403619 498778 403653
rect 498718 403253 498778 403619
rect 498718 403219 498731 403253
rect 498765 403219 498778 403253
rect 498718 402853 498778 403219
rect 498718 402819 498731 402853
rect 498765 402819 498778 402853
rect 498718 402453 498778 402819
rect 498718 402419 498731 402453
rect 498765 402419 498778 402453
rect 498718 402053 498778 402419
rect 498718 402019 498731 402053
rect 498765 402019 498778 402053
rect 498718 401868 498778 402019
rect 500598 408461 500658 408644
rect 500598 408427 500611 408461
rect 500645 408427 500658 408461
rect 500598 408061 500658 408427
rect 500598 408027 500611 408061
rect 500645 408027 500658 408061
rect 500598 407661 500658 408027
rect 500598 407627 500611 407661
rect 500645 407627 500658 407661
rect 500598 407261 500658 407627
rect 500598 407227 500611 407261
rect 500645 407227 500658 407261
rect 500598 406861 500658 407227
rect 500598 406827 500611 406861
rect 500645 406827 500658 406861
rect 500598 406461 500658 406827
rect 500598 406427 500611 406461
rect 500645 406427 500658 406461
rect 500598 406061 500658 406427
rect 500598 406027 500611 406061
rect 500645 406027 500658 406061
rect 500598 405661 500658 406027
rect 500598 405627 500611 405661
rect 500645 405627 500658 405661
rect 500598 405261 500658 405627
rect 500598 405227 500611 405261
rect 500645 405227 500658 405261
rect 500598 404861 500658 405227
rect 500598 404827 500611 404861
rect 500645 404827 500658 404861
rect 500598 404461 500658 404827
rect 500598 404427 500611 404461
rect 500645 404427 500658 404461
rect 500598 404061 500658 404427
rect 500598 404027 500611 404061
rect 500645 404027 500658 404061
rect 500598 403661 500658 404027
rect 500598 403627 500611 403661
rect 500645 403627 500658 403661
rect 500598 403261 500658 403627
rect 500598 403227 500611 403261
rect 500645 403227 500658 403261
rect 500598 402861 500658 403227
rect 500598 402827 500611 402861
rect 500645 402827 500658 402861
rect 500598 402461 500658 402827
rect 500598 402427 500611 402461
rect 500645 402427 500658 402461
rect 500598 402061 500658 402427
rect 500598 402027 500611 402061
rect 500645 402027 500658 402061
rect 500598 401661 500658 402027
rect 500598 401627 500611 401661
rect 500645 401627 500658 401661
rect 493078 401405 493138 401588
rect 493078 401371 493091 401405
rect 493125 401371 493138 401405
rect 493078 401005 493138 401371
rect 493078 400971 493091 401005
rect 493125 400971 493138 401005
rect 493078 400605 493138 400971
rect 493078 400571 493091 400605
rect 493125 400571 493138 400605
rect 493078 400205 493138 400571
rect 493078 400171 493091 400205
rect 493125 400171 493138 400205
rect 493078 399805 493138 400171
rect 493078 399771 493091 399805
rect 493125 399771 493138 399805
rect 493078 399405 493138 399771
rect 493078 399371 493091 399405
rect 493125 399371 493138 399405
rect 493078 399005 493138 399371
rect 493078 398971 493091 399005
rect 493125 398971 493138 399005
rect 493078 398605 493138 398971
rect 493078 398571 493091 398605
rect 493125 398571 493138 398605
rect 493078 398205 493138 398571
rect 493078 398171 493091 398205
rect 493125 398171 493138 398205
rect 493078 397805 493138 398171
rect 493078 397771 493091 397805
rect 493125 397771 493138 397805
rect 493078 397405 493138 397771
rect 493078 397371 493091 397405
rect 493125 397371 493138 397405
rect 493078 397005 493138 397371
rect 493078 396971 493091 397005
rect 493125 396971 493138 397005
rect 493078 396605 493138 396971
rect 493078 396571 493091 396605
rect 493125 396571 493138 396605
rect 493078 396205 493138 396571
rect 493078 396171 493091 396205
rect 493125 396171 493138 396205
rect 493078 395805 493138 396171
rect 493078 395771 493091 395805
rect 493125 395771 493138 395805
rect 493078 395405 493138 395771
rect 493078 395371 493091 395405
rect 493125 395371 493138 395405
rect 493078 395005 493138 395371
rect 493078 394971 493091 395005
rect 493125 394971 493138 395005
rect 493078 394605 493138 394971
rect 493078 394571 493091 394605
rect 493125 394571 493138 394605
rect 493078 394420 493138 394571
rect 494958 401405 495018 401588
rect 500598 401476 500658 401627
rect 502478 408461 502538 408644
rect 502478 408427 502491 408461
rect 502525 408427 502538 408461
rect 502478 408061 502538 408427
rect 502478 408027 502491 408061
rect 502525 408027 502538 408061
rect 502478 407661 502538 408027
rect 502478 407627 502491 407661
rect 502525 407627 502538 407661
rect 502478 407261 502538 407627
rect 502478 407227 502491 407261
rect 502525 407227 502538 407261
rect 502478 406861 502538 407227
rect 502478 406827 502491 406861
rect 502525 406827 502538 406861
rect 502478 406461 502538 406827
rect 502478 406427 502491 406461
rect 502525 406427 502538 406461
rect 502478 406061 502538 406427
rect 502478 406027 502491 406061
rect 502525 406027 502538 406061
rect 502478 405661 502538 406027
rect 502478 405627 502491 405661
rect 502525 405627 502538 405661
rect 502478 405261 502538 405627
rect 502478 405227 502491 405261
rect 502525 405227 502538 405261
rect 502478 404861 502538 405227
rect 502478 404827 502491 404861
rect 502525 404827 502538 404861
rect 502478 404461 502538 404827
rect 560592 404648 560860 404708
rect 560920 404648 561060 404708
rect 561120 404648 561260 404708
rect 561320 404648 561460 404708
rect 561520 404648 561660 404708
rect 561720 404648 561860 404708
rect 561920 404648 562060 404708
rect 562120 404648 562260 404708
rect 562320 404648 562460 404708
rect 562520 404648 562660 404708
rect 562720 404648 562860 404708
rect 562920 404648 563060 404708
rect 563120 404648 563260 404708
rect 563320 404648 563460 404708
rect 563520 404648 563660 404708
rect 563720 404648 563860 404708
rect 563920 404648 564060 404708
rect 564120 404648 564260 404708
rect 564320 404648 564460 404708
rect 564520 404648 564660 404708
rect 564720 404648 564860 404708
rect 564920 404648 565060 404708
rect 565120 404648 565260 404708
rect 565320 404648 565460 404708
rect 565520 404648 565660 404708
rect 565720 404648 565906 404708
rect 574448 404688 574506 404748
rect 574566 404688 574706 404748
rect 574766 404688 574906 404748
rect 574966 404688 575106 404748
rect 575166 404688 575306 404748
rect 575366 404688 575506 404748
rect 575566 404688 575706 404748
rect 575766 404688 575906 404748
rect 575966 404688 576106 404748
rect 576166 404688 576306 404748
rect 576366 404688 576506 404748
rect 576566 404688 576706 404748
rect 576766 404688 576906 404748
rect 576966 404688 577106 404748
rect 577166 404688 577306 404748
rect 577366 404688 577506 404748
rect 577566 404688 577706 404748
rect 577766 404688 577906 404748
rect 577966 404688 578106 404748
rect 578166 404688 578306 404748
rect 578366 404688 578506 404748
rect 578566 404688 578706 404748
rect 578766 404688 578906 404748
rect 578966 404688 579106 404748
rect 579166 404688 579306 404748
rect 579366 404688 579506 404748
rect 579566 404688 579834 404748
rect 575998 404646 576158 404688
rect 575998 404610 576054 404646
rect 576098 404610 576158 404646
rect 575998 404608 576158 404610
rect 577298 404646 577458 404688
rect 577298 404610 577354 404646
rect 577398 404610 577458 404646
rect 577298 404608 577458 404610
rect 578598 404646 578758 404688
rect 578598 404610 578654 404646
rect 578698 404610 578758 404646
rect 578598 404608 578758 404610
rect 579746 404598 579806 404688
rect 574258 404568 574318 404570
rect 566108 404548 566168 404550
rect 560690 404488 566168 404548
rect 502478 404427 502491 404461
rect 502525 404427 502538 404461
rect 502478 404061 502538 404427
rect 502478 404027 502491 404061
rect 502525 404027 502538 404061
rect 502478 403661 502538 404027
rect 502478 403627 502491 403661
rect 502525 403627 502538 403661
rect 502478 403261 502538 403627
rect 560701 404286 560735 404302
rect 560701 403302 560735 403310
rect 502478 403227 502491 403261
rect 502525 403227 502538 403261
rect 502478 402861 502538 403227
rect 560316 403178 560322 403282
rect 560676 403282 560735 403302
rect 560959 404286 560993 404488
rect 560959 403294 560993 403310
rect 561217 404286 561251 404302
rect 560482 403228 560735 403282
rect 561217 403228 561251 403310
rect 561475 404286 561509 404488
rect 561475 403294 561509 403310
rect 561733 404286 561767 404302
rect 561733 403228 561767 403310
rect 561991 404286 562025 404488
rect 561991 403294 562025 403310
rect 562249 404286 562283 404302
rect 562249 403228 562283 403310
rect 562507 404286 562541 404488
rect 562507 403294 562541 403310
rect 562765 404286 562799 404302
rect 562765 403228 562799 403310
rect 563023 404286 563057 404488
rect 563023 403294 563057 403310
rect 563281 404286 563315 404302
rect 563281 403228 563315 403310
rect 563539 404286 563573 404488
rect 563539 403294 563573 403310
rect 563797 404286 563831 404302
rect 563797 403228 563831 403310
rect 564055 404286 564089 404488
rect 564055 403294 564089 403310
rect 564313 404286 564347 404302
rect 564313 403228 564347 403310
rect 564571 404286 564605 404488
rect 564571 403294 564605 403310
rect 564829 404286 564863 404302
rect 564829 403228 564863 403310
rect 565087 404286 565121 404488
rect 565087 403294 565121 403310
rect 565345 404286 565379 404302
rect 565345 403228 565379 403310
rect 565603 404286 565637 404488
rect 565603 403294 565637 403310
rect 565861 404286 565895 404302
rect 565861 403294 565895 403310
rect 566074 403380 566168 404488
rect 574258 404528 579676 404568
rect 579746 404558 579756 404598
rect 579796 404558 579806 404598
rect 574258 404508 579674 404528
rect 566074 403362 566214 403380
rect 566074 403340 566226 403362
rect 560482 403178 565908 403228
rect 560316 403168 565908 403178
rect 566074 403190 566084 403340
rect 566216 403190 566226 403340
rect 566074 403170 566226 403190
rect 566074 403062 566168 403170
rect 574258 403162 574318 404508
rect 574495 404326 574529 404342
rect 574495 403208 574529 403350
rect 574753 404326 574787 404508
rect 574753 403334 574787 403350
rect 575011 404326 575045 404342
rect 575011 403208 575045 403350
rect 575269 404326 575303 404508
rect 575269 403334 575303 403350
rect 575527 404326 575561 404342
rect 575527 403208 575561 403350
rect 575785 404326 575819 404508
rect 575785 403334 575819 403350
rect 576043 404326 576077 404342
rect 576043 403208 576077 403350
rect 576301 404326 576335 404508
rect 576301 403334 576335 403350
rect 576559 404326 576593 404342
rect 576559 403208 576593 403350
rect 576817 404326 576851 404508
rect 576817 403334 576851 403350
rect 577075 404326 577109 404342
rect 577075 403208 577109 403350
rect 577333 404326 577367 404508
rect 577333 403334 577367 403350
rect 577591 404326 577625 404342
rect 577591 403208 577625 403350
rect 577849 404326 577883 404508
rect 577849 403334 577883 403350
rect 578107 404326 578141 404342
rect 578107 403208 578141 403350
rect 578365 404326 578399 404508
rect 578365 403334 578399 403350
rect 578623 404326 578657 404342
rect 578623 403208 578657 403350
rect 578881 404326 578915 404508
rect 578881 403334 578915 403350
rect 579139 404326 579173 404342
rect 579139 403208 579173 403350
rect 579397 404326 579431 404508
rect 579746 404478 579806 404558
rect 579397 403334 579431 403350
rect 579655 404326 579689 404342
rect 579655 403252 579689 403350
rect 579655 403242 579920 403252
rect 579655 403208 579820 403242
rect 502478 402827 502491 402861
rect 502525 402827 502538 402861
rect 502478 402461 502538 402827
rect 502478 402427 502491 402461
rect 502525 402427 502538 402461
rect 502478 402061 502538 402427
rect 502478 402027 502491 402061
rect 502525 402027 502538 402061
rect 502478 401661 502538 402027
rect 502478 401627 502491 401661
rect 502525 401627 502538 401661
rect 502478 401476 502538 401627
rect 504358 402779 504418 402962
rect 504358 402745 504371 402779
rect 504405 402745 504418 402779
rect 504358 402579 504418 402745
rect 504358 402545 504371 402579
rect 504405 402545 504418 402579
rect 504358 402379 504418 402545
rect 504358 402345 504371 402379
rect 504405 402345 504418 402379
rect 504358 402179 504418 402345
rect 504358 402145 504371 402179
rect 504405 402145 504418 402179
rect 504358 401979 504418 402145
rect 504358 401945 504371 401979
rect 504405 401945 504418 401979
rect 504358 401779 504418 401945
rect 504358 401745 504371 401779
rect 504405 401745 504418 401779
rect 504358 401622 504418 401745
rect 504684 402902 505972 402936
rect 504684 402868 504742 402902
rect 504776 402868 504832 402902
rect 504866 402868 504922 402902
rect 504956 402868 505012 402902
rect 505046 402868 505102 402902
rect 505136 402868 505192 402902
rect 505226 402868 505282 402902
rect 505316 402868 505372 402902
rect 505406 402868 505462 402902
rect 505496 402868 505552 402902
rect 505586 402868 505642 402902
rect 505676 402868 505732 402902
rect 505766 402868 505822 402902
rect 505856 402868 505972 402902
rect 504684 402837 505972 402868
rect 504684 402806 504783 402837
rect 504684 402772 504719 402806
rect 504753 402772 504783 402806
rect 505873 402806 505972 402837
rect 504684 402716 504783 402772
rect 504684 402682 504719 402716
rect 504753 402682 504783 402716
rect 504684 402626 504783 402682
rect 504684 402592 504719 402626
rect 504753 402592 504783 402626
rect 504684 402536 504783 402592
rect 504684 402502 504719 402536
rect 504753 402502 504783 402536
rect 504684 402446 504783 402502
rect 504684 402412 504719 402446
rect 504753 402412 504783 402446
rect 504684 402356 504783 402412
rect 504684 402322 504719 402356
rect 504753 402322 504783 402356
rect 504684 402266 504783 402322
rect 504684 402232 504719 402266
rect 504753 402232 504783 402266
rect 504684 402176 504783 402232
rect 504684 402142 504719 402176
rect 504753 402142 504783 402176
rect 504684 402086 504783 402142
rect 504684 402052 504719 402086
rect 504753 402052 504783 402086
rect 504684 401996 504783 402052
rect 504684 401962 504719 401996
rect 504753 401962 504783 401996
rect 504684 401906 504783 401962
rect 504684 401872 504719 401906
rect 504753 401872 504783 401906
rect 504684 401816 504783 401872
rect 504684 401782 504719 401816
rect 504753 401782 504783 401816
rect 504847 402754 505809 402773
rect 504847 402720 504923 402754
rect 504957 402720 505013 402754
rect 505047 402720 505103 402754
rect 505137 402720 505193 402754
rect 505227 402720 505283 402754
rect 505317 402720 505373 402754
rect 505407 402720 505463 402754
rect 505497 402720 505553 402754
rect 505587 402720 505643 402754
rect 505677 402720 505809 402754
rect 504847 402701 505809 402720
rect 504847 402642 504919 402701
rect 504847 402608 504866 402642
rect 504900 402608 504919 402642
rect 505737 402676 505809 402701
rect 505737 402642 505756 402676
rect 505790 402642 505809 402676
rect 504847 402552 504919 402608
rect 504847 402518 504866 402552
rect 504900 402518 504919 402552
rect 504847 402462 504919 402518
rect 504847 402428 504866 402462
rect 504900 402428 504919 402462
rect 504847 402372 504919 402428
rect 504847 402338 504866 402372
rect 504900 402338 504919 402372
rect 504847 402282 504919 402338
rect 504847 402248 504866 402282
rect 504900 402248 504919 402282
rect 504847 402192 504919 402248
rect 504847 402158 504866 402192
rect 504900 402158 504919 402192
rect 504847 402102 504919 402158
rect 504847 402068 504866 402102
rect 504900 402068 504919 402102
rect 504847 402012 504919 402068
rect 504847 401978 504866 402012
rect 504900 401978 504919 402012
rect 504847 401922 504919 401978
rect 504981 402578 505675 402639
rect 504981 402544 505040 402578
rect 505074 402566 505130 402578
rect 505102 402544 505130 402566
rect 505164 402566 505220 402578
rect 505164 402544 505168 402566
rect 504981 402532 505068 402544
rect 505102 402532 505168 402544
rect 505202 402544 505220 402566
rect 505254 402566 505310 402578
rect 505254 402544 505268 402566
rect 505202 402532 505268 402544
rect 505302 402544 505310 402566
rect 505344 402566 505400 402578
rect 505434 402566 505490 402578
rect 505524 402566 505580 402578
rect 505344 402544 505368 402566
rect 505434 402544 505468 402566
rect 505524 402544 505568 402566
rect 505614 402544 505675 402578
rect 505302 402532 505368 402544
rect 505402 402532 505468 402544
rect 505502 402532 505568 402544
rect 505602 402532 505675 402544
rect 504981 402488 505675 402532
rect 504981 402454 505040 402488
rect 505074 402466 505130 402488
rect 505102 402454 505130 402466
rect 505164 402466 505220 402488
rect 505164 402454 505168 402466
rect 504981 402432 505068 402454
rect 505102 402432 505168 402454
rect 505202 402454 505220 402466
rect 505254 402466 505310 402488
rect 505254 402454 505268 402466
rect 505202 402432 505268 402454
rect 505302 402454 505310 402466
rect 505344 402466 505400 402488
rect 505434 402466 505490 402488
rect 505524 402466 505580 402488
rect 505344 402454 505368 402466
rect 505434 402454 505468 402466
rect 505524 402454 505568 402466
rect 505614 402454 505675 402488
rect 505302 402432 505368 402454
rect 505402 402432 505468 402454
rect 505502 402432 505568 402454
rect 505602 402432 505675 402454
rect 504981 402398 505675 402432
rect 504981 402364 505040 402398
rect 505074 402366 505130 402398
rect 505102 402364 505130 402366
rect 505164 402366 505220 402398
rect 505164 402364 505168 402366
rect 504981 402332 505068 402364
rect 505102 402332 505168 402364
rect 505202 402364 505220 402366
rect 505254 402366 505310 402398
rect 505254 402364 505268 402366
rect 505202 402332 505268 402364
rect 505302 402364 505310 402366
rect 505344 402366 505400 402398
rect 505434 402366 505490 402398
rect 505524 402366 505580 402398
rect 505344 402364 505368 402366
rect 505434 402364 505468 402366
rect 505524 402364 505568 402366
rect 505614 402364 505675 402398
rect 505302 402332 505368 402364
rect 505402 402332 505468 402364
rect 505502 402332 505568 402364
rect 505602 402332 505675 402364
rect 504981 402308 505675 402332
rect 504981 402274 505040 402308
rect 505074 402274 505130 402308
rect 505164 402274 505220 402308
rect 505254 402274 505310 402308
rect 505344 402274 505400 402308
rect 505434 402274 505490 402308
rect 505524 402274 505580 402308
rect 505614 402274 505675 402308
rect 504981 402266 505675 402274
rect 504981 402232 505068 402266
rect 505102 402232 505168 402266
rect 505202 402232 505268 402266
rect 505302 402232 505368 402266
rect 505402 402232 505468 402266
rect 505502 402232 505568 402266
rect 505602 402232 505675 402266
rect 504981 402218 505675 402232
rect 504981 402184 505040 402218
rect 505074 402184 505130 402218
rect 505164 402184 505220 402218
rect 505254 402184 505310 402218
rect 505344 402184 505400 402218
rect 505434 402184 505490 402218
rect 505524 402184 505580 402218
rect 505614 402184 505675 402218
rect 504981 402166 505675 402184
rect 504981 402132 505068 402166
rect 505102 402132 505168 402166
rect 505202 402132 505268 402166
rect 505302 402132 505368 402166
rect 505402 402132 505468 402166
rect 505502 402132 505568 402166
rect 505602 402132 505675 402166
rect 504981 402128 505675 402132
rect 504981 402094 505040 402128
rect 505074 402094 505130 402128
rect 505164 402094 505220 402128
rect 505254 402094 505310 402128
rect 505344 402094 505400 402128
rect 505434 402094 505490 402128
rect 505524 402094 505580 402128
rect 505614 402094 505675 402128
rect 504981 402066 505675 402094
rect 504981 402038 505068 402066
rect 505102 402038 505168 402066
rect 504981 402004 505040 402038
rect 505102 402032 505130 402038
rect 505074 402004 505130 402032
rect 505164 402032 505168 402038
rect 505202 402038 505268 402066
rect 505202 402032 505220 402038
rect 505164 402004 505220 402032
rect 505254 402032 505268 402038
rect 505302 402038 505368 402066
rect 505402 402038 505468 402066
rect 505502 402038 505568 402066
rect 505602 402038 505675 402066
rect 505302 402032 505310 402038
rect 505254 402004 505310 402032
rect 505344 402032 505368 402038
rect 505434 402032 505468 402038
rect 505524 402032 505568 402038
rect 505344 402004 505400 402032
rect 505434 402004 505490 402032
rect 505524 402004 505580 402032
rect 505614 402004 505675 402038
rect 504981 401945 505675 402004
rect 505737 402586 505809 402642
rect 505737 402552 505756 402586
rect 505790 402552 505809 402586
rect 505737 402496 505809 402552
rect 505737 402462 505756 402496
rect 505790 402462 505809 402496
rect 505737 402406 505809 402462
rect 505737 402372 505756 402406
rect 505790 402372 505809 402406
rect 505737 402316 505809 402372
rect 505737 402282 505756 402316
rect 505790 402282 505809 402316
rect 505737 402226 505809 402282
rect 505737 402192 505756 402226
rect 505790 402192 505809 402226
rect 505737 402136 505809 402192
rect 505737 402102 505756 402136
rect 505790 402102 505809 402136
rect 505737 402046 505809 402102
rect 505737 402012 505756 402046
rect 505790 402012 505809 402046
rect 505737 401956 505809 402012
rect 504847 401888 504866 401922
rect 504900 401888 504919 401922
rect 504847 401883 504919 401888
rect 505737 401922 505756 401956
rect 505790 401922 505809 401956
rect 505737 401883 505809 401922
rect 504847 401864 505809 401883
rect 504847 401830 504942 401864
rect 504976 401830 505032 401864
rect 505066 401830 505122 401864
rect 505156 401830 505212 401864
rect 505246 401830 505302 401864
rect 505336 401830 505392 401864
rect 505426 401830 505482 401864
rect 505516 401830 505572 401864
rect 505606 401830 505662 401864
rect 505696 401861 505809 401864
rect 505696 401830 505765 401861
rect 504847 401827 505765 401830
rect 505799 401827 505809 401861
rect 504847 401811 505809 401827
rect 505873 402772 505906 402806
rect 505940 402772 505972 402806
rect 505873 402716 505972 402772
rect 505873 402682 505906 402716
rect 505940 402682 505972 402716
rect 505873 402626 505972 402682
rect 505873 402592 505906 402626
rect 505940 402592 505972 402626
rect 505873 402536 505972 402592
rect 505873 402502 505906 402536
rect 505940 402502 505972 402536
rect 505873 402446 505972 402502
rect 505873 402412 505906 402446
rect 505940 402412 505972 402446
rect 505873 402356 505972 402412
rect 505873 402322 505906 402356
rect 505940 402322 505972 402356
rect 505873 402266 505972 402322
rect 505873 402232 505906 402266
rect 505940 402232 505972 402266
rect 505873 402176 505972 402232
rect 505873 402142 505906 402176
rect 505940 402142 505972 402176
rect 505873 402086 505972 402142
rect 505873 402052 505906 402086
rect 505940 402052 505972 402086
rect 505873 401996 505972 402052
rect 505873 401962 505906 401996
rect 505940 401962 505972 401996
rect 505873 401906 505972 401962
rect 505873 401872 505906 401906
rect 505940 401872 505972 401906
rect 505873 401816 505972 401872
rect 504684 401747 504783 401782
rect 505873 401782 505906 401816
rect 505940 401782 505972 401816
rect 505873 401747 505972 401782
rect 504684 401715 505972 401747
rect 504684 401681 504742 401715
rect 504776 401681 504832 401715
rect 504866 401681 504922 401715
rect 504956 401681 505012 401715
rect 505046 401681 505102 401715
rect 505136 401681 505192 401715
rect 505226 401681 505282 401715
rect 505316 401681 505372 401715
rect 505406 401681 505462 401715
rect 505496 401681 505552 401715
rect 505586 401681 505642 401715
rect 505676 401681 505732 401715
rect 505766 401681 505822 401715
rect 505856 401681 505972 401715
rect 504684 401677 505972 401681
rect 504684 401648 505901 401677
rect 505935 401648 505972 401677
rect 506238 402779 506298 402962
rect 560620 402958 560680 403038
rect 560770 403002 560860 403062
rect 560920 403002 561060 403062
rect 561120 403002 561260 403062
rect 561320 403002 561460 403062
rect 561520 403002 561660 403062
rect 561720 403002 561860 403062
rect 561920 403002 562060 403062
rect 562120 403002 562260 403062
rect 562320 403002 562460 403062
rect 562520 403002 562660 403062
rect 562720 403002 562860 403062
rect 562920 403002 563060 403062
rect 563120 403002 563260 403062
rect 563320 403002 563460 403062
rect 563520 403002 563660 403062
rect 563720 403002 563860 403062
rect 563920 403002 564060 403062
rect 564120 403002 564260 403062
rect 564320 403002 564460 403062
rect 564520 403002 564660 403062
rect 564720 403002 564860 403062
rect 564920 403002 565060 403062
rect 565120 403002 565260 403062
rect 565320 403002 565460 403062
rect 565520 403002 565660 403062
rect 565720 403002 566168 403062
rect 574202 403108 574318 403162
rect 574442 403154 579820 403208
rect 579910 403154 579920 403242
rect 574442 403148 579920 403154
rect 574202 403004 574212 403108
rect 574304 403046 574318 403108
rect 574304 403004 574506 403046
rect 574202 402988 574506 403004
rect 574240 402986 574506 402988
rect 574566 402986 574706 403046
rect 574766 402986 574906 403046
rect 574966 402986 575106 403046
rect 575166 402986 575306 403046
rect 575366 402986 575506 403046
rect 575566 402986 575706 403046
rect 575766 402986 575906 403046
rect 575966 402986 576106 403046
rect 576166 402986 576306 403046
rect 576366 402986 576506 403046
rect 576566 402986 576706 403046
rect 576766 402986 576906 403046
rect 576966 402986 577106 403046
rect 577166 402986 577306 403046
rect 577366 402986 577506 403046
rect 577566 402986 577706 403046
rect 577766 402986 577906 403046
rect 577966 402986 578106 403046
rect 578166 402986 578306 403046
rect 578366 402986 578506 403046
rect 578566 402986 578706 403046
rect 578766 402986 578906 403046
rect 578966 402986 579106 403046
rect 579166 402986 579306 403046
rect 579366 402986 579506 403046
rect 579566 402986 579736 403046
rect 560620 402918 560630 402958
rect 560670 402918 560680 402958
rect 560620 402828 560680 402918
rect 561668 402926 561828 402948
rect 561668 402890 561728 402926
rect 561772 402890 561828 402926
rect 561668 402828 561828 402890
rect 562968 402926 563128 402948
rect 562968 402890 563028 402926
rect 563072 402890 563128 402926
rect 562968 402828 563128 402890
rect 564268 402926 564428 402948
rect 564268 402890 564328 402926
rect 564372 402890 564428 402926
rect 564268 402828 564428 402890
rect 506238 402745 506251 402779
rect 506285 402745 506298 402779
rect 560592 402768 560860 402828
rect 560920 402768 561060 402828
rect 561120 402768 561260 402828
rect 561320 402768 561460 402828
rect 561520 402768 561660 402828
rect 561720 402768 561860 402828
rect 561920 402768 562060 402828
rect 562120 402768 562260 402828
rect 562320 402768 562460 402828
rect 562520 402768 562660 402828
rect 562720 402768 562860 402828
rect 562920 402768 563060 402828
rect 563120 402768 563260 402828
rect 563320 402768 563460 402828
rect 563520 402768 563660 402828
rect 563720 402768 563860 402828
rect 563920 402768 564060 402828
rect 564120 402768 564260 402828
rect 564320 402768 564460 402828
rect 564520 402768 564660 402828
rect 564720 402768 564860 402828
rect 564920 402768 565060 402828
rect 565120 402768 565260 402828
rect 565320 402768 565460 402828
rect 565520 402768 565660 402828
rect 565720 402768 565906 402828
rect 574448 402808 574506 402868
rect 574566 402808 574706 402868
rect 574766 402808 574906 402868
rect 574966 402808 575106 402868
rect 575166 402808 575306 402868
rect 575366 402808 575506 402868
rect 575566 402808 575706 402868
rect 575766 402808 575906 402868
rect 575966 402808 576106 402868
rect 576166 402808 576306 402868
rect 576366 402808 576506 402868
rect 576566 402808 576706 402868
rect 576766 402808 576906 402868
rect 576966 402808 577106 402868
rect 577166 402808 577306 402868
rect 577366 402808 577506 402868
rect 577566 402808 577706 402868
rect 577766 402808 577906 402868
rect 577966 402808 578106 402868
rect 578166 402808 578306 402868
rect 578366 402808 578506 402868
rect 578566 402808 578706 402868
rect 578766 402808 578906 402868
rect 578966 402808 579106 402868
rect 579166 402808 579306 402868
rect 579366 402808 579506 402868
rect 579566 402808 579834 402868
rect 506238 402579 506298 402745
rect 506238 402545 506251 402579
rect 506285 402545 506298 402579
rect 506238 402379 506298 402545
rect 506238 402345 506251 402379
rect 506285 402345 506298 402379
rect 506238 402179 506298 402345
rect 506238 402145 506251 402179
rect 506285 402145 506298 402179
rect 506238 401979 506298 402145
rect 506238 401945 506251 401979
rect 506285 401945 506298 401979
rect 506238 401779 506298 401945
rect 506238 401745 506251 401779
rect 506285 401745 506298 401779
rect 506238 401622 506298 401745
rect 494958 401371 494971 401405
rect 495005 401371 495018 401405
rect 494958 401005 495018 401371
rect 494958 400971 494971 401005
rect 495005 400971 495018 401005
rect 494958 400605 495018 400971
rect 504358 401093 504418 401276
rect 504358 401059 504371 401093
rect 504405 401059 504418 401093
rect 494958 400571 494971 400605
rect 495005 400571 495018 400605
rect 494958 400205 495018 400571
rect 496838 400653 496898 400934
rect 498718 400906 498778 400934
rect 498508 400893 498778 400906
rect 498508 400859 498591 400893
rect 498625 400859 498778 400893
rect 498508 400846 498778 400859
rect 496838 400619 496851 400653
rect 496885 400619 496898 400653
rect 496838 400320 496898 400619
rect 496998 400367 497058 400836
rect 498318 400825 498378 400836
rect 498094 400824 498378 400825
rect 497344 400790 497371 400824
rect 497425 400790 497443 400824
rect 497493 400790 497515 400824
rect 497561 400790 497587 400824
rect 497629 400790 497659 400824
rect 497697 400790 497731 400824
rect 497765 400790 497799 400824
rect 497837 400790 497867 400824
rect 497909 400790 497935 400824
rect 497981 400790 498003 400824
rect 498053 400790 498071 400824
rect 498125 400791 498378 400824
rect 498125 400790 498152 400791
rect 498318 400573 498378 400791
rect 498544 400653 498604 400756
rect 498544 400619 498557 400653
rect 498591 400619 498604 400653
rect 498318 400539 498353 400573
rect 496998 400366 497362 400367
rect 496998 400333 497371 400366
rect 496998 400320 497058 400333
rect 497344 400332 497371 400333
rect 497425 400332 497443 400366
rect 497493 400332 497515 400366
rect 497561 400332 497587 400366
rect 497629 400332 497659 400366
rect 497697 400332 497731 400366
rect 497765 400332 497799 400366
rect 497837 400332 497867 400366
rect 497909 400332 497935 400366
rect 497981 400332 498003 400366
rect 498053 400332 498071 400366
rect 498125 400332 498152 400366
rect 498318 400320 498378 400539
rect 498544 400389 498604 400619
rect 498544 400355 498557 400389
rect 498591 400355 498604 400389
rect 498544 400320 498604 400355
rect 498718 400653 498778 400846
rect 498718 400619 498731 400653
rect 498765 400619 498778 400653
rect 498718 400320 498778 400619
rect 504358 400893 504418 401059
rect 504358 400859 504371 400893
rect 504405 400859 504418 400893
rect 504358 400693 504418 400859
rect 506238 401093 506298 401276
rect 506238 401059 506251 401093
rect 506285 401059 506298 401093
rect 506238 400893 506298 401059
rect 506238 400859 506251 400893
rect 506285 400859 506298 400893
rect 504358 400659 504371 400693
rect 504405 400659 504418 400693
rect 504358 400493 504418 400659
rect 504358 400459 504371 400493
rect 504405 400459 504418 400493
rect 494958 400171 494971 400205
rect 495005 400171 495018 400205
rect 494958 399805 495018 400171
rect 504358 400293 504418 400459
rect 506238 400693 506298 400859
rect 506238 400659 506251 400693
rect 506285 400659 506298 400693
rect 506238 400493 506298 400659
rect 506238 400459 506251 400493
rect 506285 400459 506298 400493
rect 506238 400364 506298 400459
rect 504358 400259 504371 400293
rect 504405 400259 504418 400293
rect 504358 400093 504418 400259
rect 504358 400059 504371 400093
rect 504405 400059 504418 400093
rect 494958 399771 494971 399805
rect 495005 399771 495018 399805
rect 494958 399405 495018 399771
rect 494958 399371 494971 399405
rect 495005 399371 495018 399405
rect 494958 399005 495018 399371
rect 494958 398971 494971 399005
rect 495005 398971 495018 399005
rect 494958 398605 495018 398971
rect 494958 398571 494971 398605
rect 495005 398571 495018 398605
rect 494958 398205 495018 398571
rect 494958 398171 494971 398205
rect 495005 398171 495018 398205
rect 494958 397805 495018 398171
rect 494958 397771 494971 397805
rect 495005 397771 495018 397805
rect 494958 397405 495018 397771
rect 494958 397371 494971 397405
rect 495005 397371 495018 397405
rect 494958 397005 495018 397371
rect 494958 396971 494971 397005
rect 495005 396971 495018 397005
rect 494958 396605 495018 396971
rect 494958 396571 494971 396605
rect 495005 396571 495018 396605
rect 494958 396205 495018 396571
rect 494958 396171 494971 396205
rect 495005 396171 495018 396205
rect 494958 395805 495018 396171
rect 494958 395771 494971 395805
rect 495005 395771 495018 395805
rect 494958 395405 495018 395771
rect 494958 395371 494971 395405
rect 495005 395371 495018 395405
rect 494958 395005 495018 395371
rect 494958 394971 494971 395005
rect 495005 394971 495018 395005
rect 494958 394605 495018 394971
rect 494958 394571 494971 394605
rect 495005 394571 495018 394605
rect 494958 394420 495018 394571
rect 496838 399994 496898 400022
rect 496838 399981 497108 399994
rect 496838 399947 496991 399981
rect 497025 399947 497108 399981
rect 496838 399934 497108 399947
rect 496838 399741 496898 399934
rect 498478 399895 498489 399924
rect 498523 399895 498538 399924
rect 498478 399877 498538 399895
rect 496838 399707 496851 399741
rect 496885 399707 496898 399741
rect 496838 399341 496898 399707
rect 496838 399307 496851 399341
rect 496885 399307 496898 399341
rect 496838 398946 496898 399307
rect 497018 399419 497058 399864
rect 497099 399843 497119 399877
rect 497153 399843 497187 399877
rect 497225 399843 497255 399877
rect 497297 399843 497323 399877
rect 497369 399843 497391 399877
rect 497441 399843 497459 399877
rect 497513 399843 497527 399877
rect 497585 399843 497595 399877
rect 497657 399843 497663 399877
rect 497729 399843 497731 399877
rect 497765 399843 497767 399877
rect 497833 399843 497839 399877
rect 497901 399843 497911 399877
rect 497969 399843 497983 399877
rect 498037 399843 498055 399877
rect 498105 399843 498127 399877
rect 498173 399843 498199 399877
rect 498241 399843 498271 399877
rect 498309 399843 498343 399877
rect 498377 399843 498538 399877
rect 497018 399385 497119 399419
rect 497153 399385 497187 399419
rect 497225 399385 497255 399419
rect 497297 399385 497323 399419
rect 497369 399385 497391 399419
rect 497441 399385 497459 399419
rect 497513 399385 497527 399419
rect 497585 399385 497595 399419
rect 497657 399385 497663 399419
rect 497729 399385 497731 399419
rect 497765 399385 497767 399419
rect 497833 399385 497839 399419
rect 497901 399385 497911 399419
rect 497969 399385 497983 399419
rect 498037 399385 498055 399419
rect 498105 399385 498127 399419
rect 498173 399385 498199 399419
rect 498241 399385 498271 399419
rect 498309 399385 498343 399419
rect 498377 399385 498397 399419
rect 496838 398941 496978 398946
rect 496838 398907 496851 398941
rect 496885 398907 496978 398941
rect 496838 398881 496978 398907
rect 496838 398847 496941 398881
rect 496975 398847 496978 398881
rect 496838 398786 496978 398847
rect 496838 398541 496898 398786
rect 496838 398507 496851 398541
rect 496885 398507 496898 398541
rect 496838 398141 496898 398507
rect 496838 398107 496851 398141
rect 496885 398107 496898 398141
rect 496838 397741 496898 398107
rect 496838 397707 496851 397741
rect 496885 397707 496898 397741
rect 496838 397646 496898 397707
rect 497018 398503 497058 399385
rect 498478 398961 498538 399843
rect 497099 398927 497119 398961
rect 497153 398927 497187 398961
rect 497225 398927 497255 398961
rect 497297 398927 497323 398961
rect 497369 398927 497391 398961
rect 497441 398927 497459 398961
rect 497513 398927 497527 398961
rect 497585 398927 497595 398961
rect 497657 398927 497663 398961
rect 497729 398927 497731 398961
rect 497765 398927 497767 398961
rect 497833 398927 497839 398961
rect 497901 398927 497911 398961
rect 497969 398927 497983 398961
rect 498037 398927 498055 398961
rect 498105 398927 498127 398961
rect 498173 398927 498199 398961
rect 498241 398927 498271 398961
rect 498309 398927 498343 398961
rect 498377 398927 498538 398961
rect 497018 398469 497119 398503
rect 497153 398469 497187 398503
rect 497225 398469 497255 398503
rect 497297 398469 497323 398503
rect 497369 398469 497391 398503
rect 497441 398469 497459 398503
rect 497513 398469 497527 398503
rect 497585 398469 497595 398503
rect 497657 398469 497663 398503
rect 497729 398469 497731 398503
rect 497765 398469 497767 398503
rect 497833 398469 497839 398503
rect 497901 398469 497911 398503
rect 497969 398469 497983 398503
rect 498037 398469 498055 398503
rect 498105 398469 498127 398503
rect 498173 398469 498199 398503
rect 498241 398469 498271 398503
rect 498309 398469 498343 398503
rect 498377 398469 498397 398503
rect 496838 397581 496978 397646
rect 496838 397547 496941 397581
rect 496975 397547 496978 397581
rect 496838 397486 496978 397547
rect 497018 397587 497058 398469
rect 498478 398045 498538 398927
rect 497099 398011 497119 398045
rect 497153 398011 497187 398045
rect 497225 398011 497255 398045
rect 497297 398011 497323 398045
rect 497369 398011 497391 398045
rect 497441 398011 497459 398045
rect 497513 398011 497527 398045
rect 497585 398011 497595 398045
rect 497657 398011 497663 398045
rect 497729 398011 497731 398045
rect 497765 398011 497767 398045
rect 497833 398011 497839 398045
rect 497901 398011 497911 398045
rect 497969 398011 497983 398045
rect 498037 398011 498055 398045
rect 498105 398011 498127 398045
rect 498173 398011 498199 398045
rect 498241 398011 498271 398045
rect 498309 398011 498343 398045
rect 498377 398011 498538 398045
rect 497018 397553 497119 397587
rect 497153 397553 497187 397587
rect 497225 397553 497255 397587
rect 497297 397553 497323 397587
rect 497369 397553 497391 397587
rect 497441 397553 497459 397587
rect 497513 397553 497527 397587
rect 497585 397553 497595 397587
rect 497657 397553 497663 397587
rect 497729 397553 497731 397587
rect 497765 397553 497767 397587
rect 497833 397553 497839 397587
rect 497901 397553 497911 397587
rect 497969 397553 497983 397587
rect 498037 397553 498055 397587
rect 498105 397553 498127 397587
rect 498173 397553 498199 397587
rect 498241 397553 498271 397587
rect 498309 397553 498343 397587
rect 498377 397553 498397 397587
rect 496838 397341 496898 397486
rect 496838 397307 496851 397341
rect 496885 397307 496898 397341
rect 496838 396941 496898 397307
rect 496838 396907 496851 396941
rect 496885 396907 496898 396941
rect 496838 396541 496898 396907
rect 496838 396507 496851 396541
rect 496885 396507 496898 396541
rect 496838 396346 496898 396507
rect 497018 396671 497058 397553
rect 498478 397129 498538 398011
rect 497099 397095 497119 397129
rect 497153 397095 497187 397129
rect 497225 397095 497255 397129
rect 497297 397095 497323 397129
rect 497369 397095 497391 397129
rect 497441 397095 497459 397129
rect 497513 397095 497527 397129
rect 497585 397095 497595 397129
rect 497657 397095 497663 397129
rect 497729 397095 497731 397129
rect 497765 397095 497767 397129
rect 497833 397095 497839 397129
rect 497901 397095 497911 397129
rect 497969 397095 497983 397129
rect 498037 397095 498055 397129
rect 498105 397095 498127 397129
rect 498173 397095 498199 397129
rect 498241 397095 498271 397129
rect 498309 397095 498343 397129
rect 498377 397095 498538 397129
rect 497018 396637 497119 396671
rect 497153 396637 497187 396671
rect 497225 396637 497255 396671
rect 497297 396637 497323 396671
rect 497369 396637 497391 396671
rect 497441 396637 497459 396671
rect 497513 396637 497527 396671
rect 497585 396637 497595 396671
rect 497657 396637 497663 396671
rect 497729 396637 497731 396671
rect 497765 396637 497767 396671
rect 497833 396637 497839 396671
rect 497901 396637 497911 396671
rect 497969 396637 497983 396671
rect 498037 396637 498055 396671
rect 498105 396637 498127 396671
rect 498173 396637 498199 396671
rect 498241 396637 498271 396671
rect 498309 396637 498343 396671
rect 498377 396637 498397 396671
rect 496838 396281 496978 396346
rect 496838 396247 496941 396281
rect 496975 396247 496978 396281
rect 496838 396186 496978 396247
rect 496838 396141 496898 396186
rect 496838 396107 496851 396141
rect 496885 396107 496898 396141
rect 496838 395741 496898 396107
rect 496838 395707 496851 395741
rect 496885 395707 496898 395741
rect 496838 395341 496898 395707
rect 496838 395307 496851 395341
rect 496885 395307 496898 395341
rect 496838 395046 496898 395307
rect 497018 395755 497058 396637
rect 498478 396213 498538 397095
rect 497099 396179 497119 396213
rect 497153 396179 497187 396213
rect 497225 396179 497255 396213
rect 497297 396179 497323 396213
rect 497369 396179 497391 396213
rect 497441 396179 497459 396213
rect 497513 396179 497527 396213
rect 497585 396179 497595 396213
rect 497657 396179 497663 396213
rect 497729 396179 497731 396213
rect 497765 396179 497767 396213
rect 497833 396179 497839 396213
rect 497901 396179 497911 396213
rect 497969 396179 497983 396213
rect 498037 396179 498055 396213
rect 498105 396179 498127 396213
rect 498173 396179 498199 396213
rect 498241 396179 498271 396213
rect 498309 396179 498343 396213
rect 498377 396179 498538 396213
rect 497018 395721 497119 395755
rect 497153 395721 497187 395755
rect 497225 395721 497255 395755
rect 497297 395721 497323 395755
rect 497369 395721 497391 395755
rect 497441 395721 497459 395755
rect 497513 395721 497527 395755
rect 497585 395721 497595 395755
rect 497657 395721 497663 395755
rect 497729 395721 497731 395755
rect 497765 395721 497767 395755
rect 497833 395721 497839 395755
rect 497901 395721 497911 395755
rect 497969 395721 497983 395755
rect 498037 395721 498055 395755
rect 498105 395721 498127 395755
rect 498173 395721 498199 395755
rect 498241 395721 498271 395755
rect 498309 395721 498343 395755
rect 498377 395721 498397 395755
rect 496838 394981 496978 395046
rect 496838 394947 496941 394981
rect 496975 394947 496978 394981
rect 496838 394941 496978 394947
rect 496838 394907 496851 394941
rect 496885 394907 496978 394941
rect 496838 394886 496978 394907
rect 496838 394541 496898 394886
rect 496838 394507 496851 394541
rect 496885 394507 496898 394541
rect 496838 394141 496898 394507
rect 493078 393939 493138 394122
rect 493078 393905 493091 393939
rect 493125 393905 493138 393939
rect 493078 393739 493138 393905
rect 493078 393705 493091 393739
rect 493125 393705 493138 393739
rect 493078 393539 493138 393705
rect 494958 393939 495018 394122
rect 494958 393905 494971 393939
rect 495005 393905 495018 393939
rect 494958 393739 495018 393905
rect 494958 393705 494971 393739
rect 495005 393705 495018 393739
rect 493078 393505 493091 393539
rect 493125 393505 493138 393539
rect 493078 393339 493138 393505
rect 493078 393305 493091 393339
rect 493125 393305 493138 393339
rect 493078 393139 493138 393305
rect 494958 393539 495018 393705
rect 494958 393505 494971 393539
rect 495005 393505 495018 393539
rect 494958 393339 495018 393505
rect 494958 393305 494971 393339
rect 495005 393305 495018 393339
rect 494958 393210 495018 393305
rect 493078 393105 493091 393139
rect 493125 393105 493138 393139
rect 493078 392939 493138 393105
rect 493078 392905 493091 392939
rect 493125 392905 493138 392939
rect 493078 392739 493138 392905
rect 493078 392705 493091 392739
rect 493125 392705 493138 392739
rect 493078 392539 493138 392705
rect 494018 393139 495018 393210
rect 494018 393123 494971 393139
rect 494018 392681 494057 393123
rect 494159 393105 494971 393123
rect 495005 393105 495018 393139
rect 494159 392939 495018 393105
rect 494159 392905 494971 392939
rect 495005 392905 495018 392939
rect 494159 392739 495018 392905
rect 494159 392705 494971 392739
rect 495005 392705 495018 392739
rect 494159 392681 495018 392705
rect 494018 392594 495018 392681
rect 493078 392505 493091 392539
rect 493125 392505 493138 392539
rect 493078 392339 493138 392505
rect 493078 392305 493091 392339
rect 493125 392305 493138 392339
rect 493078 392139 493138 392305
rect 493078 392105 493091 392139
rect 493125 392105 493138 392139
rect 494958 392539 495018 392594
rect 494958 392505 494971 392539
rect 495005 392505 495018 392539
rect 494958 392339 495018 392505
rect 494958 392305 494971 392339
rect 495005 392305 495018 392339
rect 494958 392139 495018 392305
rect 493078 391939 493138 392105
rect 493078 391905 493091 391939
rect 493125 391905 493138 391939
rect 493078 391682 493138 391905
rect 493913 391682 494303 392114
rect 494958 392105 494971 392139
rect 495005 392105 495018 392139
rect 494958 391939 495018 392105
rect 494958 391905 494971 391939
rect 495005 391905 495018 391939
rect 494958 391682 495018 391905
rect 496838 394107 496851 394141
rect 496885 394107 496898 394141
rect 496838 393746 496898 394107
rect 497018 394839 497058 395721
rect 498478 395297 498538 396179
rect 497099 395263 497119 395297
rect 497153 395263 497187 395297
rect 497225 395263 497255 395297
rect 497297 395263 497323 395297
rect 497369 395263 497391 395297
rect 497441 395263 497459 395297
rect 497513 395263 497527 395297
rect 497585 395263 497595 395297
rect 497657 395263 497663 395297
rect 497729 395263 497731 395297
rect 497765 395263 497767 395297
rect 497833 395263 497839 395297
rect 497901 395263 497911 395297
rect 497969 395263 497983 395297
rect 498037 395263 498055 395297
rect 498105 395263 498127 395297
rect 498173 395263 498199 395297
rect 498241 395263 498271 395297
rect 498309 395263 498343 395297
rect 498377 395263 498538 395297
rect 497018 394805 497119 394839
rect 497153 394805 497187 394839
rect 497225 394805 497255 394839
rect 497297 394805 497323 394839
rect 497369 394805 497391 394839
rect 497441 394805 497459 394839
rect 497513 394805 497527 394839
rect 497585 394805 497595 394839
rect 497657 394805 497663 394839
rect 497729 394805 497731 394839
rect 497765 394805 497767 394839
rect 497833 394805 497839 394839
rect 497901 394805 497911 394839
rect 497969 394805 497983 394839
rect 498037 394805 498055 394839
rect 498105 394805 498127 394839
rect 498173 394805 498199 394839
rect 498241 394805 498271 394839
rect 498309 394805 498343 394839
rect 498377 394805 498397 394839
rect 497018 393923 497058 394805
rect 498478 394381 498538 395263
rect 497099 394347 497119 394381
rect 497153 394347 497187 394381
rect 497225 394347 497255 394381
rect 497297 394347 497323 394381
rect 497369 394347 497391 394381
rect 497441 394347 497459 394381
rect 497513 394347 497527 394381
rect 497585 394347 497595 394381
rect 497657 394347 497663 394381
rect 497729 394347 497731 394381
rect 497765 394347 497767 394381
rect 497833 394347 497839 394381
rect 497901 394347 497911 394381
rect 497969 394347 497983 394381
rect 498037 394347 498055 394381
rect 498105 394347 498127 394381
rect 498173 394347 498199 394381
rect 498241 394347 498271 394381
rect 498309 394347 498343 394381
rect 498377 394347 498538 394381
rect 497018 393889 497119 393923
rect 497153 393889 497187 393923
rect 497225 393889 497255 393923
rect 497297 393889 497323 393923
rect 497369 393889 497391 393923
rect 497441 393889 497459 393923
rect 497513 393889 497527 393923
rect 497585 393889 497595 393923
rect 497657 393889 497663 393923
rect 497729 393889 497731 393923
rect 497765 393889 497767 393923
rect 497833 393889 497839 393923
rect 497901 393889 497911 393923
rect 497969 393889 497983 393923
rect 498037 393889 498055 393923
rect 498105 393889 498127 393923
rect 498173 393889 498199 393923
rect 498241 393889 498271 393923
rect 498309 393889 498343 393923
rect 498377 393889 498397 393923
rect 496838 393741 496978 393746
rect 496838 393707 496851 393741
rect 496885 393707 496978 393741
rect 496838 393681 496978 393707
rect 496838 393647 496941 393681
rect 496975 393647 496978 393681
rect 496838 393586 496978 393647
rect 496838 393341 496898 393586
rect 496838 393307 496851 393341
rect 496885 393307 496898 393341
rect 496838 392941 496898 393307
rect 496838 392907 496851 392941
rect 496885 392907 496898 392941
rect 496838 392541 496898 392907
rect 496838 392507 496851 392541
rect 496885 392507 496898 392541
rect 496838 392446 496898 392507
rect 497018 393007 497058 393889
rect 498478 393465 498538 394347
rect 497099 393431 497119 393465
rect 497153 393431 497187 393465
rect 497225 393431 497255 393465
rect 497297 393431 497323 393465
rect 497369 393431 497391 393465
rect 497441 393431 497459 393465
rect 497513 393431 497527 393465
rect 497585 393431 497595 393465
rect 497657 393431 497663 393465
rect 497729 393431 497731 393465
rect 497765 393431 497767 393465
rect 497833 393431 497839 393465
rect 497901 393431 497911 393465
rect 497969 393431 497983 393465
rect 498037 393431 498055 393465
rect 498105 393431 498127 393465
rect 498173 393431 498199 393465
rect 498241 393431 498271 393465
rect 498309 393431 498343 393465
rect 498377 393431 498538 393465
rect 497018 392973 497119 393007
rect 497153 392973 497187 393007
rect 497225 392973 497255 393007
rect 497297 392973 497323 393007
rect 497369 392973 497391 393007
rect 497441 392973 497459 393007
rect 497513 392973 497527 393007
rect 497585 392973 497595 393007
rect 497657 392973 497663 393007
rect 497729 392973 497731 393007
rect 497765 392973 497767 393007
rect 497833 392973 497839 393007
rect 497901 392973 497911 393007
rect 497969 392973 497983 393007
rect 498037 392973 498055 393007
rect 498105 392973 498127 393007
rect 498173 392973 498199 393007
rect 498241 392973 498271 393007
rect 498309 392973 498343 393007
rect 498377 392973 498397 393007
rect 496838 392381 496978 392446
rect 496838 392347 496941 392381
rect 496975 392347 496978 392381
rect 496838 392286 496978 392347
rect 496838 392141 496898 392286
rect 496838 392107 496851 392141
rect 496885 392107 496898 392141
rect 496838 391741 496898 392107
rect 496838 391707 496851 391741
rect 496885 391707 496898 391741
rect 496838 391341 496898 391707
rect 496838 391307 496851 391341
rect 496885 391307 496898 391341
rect 496838 391146 496898 391307
rect 497018 392091 497058 392973
rect 498478 392549 498538 393431
rect 497099 392515 497119 392549
rect 497153 392515 497187 392549
rect 497225 392515 497255 392549
rect 497297 392515 497323 392549
rect 497369 392515 497391 392549
rect 497441 392515 497459 392549
rect 497513 392515 497527 392549
rect 497585 392515 497595 392549
rect 497657 392515 497663 392549
rect 497729 392515 497731 392549
rect 497765 392515 497767 392549
rect 497833 392515 497839 392549
rect 497901 392515 497911 392549
rect 497969 392515 497983 392549
rect 498037 392515 498055 392549
rect 498105 392515 498127 392549
rect 498173 392515 498199 392549
rect 498241 392515 498271 392549
rect 498309 392515 498343 392549
rect 498377 392515 498538 392549
rect 497018 392057 497119 392091
rect 497153 392057 497187 392091
rect 497225 392057 497255 392091
rect 497297 392057 497323 392091
rect 497369 392057 497391 392091
rect 497441 392057 497459 392091
rect 497513 392057 497527 392091
rect 497585 392057 497595 392091
rect 497657 392057 497663 392091
rect 497729 392057 497731 392091
rect 497765 392057 497767 392091
rect 497833 392057 497839 392091
rect 497901 392057 497911 392091
rect 497969 392057 497983 392091
rect 498037 392057 498055 392091
rect 498105 392057 498127 392091
rect 498173 392057 498199 392091
rect 498241 392057 498271 392091
rect 498309 392057 498343 392091
rect 498377 392057 498397 392091
rect 497018 391175 497058 392057
rect 498478 391633 498538 392515
rect 497099 391599 497119 391633
rect 497153 391599 497187 391633
rect 497225 391599 497255 391633
rect 497297 391599 497323 391633
rect 497369 391599 497391 391633
rect 497441 391599 497459 391633
rect 497513 391599 497527 391633
rect 497585 391599 497595 391633
rect 497657 391599 497663 391633
rect 497729 391599 497731 391633
rect 497765 391599 497767 391633
rect 497833 391599 497839 391633
rect 497901 391599 497911 391633
rect 497969 391599 497983 391633
rect 498037 391599 498055 391633
rect 498105 391599 498127 391633
rect 498173 391599 498199 391633
rect 498241 391599 498271 391633
rect 498309 391599 498343 391633
rect 498377 391599 498538 391633
rect 493078 390853 493138 391134
rect 494958 391106 495018 391134
rect 494748 391093 495018 391106
rect 494748 391059 494831 391093
rect 494865 391059 495018 391093
rect 494748 391046 495018 391059
rect 493078 390819 493091 390853
rect 493125 390819 493138 390853
rect 493078 390520 493138 390819
rect 493238 390567 493298 391036
rect 494558 391025 494618 391036
rect 494334 391024 494618 391025
rect 493584 390990 493611 391024
rect 493665 390990 493683 391024
rect 493733 390990 493755 391024
rect 493801 390990 493827 391024
rect 493869 390990 493899 391024
rect 493937 390990 493971 391024
rect 494005 390990 494039 391024
rect 494077 390990 494107 391024
rect 494149 390990 494175 391024
rect 494221 390990 494243 391024
rect 494293 390990 494311 391024
rect 494365 390991 494618 391024
rect 494365 390990 494392 390991
rect 493238 390566 493602 390567
rect 493238 390533 493611 390566
rect 493238 390520 493298 390533
rect 493584 390532 493611 390533
rect 493665 390532 493683 390566
rect 493733 390532 493755 390566
rect 493801 390532 493827 390566
rect 493869 390532 493899 390566
rect 493937 390532 493971 390566
rect 494005 390532 494039 390566
rect 494077 390532 494107 390566
rect 494149 390532 494175 390566
rect 494221 390532 494243 390566
rect 494293 390532 494311 390566
rect 494365 390532 494392 390566
rect 494558 390520 494618 390991
rect 494784 390913 494844 390956
rect 494784 390879 494817 390913
rect 494784 390853 494844 390879
rect 494784 390819 494797 390853
rect 494831 390819 494844 390853
rect 494784 390520 494844 390819
rect 494958 390853 495018 391046
rect 494958 390819 494971 390853
rect 495005 390819 495018 390853
rect 494958 390520 495018 390819
rect 496838 391081 496978 391146
rect 496838 391047 496941 391081
rect 496975 391047 496978 391081
rect 496838 390986 496978 391047
rect 497018 391141 497119 391175
rect 497153 391141 497187 391175
rect 497225 391141 497255 391175
rect 497297 391141 497323 391175
rect 497369 391141 497391 391175
rect 497441 391141 497459 391175
rect 497513 391141 497527 391175
rect 497585 391141 497595 391175
rect 497657 391141 497663 391175
rect 497729 391141 497731 391175
rect 497765 391141 497767 391175
rect 497833 391141 497839 391175
rect 497901 391141 497911 391175
rect 497969 391141 497983 391175
rect 498037 391141 498055 391175
rect 498105 391141 498127 391175
rect 498173 391141 498199 391175
rect 498241 391141 498271 391175
rect 498309 391141 498343 391175
rect 498377 391141 498397 391175
rect 496838 390941 496898 390986
rect 496838 390907 496851 390941
rect 496885 390907 496898 390941
rect 496838 390541 496898 390907
rect 496838 390507 496851 390541
rect 496885 390507 496898 390541
rect 493078 390194 493138 390222
rect 493078 390181 493348 390194
rect 493078 390147 493231 390181
rect 493265 390147 493348 390181
rect 493078 390134 493348 390147
rect 493078 389941 493138 390134
rect 494718 390077 494778 390124
rect 493078 389907 493091 389941
rect 493125 389907 493138 389941
rect 493078 389541 493138 389907
rect 493078 389507 493091 389541
rect 493125 389507 493138 389541
rect 493078 389146 493138 389507
rect 493258 389619 493298 390064
rect 493339 390043 493359 390077
rect 493393 390043 493427 390077
rect 493465 390043 493495 390077
rect 493537 390043 493563 390077
rect 493609 390043 493631 390077
rect 493681 390043 493699 390077
rect 493753 390043 493767 390077
rect 493825 390043 493835 390077
rect 493897 390043 493903 390077
rect 493969 390043 493971 390077
rect 494005 390043 494007 390077
rect 494073 390043 494079 390077
rect 494141 390043 494151 390077
rect 494209 390043 494223 390077
rect 494277 390043 494295 390077
rect 494345 390043 494367 390077
rect 494413 390043 494439 390077
rect 494481 390043 494511 390077
rect 494549 390043 494583 390077
rect 494617 390043 494778 390077
rect 493258 389585 493359 389619
rect 493393 389585 493427 389619
rect 493465 389585 493495 389619
rect 493537 389585 493563 389619
rect 493609 389585 493631 389619
rect 493681 389585 493699 389619
rect 493753 389585 493767 389619
rect 493825 389585 493835 389619
rect 493897 389585 493903 389619
rect 493969 389585 493971 389619
rect 494005 389585 494007 389619
rect 494073 389585 494079 389619
rect 494141 389585 494151 389619
rect 494209 389585 494223 389619
rect 494277 389585 494295 389619
rect 494345 389585 494367 389619
rect 494413 389585 494439 389619
rect 494481 389585 494511 389619
rect 494549 389585 494583 389619
rect 494617 389585 494637 389619
rect 493078 389141 493218 389146
rect 493078 389107 493091 389141
rect 493125 389107 493218 389141
rect 493078 389081 493218 389107
rect 493078 389047 493181 389081
rect 493215 389047 493218 389081
rect 493078 388986 493218 389047
rect 493078 388741 493138 388986
rect 493078 388707 493091 388741
rect 493125 388707 493138 388741
rect 493078 388341 493138 388707
rect 493078 388307 493091 388341
rect 493125 388307 493138 388341
rect 493078 387941 493138 388307
rect 493078 387907 493091 387941
rect 493125 387907 493138 387941
rect 493078 387846 493138 387907
rect 493258 388703 493298 389585
rect 494718 389161 494778 390043
rect 493339 389127 493359 389161
rect 493393 389127 493427 389161
rect 493465 389127 493495 389161
rect 493537 389127 493563 389161
rect 493609 389127 493631 389161
rect 493681 389127 493699 389161
rect 493753 389127 493767 389161
rect 493825 389127 493835 389161
rect 493897 389127 493903 389161
rect 493969 389127 493971 389161
rect 494005 389127 494007 389161
rect 494073 389127 494079 389161
rect 494141 389127 494151 389161
rect 494209 389127 494223 389161
rect 494277 389127 494295 389161
rect 494345 389127 494367 389161
rect 494413 389127 494439 389161
rect 494481 389127 494511 389161
rect 494549 389127 494583 389161
rect 494617 389127 494778 389161
rect 493258 388669 493359 388703
rect 493393 388669 493427 388703
rect 493465 388669 493495 388703
rect 493537 388669 493563 388703
rect 493609 388669 493631 388703
rect 493681 388669 493699 388703
rect 493753 388669 493767 388703
rect 493825 388669 493835 388703
rect 493897 388669 493903 388703
rect 493969 388669 493971 388703
rect 494005 388669 494007 388703
rect 494073 388669 494079 388703
rect 494141 388669 494151 388703
rect 494209 388669 494223 388703
rect 494277 388669 494295 388703
rect 494345 388669 494367 388703
rect 494413 388669 494439 388703
rect 494481 388669 494511 388703
rect 494549 388669 494583 388703
rect 494617 388669 494637 388703
rect 493078 387781 493218 387846
rect 493078 387747 493181 387781
rect 493215 387747 493218 387781
rect 493078 387686 493218 387747
rect 493258 387787 493298 388669
rect 494718 388245 494778 389127
rect 493339 388211 493359 388245
rect 493393 388211 493427 388245
rect 493465 388211 493495 388245
rect 493537 388211 493563 388245
rect 493609 388211 493631 388245
rect 493681 388211 493699 388245
rect 493753 388211 493767 388245
rect 493825 388211 493835 388245
rect 493897 388211 493903 388245
rect 493969 388211 493971 388245
rect 494005 388211 494007 388245
rect 494073 388211 494079 388245
rect 494141 388211 494151 388245
rect 494209 388211 494223 388245
rect 494277 388211 494295 388245
rect 494345 388211 494367 388245
rect 494413 388211 494439 388245
rect 494481 388211 494511 388245
rect 494549 388211 494583 388245
rect 494617 388211 494778 388245
rect 493258 387753 493359 387787
rect 493393 387753 493427 387787
rect 493465 387753 493495 387787
rect 493537 387753 493563 387787
rect 493609 387753 493631 387787
rect 493681 387753 493699 387787
rect 493753 387753 493767 387787
rect 493825 387753 493835 387787
rect 493897 387753 493903 387787
rect 493969 387753 493971 387787
rect 494005 387753 494007 387787
rect 494073 387753 494079 387787
rect 494141 387753 494151 387787
rect 494209 387753 494223 387787
rect 494277 387753 494295 387787
rect 494345 387753 494367 387787
rect 494413 387753 494439 387787
rect 494481 387753 494511 387787
rect 494549 387753 494583 387787
rect 494617 387753 494637 387787
rect 493078 387541 493138 387686
rect 493078 387507 493091 387541
rect 493125 387507 493138 387541
rect 493078 387141 493138 387507
rect 493078 387107 493091 387141
rect 493125 387107 493138 387141
rect 493078 386741 493138 387107
rect 493078 386707 493091 386741
rect 493125 386707 493138 386741
rect 493078 386546 493138 386707
rect 493258 386871 493298 387753
rect 494718 387329 494778 388211
rect 493339 387295 493359 387329
rect 493393 387295 493427 387329
rect 493465 387295 493495 387329
rect 493537 387295 493563 387329
rect 493609 387295 493631 387329
rect 493681 387295 493699 387329
rect 493753 387295 493767 387329
rect 493825 387295 493835 387329
rect 493897 387295 493903 387329
rect 493969 387295 493971 387329
rect 494005 387295 494007 387329
rect 494073 387295 494079 387329
rect 494141 387295 494151 387329
rect 494209 387295 494223 387329
rect 494277 387295 494295 387329
rect 494345 387295 494367 387329
rect 494413 387295 494439 387329
rect 494481 387295 494511 387329
rect 494549 387295 494583 387329
rect 494617 387295 494778 387329
rect 493258 386837 493359 386871
rect 493393 386837 493427 386871
rect 493465 386837 493495 386871
rect 493537 386837 493563 386871
rect 493609 386837 493631 386871
rect 493681 386837 493699 386871
rect 493753 386837 493767 386871
rect 493825 386837 493835 386871
rect 493897 386837 493903 386871
rect 493969 386837 493971 386871
rect 494005 386837 494007 386871
rect 494073 386837 494079 386871
rect 494141 386837 494151 386871
rect 494209 386837 494223 386871
rect 494277 386837 494295 386871
rect 494345 386837 494367 386871
rect 494413 386837 494439 386871
rect 494481 386837 494511 386871
rect 494549 386837 494583 386871
rect 494617 386837 494637 386871
rect 493078 386481 493218 386546
rect 493078 386447 493181 386481
rect 493215 386447 493218 386481
rect 493078 386386 493218 386447
rect 493078 386341 493138 386386
rect 493078 386307 493091 386341
rect 493125 386307 493138 386341
rect 493078 385941 493138 386307
rect 493078 385907 493091 385941
rect 493125 385907 493138 385941
rect 493078 385541 493138 385907
rect 493078 385507 493091 385541
rect 493125 385507 493138 385541
rect 493078 385246 493138 385507
rect 493258 385955 493298 386837
rect 494718 386413 494778 387295
rect 493339 386379 493359 386413
rect 493393 386379 493427 386413
rect 493465 386379 493495 386413
rect 493537 386379 493563 386413
rect 493609 386379 493631 386413
rect 493681 386379 493699 386413
rect 493753 386379 493767 386413
rect 493825 386379 493835 386413
rect 493897 386379 493903 386413
rect 493969 386379 493971 386413
rect 494005 386379 494007 386413
rect 494073 386379 494079 386413
rect 494141 386379 494151 386413
rect 494209 386379 494223 386413
rect 494277 386379 494295 386413
rect 494345 386379 494367 386413
rect 494413 386379 494439 386413
rect 494481 386379 494511 386413
rect 494549 386379 494583 386413
rect 494617 386379 494778 386413
rect 493258 385921 493359 385955
rect 493393 385921 493427 385955
rect 493465 385921 493495 385955
rect 493537 385921 493563 385955
rect 493609 385921 493631 385955
rect 493681 385921 493699 385955
rect 493753 385921 493767 385955
rect 493825 385921 493835 385955
rect 493897 385921 493903 385955
rect 493969 385921 493971 385955
rect 494005 385921 494007 385955
rect 494073 385921 494079 385955
rect 494141 385921 494151 385955
rect 494209 385921 494223 385955
rect 494277 385921 494295 385955
rect 494345 385921 494367 385955
rect 494413 385921 494439 385955
rect 494481 385921 494511 385955
rect 494549 385921 494583 385955
rect 494617 385921 494637 385955
rect 493078 385181 493218 385246
rect 493078 385147 493181 385181
rect 493215 385147 493218 385181
rect 493078 385141 493218 385147
rect 493078 385107 493091 385141
rect 493125 385107 493218 385141
rect 493078 385086 493218 385107
rect 493078 384741 493138 385086
rect 493078 384707 493091 384741
rect 493125 384707 493138 384741
rect 493078 384341 493138 384707
rect 493078 384307 493091 384341
rect 493125 384307 493138 384341
rect 493078 383946 493138 384307
rect 493258 385039 493298 385921
rect 494718 385497 494778 386379
rect 493339 385463 493359 385497
rect 493393 385463 493427 385497
rect 493465 385463 493495 385497
rect 493537 385463 493563 385497
rect 493609 385463 493631 385497
rect 493681 385463 493699 385497
rect 493753 385463 493767 385497
rect 493825 385463 493835 385497
rect 493897 385463 493903 385497
rect 493969 385463 493971 385497
rect 494005 385463 494007 385497
rect 494073 385463 494079 385497
rect 494141 385463 494151 385497
rect 494209 385463 494223 385497
rect 494277 385463 494295 385497
rect 494345 385463 494367 385497
rect 494413 385463 494439 385497
rect 494481 385463 494511 385497
rect 494549 385463 494583 385497
rect 494617 385463 494778 385497
rect 494824 389941 494884 390124
rect 494824 389907 494837 389941
rect 494871 389907 494884 389941
rect 494824 389541 494884 389907
rect 494824 389507 494837 389541
rect 494871 389507 494884 389541
rect 494824 389141 494884 389507
rect 494824 389107 494837 389141
rect 494871 389107 494884 389141
rect 494824 388741 494884 389107
rect 494824 388707 494837 388741
rect 494871 388707 494884 388741
rect 494824 388341 494884 388707
rect 494824 388307 494837 388341
rect 494871 388307 494884 388341
rect 494824 387941 494884 388307
rect 494824 387907 494837 387941
rect 494871 387907 494884 387941
rect 494824 387541 494884 387907
rect 494824 387507 494837 387541
rect 494871 387507 494884 387541
rect 494824 387141 494884 387507
rect 494824 387107 494837 387141
rect 494871 387107 494884 387141
rect 494824 386741 494884 387107
rect 494824 386707 494837 386741
rect 494871 386707 494884 386741
rect 494824 386341 494884 386707
rect 494824 386307 494837 386341
rect 494871 386307 494884 386341
rect 494824 385941 494884 386307
rect 494824 385907 494837 385941
rect 494871 385907 494884 385941
rect 494824 385541 494884 385907
rect 494824 385507 494837 385541
rect 494871 385507 494884 385541
rect 494824 385485 494884 385507
rect 493258 385005 493359 385039
rect 493393 385005 493427 385039
rect 493465 385005 493495 385039
rect 493537 385005 493563 385039
rect 493609 385005 493631 385039
rect 493681 385005 493699 385039
rect 493753 385005 493767 385039
rect 493825 385005 493835 385039
rect 493897 385005 493903 385039
rect 493969 385005 493971 385039
rect 494005 385005 494007 385039
rect 494073 385005 494079 385039
rect 494141 385005 494151 385039
rect 494209 385005 494223 385039
rect 494277 385005 494295 385039
rect 494345 385005 494367 385039
rect 494413 385005 494439 385039
rect 494481 385005 494511 385039
rect 494549 385005 494583 385039
rect 494617 385005 494637 385039
rect 493258 384123 493298 385005
rect 494718 384581 494778 385463
rect 494851 385451 494884 385485
rect 493339 384547 493359 384581
rect 493393 384547 493427 384581
rect 493465 384547 493495 384581
rect 493537 384547 493563 384581
rect 493609 384547 493631 384581
rect 493681 384547 493699 384581
rect 493753 384547 493767 384581
rect 493825 384547 493835 384581
rect 493897 384547 493903 384581
rect 493969 384547 493971 384581
rect 494005 384547 494007 384581
rect 494073 384547 494079 384581
rect 494141 384547 494151 384581
rect 494209 384547 494223 384581
rect 494277 384547 494295 384581
rect 494345 384547 494367 384581
rect 494413 384547 494439 384581
rect 494481 384547 494511 384581
rect 494549 384547 494583 384581
rect 494617 384547 494778 384581
rect 493258 384089 493359 384123
rect 493393 384089 493427 384123
rect 493465 384089 493495 384123
rect 493537 384089 493563 384123
rect 493609 384089 493631 384123
rect 493681 384089 493699 384123
rect 493753 384089 493767 384123
rect 493825 384089 493835 384123
rect 493897 384089 493903 384123
rect 493969 384089 493971 384123
rect 494005 384089 494007 384123
rect 494073 384089 494079 384123
rect 494141 384089 494151 384123
rect 494209 384089 494223 384123
rect 494277 384089 494295 384123
rect 494345 384089 494367 384123
rect 494413 384089 494439 384123
rect 494481 384089 494511 384123
rect 494549 384089 494583 384123
rect 494617 384089 494637 384123
rect 493078 383941 493218 383946
rect 493078 383907 493091 383941
rect 493125 383907 493218 383941
rect 493078 383881 493218 383907
rect 493078 383847 493181 383881
rect 493215 383847 493218 383881
rect 493078 383786 493218 383847
rect 493078 383541 493138 383786
rect 493078 383507 493091 383541
rect 493125 383507 493138 383541
rect 493078 383141 493138 383507
rect 493078 383107 493091 383141
rect 493125 383107 493138 383141
rect 493078 382741 493138 383107
rect 493078 382707 493091 382741
rect 493125 382707 493138 382741
rect 493078 382646 493138 382707
rect 493258 383207 493298 384089
rect 494718 383665 494778 384547
rect 493339 383631 493359 383665
rect 493393 383631 493427 383665
rect 493465 383631 493495 383665
rect 493537 383631 493563 383665
rect 493609 383631 493631 383665
rect 493681 383631 493699 383665
rect 493753 383631 493767 383665
rect 493825 383631 493835 383665
rect 493897 383631 493903 383665
rect 493969 383631 493971 383665
rect 494005 383631 494007 383665
rect 494073 383631 494079 383665
rect 494141 383631 494151 383665
rect 494209 383631 494223 383665
rect 494277 383631 494295 383665
rect 494345 383631 494367 383665
rect 494413 383631 494439 383665
rect 494481 383631 494511 383665
rect 494549 383631 494583 383665
rect 494617 383631 494778 383665
rect 493258 383173 493359 383207
rect 493393 383173 493427 383207
rect 493465 383173 493495 383207
rect 493537 383173 493563 383207
rect 493609 383173 493631 383207
rect 493681 383173 493699 383207
rect 493753 383173 493767 383207
rect 493825 383173 493835 383207
rect 493897 383173 493903 383207
rect 493969 383173 493971 383207
rect 494005 383173 494007 383207
rect 494073 383173 494079 383207
rect 494141 383173 494151 383207
rect 494209 383173 494223 383207
rect 494277 383173 494295 383207
rect 494345 383173 494367 383207
rect 494413 383173 494439 383207
rect 494481 383173 494511 383207
rect 494549 383173 494583 383207
rect 494617 383173 494637 383207
rect 493078 382581 493218 382646
rect 493078 382547 493181 382581
rect 493215 382547 493218 382581
rect 493078 382486 493218 382547
rect 493078 382341 493138 382486
rect 493078 382307 493091 382341
rect 493125 382307 493138 382341
rect 493078 381941 493138 382307
rect 493078 381907 493091 381941
rect 493125 381907 493138 381941
rect 493078 381541 493138 381907
rect 493078 381507 493091 381541
rect 493125 381507 493138 381541
rect 493078 381346 493138 381507
rect 493258 382291 493298 383173
rect 494718 382749 494778 383631
rect 493339 382715 493359 382749
rect 493393 382715 493427 382749
rect 493465 382715 493495 382749
rect 493537 382715 493563 382749
rect 493609 382715 493631 382749
rect 493681 382715 493699 382749
rect 493753 382715 493767 382749
rect 493825 382715 493835 382749
rect 493897 382715 493903 382749
rect 493969 382715 493971 382749
rect 494005 382715 494007 382749
rect 494073 382715 494079 382749
rect 494141 382715 494151 382749
rect 494209 382715 494223 382749
rect 494277 382715 494295 382749
rect 494345 382715 494367 382749
rect 494413 382715 494439 382749
rect 494481 382715 494511 382749
rect 494549 382715 494583 382749
rect 494617 382715 494778 382749
rect 493258 382257 493359 382291
rect 493393 382257 493427 382291
rect 493465 382257 493495 382291
rect 493537 382257 493563 382291
rect 493609 382257 493631 382291
rect 493681 382257 493699 382291
rect 493753 382257 493767 382291
rect 493825 382257 493835 382291
rect 493897 382257 493903 382291
rect 493969 382257 493971 382291
rect 494005 382257 494007 382291
rect 494073 382257 494079 382291
rect 494141 382257 494151 382291
rect 494209 382257 494223 382291
rect 494277 382257 494295 382291
rect 494345 382257 494367 382291
rect 494413 382257 494439 382291
rect 494481 382257 494511 382291
rect 494549 382257 494583 382291
rect 494617 382257 494637 382291
rect 493258 381375 493298 382257
rect 494718 381833 494778 382715
rect 493339 381799 493359 381833
rect 493393 381799 493427 381833
rect 493465 381799 493495 381833
rect 493537 381799 493563 381833
rect 493609 381799 493631 381833
rect 493681 381799 493699 381833
rect 493753 381799 493767 381833
rect 493825 381799 493835 381833
rect 493897 381799 493903 381833
rect 493969 381799 493971 381833
rect 494005 381799 494007 381833
rect 494073 381799 494079 381833
rect 494141 381799 494151 381833
rect 494209 381799 494223 381833
rect 494277 381799 494295 381833
rect 494345 381799 494367 381833
rect 494413 381799 494439 381833
rect 494481 381799 494511 381833
rect 494549 381799 494583 381833
rect 494617 381799 494778 381833
rect 493078 381281 493218 381346
rect 493078 381247 493181 381281
rect 493215 381247 493218 381281
rect 493078 381186 493218 381247
rect 493258 381341 493359 381375
rect 493393 381341 493427 381375
rect 493465 381341 493495 381375
rect 493537 381341 493563 381375
rect 493609 381341 493631 381375
rect 493681 381341 493699 381375
rect 493753 381341 493767 381375
rect 493825 381341 493835 381375
rect 493897 381341 493903 381375
rect 493969 381341 493971 381375
rect 494005 381341 494007 381375
rect 494073 381341 494079 381375
rect 494141 381341 494151 381375
rect 494209 381341 494223 381375
rect 494277 381341 494295 381375
rect 494345 381341 494367 381375
rect 494413 381341 494439 381375
rect 494481 381341 494511 381375
rect 494549 381341 494583 381375
rect 494617 381341 494637 381375
rect 493078 381141 493138 381186
rect 493078 381107 493091 381141
rect 493125 381107 493138 381141
rect 493078 380741 493138 381107
rect 493078 380707 493091 380741
rect 493125 380707 493138 380741
rect 493078 380341 493138 380707
rect 493078 380307 493091 380341
rect 493125 380307 493138 380341
rect 493078 380046 493138 380307
rect 493258 380459 493298 381341
rect 494718 380917 494778 381799
rect 493339 380883 493359 380917
rect 493393 380883 493427 380917
rect 493465 380883 493495 380917
rect 493537 380883 493563 380917
rect 493609 380883 493631 380917
rect 493681 380883 493699 380917
rect 493753 380883 493767 380917
rect 493825 380883 493835 380917
rect 493897 380883 493903 380917
rect 493969 380883 493971 380917
rect 494005 380883 494007 380917
rect 494073 380883 494079 380917
rect 494141 380883 494151 380917
rect 494209 380883 494223 380917
rect 494277 380883 494295 380917
rect 494345 380883 494367 380917
rect 494413 380883 494439 380917
rect 494481 380883 494511 380917
rect 494549 380883 494583 380917
rect 494617 380883 494778 380917
rect 493258 380425 493359 380459
rect 493393 380425 493427 380459
rect 493465 380425 493495 380459
rect 493537 380425 493563 380459
rect 493609 380425 493631 380459
rect 493681 380425 493699 380459
rect 493753 380425 493767 380459
rect 493825 380425 493835 380459
rect 493897 380425 493903 380459
rect 493969 380425 493971 380459
rect 494005 380425 494007 380459
rect 494073 380425 494079 380459
rect 494141 380425 494151 380459
rect 494209 380425 494223 380459
rect 494277 380425 494295 380459
rect 494345 380425 494367 380459
rect 494413 380425 494439 380459
rect 494481 380425 494511 380459
rect 494549 380425 494583 380459
rect 494617 380425 494637 380459
rect 493078 379981 493218 380046
rect 493078 379947 493181 379981
rect 493215 379947 493218 379981
rect 493078 379941 493218 379947
rect 493078 379907 493091 379941
rect 493125 379907 493218 379941
rect 493078 379886 493218 379907
rect 493078 379541 493138 379886
rect 493078 379507 493091 379541
rect 493125 379507 493138 379541
rect 493078 379141 493138 379507
rect 493078 379107 493091 379141
rect 493125 379107 493138 379141
rect 493078 378746 493138 379107
rect 493258 379543 493298 380425
rect 494718 380001 494778 380883
rect 493339 379967 493359 380001
rect 493393 379967 493427 380001
rect 493465 379967 493495 380001
rect 493537 379967 493563 380001
rect 493609 379967 493631 380001
rect 493681 379967 493699 380001
rect 493753 379967 493767 380001
rect 493825 379967 493835 380001
rect 493897 379967 493903 380001
rect 493969 379967 493971 380001
rect 494005 379967 494007 380001
rect 494073 379967 494079 380001
rect 494141 379967 494151 380001
rect 494209 379967 494223 380001
rect 494277 379967 494295 380001
rect 494345 379967 494367 380001
rect 494413 379967 494439 380001
rect 494481 379967 494511 380001
rect 494549 379967 494583 380001
rect 494617 379967 494778 380001
rect 493258 379509 493359 379543
rect 493393 379509 493427 379543
rect 493465 379509 493495 379543
rect 493537 379509 493563 379543
rect 493609 379509 493631 379543
rect 493681 379509 493699 379543
rect 493753 379509 493767 379543
rect 493825 379509 493835 379543
rect 493897 379509 493903 379543
rect 493969 379509 493971 379543
rect 494005 379509 494007 379543
rect 494073 379509 494079 379543
rect 494141 379509 494151 379543
rect 494209 379509 494223 379543
rect 494277 379509 494295 379543
rect 494345 379509 494367 379543
rect 494413 379509 494439 379543
rect 494481 379509 494511 379543
rect 494549 379509 494583 379543
rect 494617 379509 494637 379543
rect 493078 378741 493218 378746
rect 493078 378707 493091 378741
rect 493125 378707 493218 378741
rect 493078 378681 493218 378707
rect 493078 378647 493181 378681
rect 493215 378647 493218 378681
rect 493078 378586 493218 378647
rect 493258 378627 493298 379509
rect 494718 379085 494778 379967
rect 493339 379051 493359 379085
rect 493393 379051 493427 379085
rect 493465 379051 493495 379085
rect 493537 379051 493563 379085
rect 493609 379051 493631 379085
rect 493681 379051 493699 379085
rect 493753 379051 493767 379085
rect 493825 379051 493835 379085
rect 493897 379051 493903 379085
rect 493969 379051 493971 379085
rect 494005 379051 494007 379085
rect 494073 379051 494079 379085
rect 494141 379051 494151 379085
rect 494209 379051 494223 379085
rect 494277 379051 494295 379085
rect 494345 379051 494367 379085
rect 494413 379051 494439 379085
rect 494481 379051 494511 379085
rect 494549 379051 494583 379085
rect 494617 379051 494778 379085
rect 493258 378593 493359 378627
rect 493393 378593 493427 378627
rect 493465 378593 493495 378627
rect 493537 378593 493563 378627
rect 493609 378593 493631 378627
rect 493681 378593 493699 378627
rect 493753 378593 493767 378627
rect 493825 378593 493835 378627
rect 493897 378593 493903 378627
rect 493969 378593 493971 378627
rect 494005 378593 494007 378627
rect 494073 378593 494079 378627
rect 494141 378593 494151 378627
rect 494209 378593 494223 378627
rect 494277 378593 494295 378627
rect 494345 378593 494367 378627
rect 494413 378593 494439 378627
rect 494481 378593 494511 378627
rect 494549 378593 494583 378627
rect 494617 378593 494637 378627
rect 493078 378341 493138 378586
rect 493078 378307 493091 378341
rect 493125 378307 493138 378341
rect 493078 377941 493138 378307
rect 493078 377907 493091 377941
rect 493125 377907 493138 377941
rect 493078 377541 493138 377907
rect 493078 377507 493091 377541
rect 493125 377507 493138 377541
rect 493078 377446 493138 377507
rect 493258 377711 493298 378593
rect 494718 378169 494778 379051
rect 493339 378135 493359 378169
rect 493393 378135 493427 378169
rect 493465 378135 493495 378169
rect 493537 378135 493563 378169
rect 493609 378135 493631 378169
rect 493681 378135 493699 378169
rect 493753 378135 493767 378169
rect 493825 378135 493835 378169
rect 493897 378135 493903 378169
rect 493969 378135 493971 378169
rect 494005 378135 494007 378169
rect 494073 378135 494079 378169
rect 494141 378135 494151 378169
rect 494209 378135 494223 378169
rect 494277 378135 494295 378169
rect 494345 378135 494367 378169
rect 494413 378135 494439 378169
rect 494481 378135 494511 378169
rect 494549 378135 494583 378169
rect 494617 378135 494778 378169
rect 493258 377677 493359 377711
rect 493393 377677 493427 377711
rect 493465 377677 493495 377711
rect 493537 377677 493563 377711
rect 493609 377677 493631 377711
rect 493681 377677 493699 377711
rect 493753 377677 493767 377711
rect 493825 377677 493835 377711
rect 493897 377677 493903 377711
rect 493969 377677 493971 377711
rect 494005 377677 494007 377711
rect 494073 377677 494079 377711
rect 494141 377677 494151 377711
rect 494209 377677 494223 377711
rect 494277 377677 494295 377711
rect 494345 377677 494367 377711
rect 494413 377677 494439 377711
rect 494481 377677 494511 377711
rect 494549 377677 494583 377711
rect 494617 377677 494637 377711
rect 493078 377381 493218 377446
rect 493078 377347 493181 377381
rect 493215 377347 493218 377381
rect 493078 377286 493218 377347
rect 493078 377141 493138 377286
rect 493078 377107 493091 377141
rect 493125 377107 493138 377141
rect 493078 376741 493138 377107
rect 493078 376707 493091 376741
rect 493125 376707 493138 376741
rect 493078 376341 493138 376707
rect 493078 376307 493091 376341
rect 493125 376307 493138 376341
rect 493078 376146 493138 376307
rect 493258 376795 493298 377677
rect 494718 377253 494778 378135
rect 493339 377219 493359 377253
rect 493393 377219 493427 377253
rect 493465 377219 493495 377253
rect 493537 377219 493563 377253
rect 493609 377219 493631 377253
rect 493681 377219 493699 377253
rect 493753 377219 493767 377253
rect 493825 377219 493835 377253
rect 493897 377219 493903 377253
rect 493969 377219 493971 377253
rect 494005 377219 494007 377253
rect 494073 377219 494079 377253
rect 494141 377219 494151 377253
rect 494209 377219 494223 377253
rect 494277 377219 494295 377253
rect 494345 377219 494367 377253
rect 494413 377219 494439 377253
rect 494481 377219 494511 377253
rect 494549 377219 494583 377253
rect 494617 377219 494778 377253
rect 493258 376761 493359 376795
rect 493393 376761 493427 376795
rect 493465 376761 493495 376795
rect 493537 376761 493563 376795
rect 493609 376761 493631 376795
rect 493681 376761 493699 376795
rect 493753 376761 493767 376795
rect 493825 376761 493835 376795
rect 493897 376761 493903 376795
rect 493969 376761 493971 376795
rect 494005 376761 494007 376795
rect 494073 376761 494079 376795
rect 494141 376761 494151 376795
rect 494209 376761 494223 376795
rect 494277 376761 494295 376795
rect 494345 376761 494367 376795
rect 494413 376761 494439 376795
rect 494481 376761 494511 376795
rect 494549 376761 494583 376795
rect 494617 376761 494637 376795
rect 493078 376081 493218 376146
rect 493078 376047 493181 376081
rect 493215 376047 493218 376081
rect 493078 375986 493218 376047
rect 493078 375941 493138 375986
rect 493078 375907 493091 375941
rect 493125 375907 493138 375941
rect 493078 375541 493138 375907
rect 493078 375507 493091 375541
rect 493125 375507 493138 375541
rect 493078 375141 493138 375507
rect 493078 375107 493091 375141
rect 493125 375107 493138 375141
rect 493078 374846 493138 375107
rect 493258 375879 493298 376761
rect 494718 376337 494778 377219
rect 493339 376303 493359 376337
rect 493393 376303 493427 376337
rect 493465 376303 493495 376337
rect 493537 376303 493563 376337
rect 493609 376303 493631 376337
rect 493681 376303 493699 376337
rect 493753 376303 493767 376337
rect 493825 376303 493835 376337
rect 493897 376303 493903 376337
rect 493969 376303 493971 376337
rect 494005 376303 494007 376337
rect 494073 376303 494079 376337
rect 494141 376303 494151 376337
rect 494209 376303 494223 376337
rect 494277 376303 494295 376337
rect 494345 376303 494367 376337
rect 494413 376303 494439 376337
rect 494481 376303 494511 376337
rect 494549 376303 494583 376337
rect 494617 376303 494778 376337
rect 493258 375845 493359 375879
rect 493393 375845 493427 375879
rect 493465 375845 493495 375879
rect 493537 375845 493563 375879
rect 493609 375845 493631 375879
rect 493681 375845 493699 375879
rect 493753 375845 493767 375879
rect 493825 375845 493835 375879
rect 493897 375845 493903 375879
rect 493969 375845 493971 375879
rect 494005 375845 494007 375879
rect 494073 375845 494079 375879
rect 494141 375845 494151 375879
rect 494209 375845 494223 375879
rect 494277 375845 494295 375879
rect 494345 375845 494367 375879
rect 494413 375845 494439 375879
rect 494481 375845 494511 375879
rect 494549 375845 494583 375879
rect 494617 375845 494637 375879
rect 493258 374963 493298 375845
rect 494718 375421 494778 376303
rect 493339 375387 493359 375421
rect 493393 375387 493427 375421
rect 493465 375387 493495 375421
rect 493537 375387 493563 375421
rect 493609 375387 493631 375421
rect 493681 375387 493699 375421
rect 493753 375387 493767 375421
rect 493825 375387 493835 375421
rect 493897 375387 493903 375421
rect 493969 375387 493971 375421
rect 494005 375387 494007 375421
rect 494073 375387 494079 375421
rect 494141 375387 494151 375421
rect 494209 375387 494223 375421
rect 494277 375387 494295 375421
rect 494345 375387 494367 375421
rect 494413 375387 494439 375421
rect 494481 375387 494511 375421
rect 494549 375387 494583 375421
rect 494617 375387 494778 375421
rect 493258 374929 493359 374963
rect 493393 374929 493427 374963
rect 493465 374929 493495 374963
rect 493537 374929 493563 374963
rect 493609 374929 493631 374963
rect 493681 374929 493699 374963
rect 493753 374929 493767 374963
rect 493825 374929 493835 374963
rect 493897 374929 493903 374963
rect 493969 374929 493971 374963
rect 494005 374929 494007 374963
rect 494073 374929 494079 374963
rect 494141 374929 494151 374963
rect 494209 374929 494223 374963
rect 494277 374929 494295 374963
rect 494345 374929 494367 374963
rect 494413 374929 494439 374963
rect 494481 374929 494511 374963
rect 494549 374929 494583 374963
rect 494617 374929 494637 374963
rect 493078 374781 493218 374846
rect 493078 374747 493181 374781
rect 493215 374747 493218 374781
rect 493078 374741 493218 374747
rect 493078 374707 493091 374741
rect 493125 374707 493218 374741
rect 493078 374686 493218 374707
rect 493078 374341 493138 374686
rect 493078 374307 493091 374341
rect 493125 374307 493138 374341
rect 493078 373941 493138 374307
rect 493078 373907 493091 373941
rect 493125 373907 493138 373941
rect 493078 373546 493138 373907
rect 493258 374047 493298 374929
rect 494718 374505 494778 375387
rect 493339 374471 493359 374505
rect 493393 374471 493427 374505
rect 493465 374471 493495 374505
rect 493537 374471 493563 374505
rect 493609 374471 493631 374505
rect 493681 374471 493699 374505
rect 493753 374471 493767 374505
rect 493825 374471 493835 374505
rect 493897 374471 493903 374505
rect 493969 374471 493971 374505
rect 494005 374471 494007 374505
rect 494073 374471 494079 374505
rect 494141 374471 494151 374505
rect 494209 374471 494223 374505
rect 494277 374471 494295 374505
rect 494345 374471 494367 374505
rect 494413 374471 494439 374505
rect 494481 374471 494511 374505
rect 494549 374471 494583 374505
rect 494617 374471 494778 374505
rect 493258 374013 493359 374047
rect 493393 374013 493427 374047
rect 493465 374013 493495 374047
rect 493537 374013 493563 374047
rect 493609 374013 493631 374047
rect 493681 374013 493699 374047
rect 493753 374013 493767 374047
rect 493825 374013 493835 374047
rect 493897 374013 493903 374047
rect 493969 374013 493971 374047
rect 494005 374013 494007 374047
rect 494073 374013 494079 374047
rect 494141 374013 494151 374047
rect 494209 374013 494223 374047
rect 494277 374013 494295 374047
rect 494345 374013 494367 374047
rect 494413 374013 494439 374047
rect 494481 374013 494511 374047
rect 494549 374013 494583 374047
rect 494617 374013 494637 374047
rect 493078 373541 493218 373546
rect 493078 373507 493091 373541
rect 493125 373507 493218 373541
rect 493078 373481 493218 373507
rect 493078 373447 493181 373481
rect 493215 373447 493218 373481
rect 493078 373386 493218 373447
rect 493078 373141 493138 373386
rect 493078 373107 493091 373141
rect 493125 373107 493138 373141
rect 493078 372741 493138 373107
rect 493078 372707 493091 372741
rect 493125 372707 493138 372741
rect 493078 372341 493138 372707
rect 493078 372307 493091 372341
rect 493125 372307 493138 372341
rect 493078 372246 493138 372307
rect 493258 373131 493298 374013
rect 494718 373589 494778 374471
rect 493339 373555 493359 373589
rect 493393 373555 493427 373589
rect 493465 373555 493495 373589
rect 493537 373555 493563 373589
rect 493609 373555 493631 373589
rect 493681 373555 493699 373589
rect 493753 373555 493767 373589
rect 493825 373555 493835 373589
rect 493897 373555 493903 373589
rect 493969 373555 493971 373589
rect 494005 373555 494007 373589
rect 494073 373555 494079 373589
rect 494141 373555 494151 373589
rect 494209 373555 494223 373589
rect 494277 373555 494295 373589
rect 494345 373555 494367 373589
rect 494413 373555 494439 373589
rect 494481 373555 494511 373589
rect 494549 373555 494583 373589
rect 494617 373555 494778 373589
rect 493258 373097 493359 373131
rect 493393 373097 493427 373131
rect 493465 373097 493495 373131
rect 493537 373097 493563 373131
rect 493609 373097 493631 373131
rect 493681 373097 493699 373131
rect 493753 373097 493767 373131
rect 493825 373097 493835 373131
rect 493897 373097 493903 373131
rect 493969 373097 493971 373131
rect 494005 373097 494007 373131
rect 494073 373097 494079 373131
rect 494141 373097 494151 373131
rect 494209 373097 494223 373131
rect 494277 373097 494295 373131
rect 494345 373097 494367 373131
rect 494413 373097 494439 373131
rect 494481 373097 494511 373131
rect 494549 373097 494583 373131
rect 494617 373097 494637 373131
rect 493078 372181 493218 372246
rect 493078 372147 493181 372181
rect 493215 372147 493218 372181
rect 493078 372086 493218 372147
rect 493258 372215 493298 373097
rect 494718 372673 494778 373555
rect 493339 372639 493359 372673
rect 493393 372639 493427 372673
rect 493465 372639 493495 372673
rect 493537 372639 493563 372673
rect 493609 372639 493631 372673
rect 493681 372639 493699 372673
rect 493753 372639 493767 372673
rect 493825 372639 493835 372673
rect 493897 372639 493903 372673
rect 493969 372639 493971 372673
rect 494005 372639 494007 372673
rect 494073 372639 494079 372673
rect 494141 372639 494151 372673
rect 494209 372639 494223 372673
rect 494277 372639 494295 372673
rect 494345 372639 494367 372673
rect 494413 372639 494439 372673
rect 494481 372639 494511 372673
rect 494549 372639 494583 372673
rect 494617 372639 494778 372673
rect 493258 372181 493359 372215
rect 493393 372181 493427 372215
rect 493465 372181 493495 372215
rect 493537 372181 493563 372215
rect 493609 372181 493631 372215
rect 493681 372181 493699 372215
rect 493753 372181 493767 372215
rect 493825 372181 493835 372215
rect 493897 372181 493903 372215
rect 493969 372181 493971 372215
rect 494005 372181 494007 372215
rect 494073 372181 494079 372215
rect 494141 372181 494151 372215
rect 494209 372181 494223 372215
rect 494277 372181 494295 372215
rect 494345 372181 494367 372215
rect 494413 372181 494439 372215
rect 494481 372181 494511 372215
rect 494549 372181 494583 372215
rect 494617 372181 494637 372215
rect 493078 371941 493138 372086
rect 493078 371907 493091 371941
rect 493125 371907 493138 371941
rect 493078 371541 493138 371907
rect 493078 371507 493091 371541
rect 493125 371507 493138 371541
rect 493078 371141 493138 371507
rect 493078 371107 493091 371141
rect 493125 371107 493138 371141
rect 493078 370946 493138 371107
rect 493258 371299 493298 372181
rect 494718 371757 494778 372639
rect 493339 371723 493359 371757
rect 493393 371723 493427 371757
rect 493465 371723 493495 371757
rect 493537 371723 493563 371757
rect 493609 371723 493631 371757
rect 493681 371723 493699 371757
rect 493753 371723 493767 371757
rect 493825 371723 493835 371757
rect 493897 371723 493903 371757
rect 493969 371723 493971 371757
rect 494005 371723 494007 371757
rect 494073 371723 494079 371757
rect 494141 371723 494151 371757
rect 494209 371723 494223 371757
rect 494277 371723 494295 371757
rect 494345 371723 494367 371757
rect 494413 371723 494439 371757
rect 494481 371723 494511 371757
rect 494549 371723 494583 371757
rect 494617 371723 494778 371757
rect 493258 371265 493359 371299
rect 493393 371265 493427 371299
rect 493465 371265 493495 371299
rect 493537 371265 493563 371299
rect 493609 371265 493631 371299
rect 493681 371265 493699 371299
rect 493753 371265 493767 371299
rect 493825 371265 493835 371299
rect 493897 371265 493903 371299
rect 493969 371265 493971 371299
rect 494005 371265 494007 371299
rect 494073 371265 494079 371299
rect 494141 371265 494151 371299
rect 494209 371265 494223 371299
rect 494277 371265 494295 371299
rect 494345 371265 494367 371299
rect 494413 371265 494439 371299
rect 494481 371265 494511 371299
rect 494549 371265 494583 371299
rect 494617 371265 494637 371299
rect 493078 370881 493218 370946
rect 493078 370847 493181 370881
rect 493215 370847 493218 370881
rect 493078 370786 493218 370847
rect 493078 370741 493138 370786
rect 493078 370707 493091 370741
rect 493125 370707 493138 370741
rect 493078 370341 493138 370707
rect 493078 370307 493091 370341
rect 493125 370307 493138 370341
rect 493078 369941 493138 370307
rect 493078 369907 493091 369941
rect 493125 369907 493138 369941
rect 493078 369646 493138 369907
rect 493258 370383 493298 371265
rect 494718 370841 494778 371723
rect 493339 370807 493359 370841
rect 493393 370807 493427 370841
rect 493465 370807 493495 370841
rect 493537 370807 493563 370841
rect 493609 370807 493631 370841
rect 493681 370807 493699 370841
rect 493753 370807 493767 370841
rect 493825 370807 493835 370841
rect 493897 370807 493903 370841
rect 493969 370807 493971 370841
rect 494005 370807 494007 370841
rect 494073 370807 494079 370841
rect 494141 370807 494151 370841
rect 494209 370807 494223 370841
rect 494277 370807 494295 370841
rect 494345 370807 494367 370841
rect 494413 370807 494439 370841
rect 494481 370807 494511 370841
rect 494549 370807 494583 370841
rect 494617 370807 494778 370841
rect 493258 370349 493359 370383
rect 493393 370349 493427 370383
rect 493465 370349 493495 370383
rect 493537 370349 493563 370383
rect 493609 370349 493631 370383
rect 493681 370349 493699 370383
rect 493753 370349 493767 370383
rect 493825 370349 493835 370383
rect 493897 370349 493903 370383
rect 493969 370349 493971 370383
rect 494005 370349 494007 370383
rect 494073 370349 494079 370383
rect 494141 370349 494151 370383
rect 494209 370349 494223 370383
rect 494277 370349 494295 370383
rect 494345 370349 494367 370383
rect 494413 370349 494439 370383
rect 494481 370349 494511 370383
rect 494549 370349 494583 370383
rect 494617 370349 494637 370383
rect 493078 369581 493218 369646
rect 493078 369547 493181 369581
rect 493215 369547 493218 369581
rect 493078 369541 493218 369547
rect 493078 369507 493091 369541
rect 493125 369507 493218 369541
rect 493078 369486 493218 369507
rect 493078 369141 493138 369486
rect 493078 369107 493091 369141
rect 493125 369107 493138 369141
rect 493078 368741 493138 369107
rect 493078 368707 493091 368741
rect 493125 368707 493138 368741
rect 493078 368346 493138 368707
rect 493258 369467 493298 370349
rect 494718 369925 494778 370807
rect 493339 369891 493359 369925
rect 493393 369891 493427 369925
rect 493465 369891 493495 369925
rect 493537 369891 493563 369925
rect 493609 369891 493631 369925
rect 493681 369891 493699 369925
rect 493753 369891 493767 369925
rect 493825 369891 493835 369925
rect 493897 369891 493903 369925
rect 493969 369891 493971 369925
rect 494005 369891 494007 369925
rect 494073 369891 494079 369925
rect 494141 369891 494151 369925
rect 494209 369891 494223 369925
rect 494277 369891 494295 369925
rect 494345 369891 494367 369925
rect 494413 369891 494439 369925
rect 494481 369891 494511 369925
rect 494549 369891 494583 369925
rect 494617 369891 494778 369925
rect 493258 369433 493359 369467
rect 493393 369433 493427 369467
rect 493465 369433 493495 369467
rect 493537 369433 493563 369467
rect 493609 369433 493631 369467
rect 493681 369433 493699 369467
rect 493753 369433 493767 369467
rect 493825 369433 493835 369467
rect 493897 369433 493903 369467
rect 493969 369433 493971 369467
rect 494005 369433 494007 369467
rect 494073 369433 494079 369467
rect 494141 369433 494151 369467
rect 494209 369433 494223 369467
rect 494277 369433 494295 369467
rect 494345 369433 494367 369467
rect 494413 369433 494439 369467
rect 494481 369433 494511 369467
rect 494549 369433 494583 369467
rect 494617 369433 494637 369467
rect 493258 368551 493298 369433
rect 494718 369009 494778 369891
rect 493339 368975 493359 369009
rect 493393 368975 493427 369009
rect 493465 368975 493495 369009
rect 493537 368975 493563 369009
rect 493609 368975 493631 369009
rect 493681 368975 493699 369009
rect 493753 368975 493767 369009
rect 493825 368975 493835 369009
rect 493897 368975 493903 369009
rect 493969 368975 493971 369009
rect 494005 368975 494007 369009
rect 494073 368975 494079 369009
rect 494141 368975 494151 369009
rect 494209 368975 494223 369009
rect 494277 368975 494295 369009
rect 494345 368975 494367 369009
rect 494413 368975 494439 369009
rect 494481 368975 494511 369009
rect 494549 368975 494583 369009
rect 494617 368975 494778 369009
rect 493258 368517 493359 368551
rect 493393 368517 493427 368551
rect 493465 368517 493495 368551
rect 493537 368517 493563 368551
rect 493609 368517 493631 368551
rect 493681 368517 493699 368551
rect 493753 368517 493767 368551
rect 493825 368517 493835 368551
rect 493897 368517 493903 368551
rect 493969 368517 493971 368551
rect 494005 368517 494007 368551
rect 494073 368517 494079 368551
rect 494141 368517 494151 368551
rect 494209 368517 494223 368551
rect 494277 368517 494295 368551
rect 494345 368517 494367 368551
rect 494413 368517 494439 368551
rect 494481 368517 494511 368551
rect 494549 368517 494583 368551
rect 494617 368517 494637 368551
rect 493078 368341 493218 368346
rect 493078 368307 493091 368341
rect 493125 368307 493218 368341
rect 493078 368281 493218 368307
rect 493078 368247 493181 368281
rect 493215 368247 493218 368281
rect 493078 368186 493218 368247
rect 493078 367941 493138 368186
rect 493078 367907 493091 367941
rect 493125 367907 493138 367941
rect 493078 367541 493138 367907
rect 493078 367507 493091 367541
rect 493125 367507 493138 367541
rect 493078 367141 493138 367507
rect 493078 367107 493091 367141
rect 493125 367107 493138 367141
rect 493078 367046 493138 367107
rect 493258 367635 493298 368517
rect 494718 368093 494778 368975
rect 493339 368059 493359 368093
rect 493393 368059 493427 368093
rect 493465 368059 493495 368093
rect 493537 368059 493563 368093
rect 493609 368059 493631 368093
rect 493681 368059 493699 368093
rect 493753 368059 493767 368093
rect 493825 368059 493835 368093
rect 493897 368059 493903 368093
rect 493969 368059 493971 368093
rect 494005 368059 494007 368093
rect 494073 368059 494079 368093
rect 494141 368059 494151 368093
rect 494209 368059 494223 368093
rect 494277 368059 494295 368093
rect 494345 368059 494367 368093
rect 494413 368059 494439 368093
rect 494481 368059 494511 368093
rect 494549 368059 494583 368093
rect 494617 368059 494778 368093
rect 493258 367601 493359 367635
rect 493393 367601 493427 367635
rect 493465 367601 493495 367635
rect 493537 367601 493563 367635
rect 493609 367601 493631 367635
rect 493681 367601 493699 367635
rect 493753 367601 493767 367635
rect 493825 367601 493835 367635
rect 493897 367601 493903 367635
rect 493969 367601 493971 367635
rect 494005 367601 494007 367635
rect 494073 367601 494079 367635
rect 494141 367601 494151 367635
rect 494209 367601 494223 367635
rect 494277 367601 494295 367635
rect 494345 367601 494367 367635
rect 494413 367601 494439 367635
rect 494481 367601 494511 367635
rect 494549 367601 494583 367635
rect 494617 367601 494637 367635
rect 493078 366981 493218 367046
rect 493078 366947 493181 366981
rect 493215 366947 493218 366981
rect 493078 366886 493218 366947
rect 493078 366741 493138 366886
rect 493078 366707 493091 366741
rect 493125 366707 493138 366741
rect 493078 366341 493138 366707
rect 493078 366307 493091 366341
rect 493125 366307 493138 366341
rect 493078 365941 493138 366307
rect 493078 365907 493091 365941
rect 493125 365907 493138 365941
rect 493078 365746 493138 365907
rect 493258 366719 493298 367601
rect 494718 367177 494778 368059
rect 493339 367143 493359 367177
rect 493393 367143 493427 367177
rect 493465 367143 493495 367177
rect 493537 367143 493563 367177
rect 493609 367143 493631 367177
rect 493681 367143 493699 367177
rect 493753 367143 493767 367177
rect 493825 367143 493835 367177
rect 493897 367143 493903 367177
rect 493969 367143 493971 367177
rect 494005 367143 494007 367177
rect 494073 367143 494079 367177
rect 494141 367143 494151 367177
rect 494209 367143 494223 367177
rect 494277 367143 494295 367177
rect 494345 367143 494367 367177
rect 494413 367143 494439 367177
rect 494481 367143 494511 367177
rect 494549 367143 494583 367177
rect 494617 367143 494778 367177
rect 493258 366685 493359 366719
rect 493393 366685 493427 366719
rect 493465 366685 493495 366719
rect 493537 366685 493563 366719
rect 493609 366685 493631 366719
rect 493681 366685 493699 366719
rect 493753 366685 493767 366719
rect 493825 366685 493835 366719
rect 493897 366685 493903 366719
rect 493969 366685 493971 366719
rect 494005 366685 494007 366719
rect 494073 366685 494079 366719
rect 494141 366685 494151 366719
rect 494209 366685 494223 366719
rect 494277 366685 494295 366719
rect 494345 366685 494367 366719
rect 494413 366685 494439 366719
rect 494481 366685 494511 366719
rect 494549 366685 494583 366719
rect 494617 366685 494637 366719
rect 493258 365803 493298 366685
rect 494718 366261 494778 367143
rect 493339 366227 493359 366261
rect 493393 366227 493427 366261
rect 493465 366227 493495 366261
rect 493537 366227 493563 366261
rect 493609 366227 493631 366261
rect 493681 366227 493699 366261
rect 493753 366227 493767 366261
rect 493825 366227 493835 366261
rect 493897 366227 493903 366261
rect 493969 366227 493971 366261
rect 494005 366227 494007 366261
rect 494073 366227 494079 366261
rect 494141 366227 494151 366261
rect 494209 366227 494223 366261
rect 494277 366227 494295 366261
rect 494345 366227 494367 366261
rect 494413 366227 494439 366261
rect 494481 366227 494511 366261
rect 494549 366227 494583 366261
rect 494617 366227 494778 366261
rect 493258 365769 493359 365803
rect 493393 365769 493427 365803
rect 493465 365769 493495 365803
rect 493537 365769 493563 365803
rect 493609 365769 493631 365803
rect 493681 365769 493699 365803
rect 493753 365769 493767 365803
rect 493825 365769 493835 365803
rect 493897 365769 493903 365803
rect 493969 365769 493971 365803
rect 494005 365769 494007 365803
rect 494073 365769 494079 365803
rect 494141 365769 494151 365803
rect 494209 365769 494223 365803
rect 494277 365769 494295 365803
rect 494345 365769 494367 365803
rect 494413 365769 494439 365803
rect 494481 365769 494511 365803
rect 494549 365769 494583 365803
rect 494617 365769 494637 365803
rect 493078 365681 493218 365746
rect 493078 365647 493181 365681
rect 493215 365647 493218 365681
rect 493078 365586 493218 365647
rect 493078 365541 493138 365586
rect 493078 365507 493091 365541
rect 493125 365507 493138 365541
rect 493078 365141 493138 365507
rect 493078 365107 493091 365141
rect 493125 365107 493138 365141
rect 493078 364741 493138 365107
rect 493078 364707 493091 364741
rect 493125 364707 493138 364741
rect 493078 364446 493138 364707
rect 493258 364887 493298 365769
rect 494718 365345 494778 366227
rect 493339 365311 493359 365345
rect 493393 365311 493427 365345
rect 493465 365311 493495 365345
rect 493537 365311 493563 365345
rect 493609 365311 493631 365345
rect 493681 365311 493699 365345
rect 493753 365311 493767 365345
rect 493825 365311 493835 365345
rect 493897 365311 493903 365345
rect 493969 365311 493971 365345
rect 494005 365311 494007 365345
rect 494073 365311 494079 365345
rect 494141 365311 494151 365345
rect 494209 365311 494223 365345
rect 494277 365311 494295 365345
rect 494345 365311 494367 365345
rect 494413 365311 494439 365345
rect 494481 365311 494511 365345
rect 494549 365311 494583 365345
rect 494617 365311 494778 365345
rect 493258 364853 493359 364887
rect 493393 364853 493427 364887
rect 493465 364853 493495 364887
rect 493537 364853 493563 364887
rect 493609 364853 493631 364887
rect 493681 364853 493699 364887
rect 493753 364853 493767 364887
rect 493825 364853 493835 364887
rect 493897 364853 493903 364887
rect 493969 364853 493971 364887
rect 494005 364853 494007 364887
rect 494073 364853 494079 364887
rect 494141 364853 494151 364887
rect 494209 364853 494223 364887
rect 494277 364853 494295 364887
rect 494345 364853 494367 364887
rect 494413 364853 494439 364887
rect 494481 364853 494511 364887
rect 494549 364853 494583 364887
rect 494617 364853 494637 364887
rect 493078 364381 493218 364446
rect 493078 364347 493181 364381
rect 493215 364347 493218 364381
rect 493078 364341 493218 364347
rect 493078 364307 493091 364341
rect 493125 364307 493218 364341
rect 493078 364286 493218 364307
rect 493078 363941 493138 364286
rect 493078 363907 493091 363941
rect 493125 363907 493138 363941
rect 493078 363541 493138 363907
rect 493078 363507 493091 363541
rect 493125 363507 493138 363541
rect 493078 363141 493138 363507
rect 493078 363107 493091 363141
rect 493125 363107 493138 363141
rect 493078 362741 493138 363107
rect 493078 362707 493091 362741
rect 493125 362707 493138 362741
rect 493078 362516 493138 362707
rect 493258 363971 493298 364853
rect 494718 364429 494778 365311
rect 493339 364395 493359 364429
rect 493393 364395 493427 364429
rect 493465 364395 493495 364429
rect 493537 364395 493563 364429
rect 493609 364395 493631 364429
rect 493681 364395 493699 364429
rect 493753 364395 493767 364429
rect 493825 364395 493835 364429
rect 493897 364395 493903 364429
rect 493969 364395 493971 364429
rect 494005 364395 494007 364429
rect 494073 364395 494079 364429
rect 494141 364395 494151 364429
rect 494209 364395 494223 364429
rect 494277 364395 494295 364429
rect 494345 364395 494367 364429
rect 494413 364395 494439 364429
rect 494481 364395 494511 364429
rect 494549 364395 494583 364429
rect 494617 364395 494778 364429
rect 493258 363937 493359 363971
rect 493393 363937 493427 363971
rect 493465 363937 493495 363971
rect 493537 363937 493563 363971
rect 493609 363937 493631 363971
rect 493681 363937 493699 363971
rect 493753 363937 493767 363971
rect 493825 363937 493835 363971
rect 493897 363937 493903 363971
rect 493969 363937 493971 363971
rect 494005 363937 494007 363971
rect 494073 363937 494079 363971
rect 494141 363937 494151 363971
rect 494209 363937 494223 363971
rect 494277 363937 494295 363971
rect 494345 363937 494367 363971
rect 494413 363937 494439 363971
rect 494481 363937 494511 363971
rect 494549 363937 494583 363971
rect 494617 363937 494637 363971
rect 493258 363055 493298 363937
rect 494718 363513 494778 364395
rect 493339 363479 493359 363513
rect 493393 363479 493427 363513
rect 493465 363479 493495 363513
rect 493537 363479 493563 363513
rect 493609 363479 493631 363513
rect 493681 363479 493699 363513
rect 493753 363479 493767 363513
rect 493825 363479 493835 363513
rect 493897 363479 493903 363513
rect 493969 363479 493971 363513
rect 494005 363479 494007 363513
rect 494073 363479 494079 363513
rect 494141 363479 494151 363513
rect 494209 363479 494223 363513
rect 494277 363479 494295 363513
rect 494345 363479 494367 363513
rect 494413 363479 494439 363513
rect 494481 363479 494511 363513
rect 494549 363479 494583 363513
rect 494617 363479 494778 363513
rect 493258 363021 493359 363055
rect 493393 363021 493427 363055
rect 493465 363021 493495 363055
rect 493537 363021 493563 363055
rect 493609 363021 493631 363055
rect 493681 363021 493699 363055
rect 493753 363021 493767 363055
rect 493825 363021 493835 363055
rect 493897 363021 493903 363055
rect 493969 363021 493971 363055
rect 494005 363021 494007 363055
rect 494073 363021 494079 363055
rect 494141 363021 494151 363055
rect 494209 363021 494223 363055
rect 494277 363021 494295 363055
rect 494345 363021 494367 363055
rect 494413 363021 494439 363055
rect 494481 363021 494511 363055
rect 494549 363021 494583 363055
rect 494617 363021 494637 363055
rect 493258 362516 493298 363021
rect 494718 362597 494778 363479
rect 493339 362563 493359 362597
rect 493393 362563 493427 362597
rect 493465 362563 493495 362597
rect 493537 362563 493563 362597
rect 493609 362563 493631 362597
rect 493681 362563 493699 362597
rect 493753 362563 493767 362597
rect 493825 362563 493835 362597
rect 493897 362563 493903 362597
rect 493969 362563 493971 362597
rect 494005 362563 494007 362597
rect 494073 362563 494079 362597
rect 494141 362563 494151 362597
rect 494209 362563 494223 362597
rect 494277 362563 494295 362597
rect 494345 362563 494367 362597
rect 494413 362563 494439 362597
rect 494481 362563 494511 362597
rect 494549 362563 494583 362597
rect 494617 362563 494778 362597
rect 494718 362516 494778 362563
rect 494824 385141 494884 385451
rect 494824 385107 494837 385141
rect 494871 385107 494884 385141
rect 494824 384741 494884 385107
rect 494824 384707 494837 384741
rect 494871 384707 494884 384741
rect 494824 384341 494884 384707
rect 494824 384307 494837 384341
rect 494871 384307 494884 384341
rect 494824 383941 494884 384307
rect 494824 383907 494837 383941
rect 494871 383907 494884 383941
rect 494824 383541 494884 383907
rect 494824 383507 494837 383541
rect 494871 383507 494884 383541
rect 494824 383141 494884 383507
rect 494824 383107 494837 383141
rect 494871 383107 494884 383141
rect 494824 382741 494884 383107
rect 494824 382707 494837 382741
rect 494871 382707 494884 382741
rect 494824 382341 494884 382707
rect 494824 382307 494837 382341
rect 494871 382307 494884 382341
rect 494824 381941 494884 382307
rect 494824 381907 494837 381941
rect 494871 381907 494884 381941
rect 494824 381541 494884 381907
rect 494824 381507 494837 381541
rect 494871 381507 494884 381541
rect 494824 381141 494884 381507
rect 494824 381107 494837 381141
rect 494871 381107 494884 381141
rect 494824 380741 494884 381107
rect 494824 380707 494837 380741
rect 494871 380707 494884 380741
rect 494824 380341 494884 380707
rect 494824 380307 494837 380341
rect 494871 380307 494884 380341
rect 494824 379941 494884 380307
rect 494824 379907 494837 379941
rect 494871 379907 494884 379941
rect 494824 379541 494884 379907
rect 494824 379507 494837 379541
rect 494871 379507 494884 379541
rect 494824 379141 494884 379507
rect 494824 379107 494837 379141
rect 494871 379107 494884 379141
rect 494824 378741 494884 379107
rect 494824 378707 494837 378741
rect 494871 378707 494884 378741
rect 494824 378341 494884 378707
rect 494824 378307 494837 378341
rect 494871 378307 494884 378341
rect 494824 377941 494884 378307
rect 494824 377907 494837 377941
rect 494871 377907 494884 377941
rect 494824 377541 494884 377907
rect 494824 377507 494837 377541
rect 494871 377507 494884 377541
rect 494824 377141 494884 377507
rect 494824 377107 494837 377141
rect 494871 377107 494884 377141
rect 494824 376741 494884 377107
rect 494824 376707 494837 376741
rect 494871 376707 494884 376741
rect 494824 376341 494884 376707
rect 494824 376307 494837 376341
rect 494871 376307 494884 376341
rect 494824 375941 494884 376307
rect 494824 375907 494837 375941
rect 494871 375907 494884 375941
rect 494824 375541 494884 375907
rect 494824 375507 494837 375541
rect 494871 375507 494884 375541
rect 494824 375141 494884 375507
rect 494824 375107 494837 375141
rect 494871 375107 494884 375141
rect 494824 374741 494884 375107
rect 494824 374707 494837 374741
rect 494871 374707 494884 374741
rect 494824 374341 494884 374707
rect 494824 374307 494837 374341
rect 494871 374307 494884 374341
rect 494824 373941 494884 374307
rect 494824 373907 494837 373941
rect 494871 373907 494884 373941
rect 494824 373541 494884 373907
rect 494824 373507 494837 373541
rect 494871 373507 494884 373541
rect 494824 373141 494884 373507
rect 494824 373107 494837 373141
rect 494871 373107 494884 373141
rect 494824 372741 494884 373107
rect 494824 372707 494837 372741
rect 494871 372707 494884 372741
rect 494824 372341 494884 372707
rect 494824 372307 494837 372341
rect 494871 372307 494884 372341
rect 494824 371941 494884 372307
rect 494824 371907 494837 371941
rect 494871 371907 494884 371941
rect 494824 371541 494884 371907
rect 494824 371507 494837 371541
rect 494871 371507 494884 371541
rect 494824 371141 494884 371507
rect 494824 371107 494837 371141
rect 494871 371107 494884 371141
rect 494824 370741 494884 371107
rect 494824 370707 494837 370741
rect 494871 370707 494884 370741
rect 494824 370341 494884 370707
rect 494824 370307 494837 370341
rect 494871 370307 494884 370341
rect 494824 369941 494884 370307
rect 494824 369907 494837 369941
rect 494871 369907 494884 369941
rect 494824 369541 494884 369907
rect 494824 369507 494837 369541
rect 494871 369507 494884 369541
rect 494824 369141 494884 369507
rect 494824 369107 494837 369141
rect 494871 369107 494884 369141
rect 494824 368741 494884 369107
rect 494824 368707 494837 368741
rect 494871 368707 494884 368741
rect 494824 368341 494884 368707
rect 494824 368307 494837 368341
rect 494871 368307 494884 368341
rect 494824 367941 494884 368307
rect 494824 367907 494837 367941
rect 494871 367907 494884 367941
rect 494824 367541 494884 367907
rect 494824 367507 494837 367541
rect 494871 367507 494884 367541
rect 494824 367141 494884 367507
rect 494824 367107 494837 367141
rect 494871 367107 494884 367141
rect 494824 366741 494884 367107
rect 494824 366707 494837 366741
rect 494871 366707 494884 366741
rect 494824 366341 494884 366707
rect 494824 366307 494837 366341
rect 494871 366307 494884 366341
rect 494824 365941 494884 366307
rect 494824 365907 494837 365941
rect 494871 365907 494884 365941
rect 494824 365541 494884 365907
rect 494824 365507 494837 365541
rect 494871 365507 494884 365541
rect 494824 365141 494884 365507
rect 494824 365107 494837 365141
rect 494871 365107 494884 365141
rect 494824 364741 494884 365107
rect 494824 364707 494837 364741
rect 494871 364707 494884 364741
rect 494824 364341 494884 364707
rect 494824 364307 494837 364341
rect 494871 364307 494884 364341
rect 494824 363941 494884 364307
rect 494824 363907 494837 363941
rect 494871 363907 494884 363941
rect 494824 363541 494884 363907
rect 494824 363507 494837 363541
rect 494871 363507 494884 363541
rect 494824 363141 494884 363507
rect 494824 363107 494837 363141
rect 494871 363107 494884 363141
rect 494824 362741 494884 363107
rect 494824 362707 494837 362741
rect 494871 362707 494884 362741
rect 494824 362516 494884 362707
rect 494958 389941 495018 390222
rect 494958 389907 494971 389941
rect 495005 389907 495018 389941
rect 494958 389541 495018 389907
rect 494958 389507 494971 389541
rect 495005 389507 495018 389541
rect 494958 389141 495018 389507
rect 494958 389107 494971 389141
rect 495005 389107 495018 389141
rect 494958 388741 495018 389107
rect 494958 388707 494971 388741
rect 495005 388707 495018 388741
rect 494958 388341 495018 388707
rect 494958 388307 494971 388341
rect 495005 388307 495018 388341
rect 494958 387941 495018 388307
rect 494958 387907 494971 387941
rect 495005 387907 495018 387941
rect 494958 387541 495018 387907
rect 494958 387507 494971 387541
rect 495005 387507 495018 387541
rect 494958 387141 495018 387507
rect 494958 387107 494971 387141
rect 495005 387107 495018 387141
rect 494958 386741 495018 387107
rect 494958 386707 494971 386741
rect 495005 386707 495018 386741
rect 494958 386341 495018 386707
rect 494958 386307 494971 386341
rect 495005 386307 495018 386341
rect 494958 385941 495018 386307
rect 494958 385907 494971 385941
rect 495005 385907 495018 385941
rect 494958 385541 495018 385907
rect 494958 385507 494971 385541
rect 495005 385507 495018 385541
rect 494958 385141 495018 385507
rect 494958 385107 494971 385141
rect 495005 385107 495018 385141
rect 494958 384741 495018 385107
rect 494958 384707 494971 384741
rect 495005 384707 495018 384741
rect 494958 384341 495018 384707
rect 494958 384307 494971 384341
rect 495005 384307 495018 384341
rect 494958 383941 495018 384307
rect 494958 383907 494971 383941
rect 495005 383907 495018 383941
rect 494958 383541 495018 383907
rect 494958 383507 494971 383541
rect 495005 383507 495018 383541
rect 494958 383141 495018 383507
rect 494958 383107 494971 383141
rect 495005 383107 495018 383141
rect 494958 382741 495018 383107
rect 494958 382707 494971 382741
rect 495005 382707 495018 382741
rect 494958 382341 495018 382707
rect 494958 382307 494971 382341
rect 495005 382307 495018 382341
rect 494958 381941 495018 382307
rect 494958 381907 494971 381941
rect 495005 381907 495018 381941
rect 494958 381541 495018 381907
rect 494958 381507 494971 381541
rect 495005 381507 495018 381541
rect 494958 381141 495018 381507
rect 494958 381107 494971 381141
rect 495005 381107 495018 381141
rect 494958 380741 495018 381107
rect 494958 380707 494971 380741
rect 495005 380707 495018 380741
rect 494958 380341 495018 380707
rect 494958 380307 494971 380341
rect 495005 380307 495018 380341
rect 494958 379941 495018 380307
rect 494958 379907 494971 379941
rect 495005 379907 495018 379941
rect 494958 379541 495018 379907
rect 494958 379507 494971 379541
rect 495005 379507 495018 379541
rect 494958 379141 495018 379507
rect 494958 379107 494971 379141
rect 495005 379107 495018 379141
rect 494958 378741 495018 379107
rect 494958 378707 494971 378741
rect 495005 378707 495018 378741
rect 494958 378341 495018 378707
rect 494958 378307 494971 378341
rect 495005 378307 495018 378341
rect 494958 377941 495018 378307
rect 494958 377907 494971 377941
rect 495005 377907 495018 377941
rect 494958 377541 495018 377907
rect 494958 377507 494971 377541
rect 495005 377507 495018 377541
rect 494958 377141 495018 377507
rect 494958 377107 494971 377141
rect 495005 377107 495018 377141
rect 494958 376741 495018 377107
rect 494958 376707 494971 376741
rect 495005 376707 495018 376741
rect 494958 376341 495018 376707
rect 494958 376307 494971 376341
rect 495005 376307 495018 376341
rect 494958 375941 495018 376307
rect 494958 375907 494971 375941
rect 495005 375907 495018 375941
rect 494958 375541 495018 375907
rect 494958 375507 494971 375541
rect 495005 375507 495018 375541
rect 494958 375141 495018 375507
rect 494958 375107 494971 375141
rect 495005 375107 495018 375141
rect 494958 374741 495018 375107
rect 494958 374707 494971 374741
rect 495005 374707 495018 374741
rect 494958 374341 495018 374707
rect 494958 374307 494971 374341
rect 495005 374307 495018 374341
rect 494958 373941 495018 374307
rect 494958 373907 494971 373941
rect 495005 373907 495018 373941
rect 494958 373541 495018 373907
rect 494958 373507 494971 373541
rect 495005 373507 495018 373541
rect 494958 373141 495018 373507
rect 494958 373107 494971 373141
rect 495005 373107 495018 373141
rect 494958 372741 495018 373107
rect 494958 372707 494971 372741
rect 495005 372707 495018 372741
rect 494958 372341 495018 372707
rect 494958 372307 494971 372341
rect 495005 372307 495018 372341
rect 496838 390141 496898 390507
rect 496838 390107 496851 390141
rect 496885 390107 496898 390141
rect 496838 389846 496898 390107
rect 497018 390259 497058 391141
rect 498478 390717 498538 391599
rect 497099 390683 497119 390717
rect 497153 390683 497187 390717
rect 497225 390683 497255 390717
rect 497297 390683 497323 390717
rect 497369 390683 497391 390717
rect 497441 390683 497459 390717
rect 497513 390683 497527 390717
rect 497585 390683 497595 390717
rect 497657 390683 497663 390717
rect 497729 390683 497731 390717
rect 497765 390683 497767 390717
rect 497833 390683 497839 390717
rect 497901 390683 497911 390717
rect 497969 390683 497983 390717
rect 498037 390683 498055 390717
rect 498105 390683 498127 390717
rect 498173 390683 498199 390717
rect 498241 390683 498271 390717
rect 498309 390683 498343 390717
rect 498377 390683 498538 390717
rect 497018 390225 497119 390259
rect 497153 390225 497187 390259
rect 497225 390225 497255 390259
rect 497297 390225 497323 390259
rect 497369 390225 497391 390259
rect 497441 390225 497459 390259
rect 497513 390225 497527 390259
rect 497585 390225 497595 390259
rect 497657 390225 497663 390259
rect 497729 390225 497731 390259
rect 497765 390225 497767 390259
rect 497833 390225 497839 390259
rect 497901 390225 497911 390259
rect 497969 390225 497983 390259
rect 498037 390225 498055 390259
rect 498105 390225 498127 390259
rect 498173 390225 498199 390259
rect 498241 390225 498271 390259
rect 498309 390225 498343 390259
rect 498377 390225 498397 390259
rect 496838 389781 496978 389846
rect 496838 389747 496941 389781
rect 496975 389747 496978 389781
rect 496838 389741 496978 389747
rect 496838 389707 496851 389741
rect 496885 389707 496978 389741
rect 496838 389686 496978 389707
rect 496838 389341 496898 389686
rect 496838 389307 496851 389341
rect 496885 389307 496898 389341
rect 496838 388941 496898 389307
rect 496838 388907 496851 388941
rect 496885 388907 496898 388941
rect 496838 388546 496898 388907
rect 497018 389343 497058 390225
rect 498478 389801 498538 390683
rect 497099 389767 497119 389801
rect 497153 389767 497187 389801
rect 497225 389767 497255 389801
rect 497297 389767 497323 389801
rect 497369 389767 497391 389801
rect 497441 389767 497459 389801
rect 497513 389767 497527 389801
rect 497585 389767 497595 389801
rect 497657 389767 497663 389801
rect 497729 389767 497731 389801
rect 497765 389767 497767 389801
rect 497833 389767 497839 389801
rect 497901 389767 497911 389801
rect 497969 389767 497983 389801
rect 498037 389767 498055 389801
rect 498105 389767 498127 389801
rect 498173 389767 498199 389801
rect 498241 389767 498271 389801
rect 498309 389767 498343 389801
rect 498377 389767 498538 389801
rect 497018 389309 497119 389343
rect 497153 389309 497187 389343
rect 497225 389309 497255 389343
rect 497297 389309 497323 389343
rect 497369 389309 497391 389343
rect 497441 389309 497459 389343
rect 497513 389309 497527 389343
rect 497585 389309 497595 389343
rect 497657 389309 497663 389343
rect 497729 389309 497731 389343
rect 497765 389309 497767 389343
rect 497833 389309 497839 389343
rect 497901 389309 497911 389343
rect 497969 389309 497983 389343
rect 498037 389309 498055 389343
rect 498105 389309 498127 389343
rect 498173 389309 498199 389343
rect 498241 389309 498271 389343
rect 498309 389309 498343 389343
rect 498377 389309 498397 389343
rect 496838 388541 496978 388546
rect 496838 388507 496851 388541
rect 496885 388507 496978 388541
rect 496838 388481 496978 388507
rect 496838 388447 496941 388481
rect 496975 388447 496978 388481
rect 496838 388386 496978 388447
rect 497018 388427 497058 389309
rect 498478 388885 498538 389767
rect 497099 388851 497119 388885
rect 497153 388851 497187 388885
rect 497225 388851 497255 388885
rect 497297 388851 497323 388885
rect 497369 388851 497391 388885
rect 497441 388851 497459 388885
rect 497513 388851 497527 388885
rect 497585 388851 497595 388885
rect 497657 388851 497663 388885
rect 497729 388851 497731 388885
rect 497765 388851 497767 388885
rect 497833 388851 497839 388885
rect 497901 388851 497911 388885
rect 497969 388851 497983 388885
rect 498037 388851 498055 388885
rect 498105 388851 498127 388885
rect 498173 388851 498199 388885
rect 498241 388851 498271 388885
rect 498309 388851 498343 388885
rect 498377 388851 498538 388885
rect 497018 388393 497119 388427
rect 497153 388393 497187 388427
rect 497225 388393 497255 388427
rect 497297 388393 497323 388427
rect 497369 388393 497391 388427
rect 497441 388393 497459 388427
rect 497513 388393 497527 388427
rect 497585 388393 497595 388427
rect 497657 388393 497663 388427
rect 497729 388393 497731 388427
rect 497765 388393 497767 388427
rect 497833 388393 497839 388427
rect 497901 388393 497911 388427
rect 497969 388393 497983 388427
rect 498037 388393 498055 388427
rect 498105 388393 498127 388427
rect 498173 388393 498199 388427
rect 498241 388393 498271 388427
rect 498309 388393 498343 388427
rect 498377 388393 498397 388427
rect 496838 388141 496898 388386
rect 496838 388107 496851 388141
rect 496885 388107 496898 388141
rect 496838 387741 496898 388107
rect 496838 387707 496851 387741
rect 496885 387707 496898 387741
rect 496838 387341 496898 387707
rect 496838 387307 496851 387341
rect 496885 387307 496898 387341
rect 496838 387246 496898 387307
rect 497018 387511 497058 388393
rect 498478 387969 498538 388851
rect 497099 387935 497119 387969
rect 497153 387935 497187 387969
rect 497225 387935 497255 387969
rect 497297 387935 497323 387969
rect 497369 387935 497391 387969
rect 497441 387935 497459 387969
rect 497513 387935 497527 387969
rect 497585 387935 497595 387969
rect 497657 387935 497663 387969
rect 497729 387935 497731 387969
rect 497765 387935 497767 387969
rect 497833 387935 497839 387969
rect 497901 387935 497911 387969
rect 497969 387935 497983 387969
rect 498037 387935 498055 387969
rect 498105 387935 498127 387969
rect 498173 387935 498199 387969
rect 498241 387935 498271 387969
rect 498309 387935 498343 387969
rect 498377 387935 498538 387969
rect 497018 387477 497119 387511
rect 497153 387477 497187 387511
rect 497225 387477 497255 387511
rect 497297 387477 497323 387511
rect 497369 387477 497391 387511
rect 497441 387477 497459 387511
rect 497513 387477 497527 387511
rect 497585 387477 497595 387511
rect 497657 387477 497663 387511
rect 497729 387477 497731 387511
rect 497765 387477 497767 387511
rect 497833 387477 497839 387511
rect 497901 387477 497911 387511
rect 497969 387477 497983 387511
rect 498037 387477 498055 387511
rect 498105 387477 498127 387511
rect 498173 387477 498199 387511
rect 498241 387477 498271 387511
rect 498309 387477 498343 387511
rect 498377 387477 498397 387511
rect 496838 387181 496978 387246
rect 496838 387147 496941 387181
rect 496975 387147 496978 387181
rect 496838 387086 496978 387147
rect 496838 386941 496898 387086
rect 496838 386907 496851 386941
rect 496885 386907 496898 386941
rect 496838 386541 496898 386907
rect 496838 386507 496851 386541
rect 496885 386507 496898 386541
rect 496838 386141 496898 386507
rect 496838 386107 496851 386141
rect 496885 386107 496898 386141
rect 496838 385946 496898 386107
rect 497018 386595 497058 387477
rect 498478 387053 498538 387935
rect 497099 387019 497119 387053
rect 497153 387019 497187 387053
rect 497225 387019 497255 387053
rect 497297 387019 497323 387053
rect 497369 387019 497391 387053
rect 497441 387019 497459 387053
rect 497513 387019 497527 387053
rect 497585 387019 497595 387053
rect 497657 387019 497663 387053
rect 497729 387019 497731 387053
rect 497765 387019 497767 387053
rect 497833 387019 497839 387053
rect 497901 387019 497911 387053
rect 497969 387019 497983 387053
rect 498037 387019 498055 387053
rect 498105 387019 498127 387053
rect 498173 387019 498199 387053
rect 498241 387019 498271 387053
rect 498309 387019 498343 387053
rect 498377 387019 498538 387053
rect 497018 386561 497119 386595
rect 497153 386561 497187 386595
rect 497225 386561 497255 386595
rect 497297 386561 497323 386595
rect 497369 386561 497391 386595
rect 497441 386561 497459 386595
rect 497513 386561 497527 386595
rect 497585 386561 497595 386595
rect 497657 386561 497663 386595
rect 497729 386561 497731 386595
rect 497765 386561 497767 386595
rect 497833 386561 497839 386595
rect 497901 386561 497911 386595
rect 497969 386561 497983 386595
rect 498037 386561 498055 386595
rect 498105 386561 498127 386595
rect 498173 386561 498199 386595
rect 498241 386561 498271 386595
rect 498309 386561 498343 386595
rect 498377 386561 498397 386595
rect 496838 385881 496978 385946
rect 496838 385847 496941 385881
rect 496975 385847 496978 385881
rect 496838 385786 496978 385847
rect 496838 385741 496898 385786
rect 496838 385707 496851 385741
rect 496885 385707 496898 385741
rect 496838 385341 496898 385707
rect 496838 385307 496851 385341
rect 496885 385307 496898 385341
rect 496838 384941 496898 385307
rect 496838 384907 496851 384941
rect 496885 384907 496898 384941
rect 496838 384646 496898 384907
rect 497018 385679 497058 386561
rect 498478 386137 498538 387019
rect 497099 386103 497119 386137
rect 497153 386103 497187 386137
rect 497225 386103 497255 386137
rect 497297 386103 497323 386137
rect 497369 386103 497391 386137
rect 497441 386103 497459 386137
rect 497513 386103 497527 386137
rect 497585 386103 497595 386137
rect 497657 386103 497663 386137
rect 497729 386103 497731 386137
rect 497765 386103 497767 386137
rect 497833 386103 497839 386137
rect 497901 386103 497911 386137
rect 497969 386103 497983 386137
rect 498037 386103 498055 386137
rect 498105 386103 498127 386137
rect 498173 386103 498199 386137
rect 498241 386103 498271 386137
rect 498309 386103 498343 386137
rect 498377 386103 498538 386137
rect 497018 385645 497119 385679
rect 497153 385645 497187 385679
rect 497225 385645 497255 385679
rect 497297 385645 497323 385679
rect 497369 385645 497391 385679
rect 497441 385645 497459 385679
rect 497513 385645 497527 385679
rect 497585 385645 497595 385679
rect 497657 385645 497663 385679
rect 497729 385645 497731 385679
rect 497765 385645 497767 385679
rect 497833 385645 497839 385679
rect 497901 385645 497911 385679
rect 497969 385645 497983 385679
rect 498037 385645 498055 385679
rect 498105 385645 498127 385679
rect 498173 385645 498199 385679
rect 498241 385645 498271 385679
rect 498309 385645 498343 385679
rect 498377 385645 498397 385679
rect 497018 384763 497058 385645
rect 498478 385221 498538 386103
rect 497099 385187 497119 385221
rect 497153 385187 497187 385221
rect 497225 385187 497255 385221
rect 497297 385187 497323 385221
rect 497369 385187 497391 385221
rect 497441 385187 497459 385221
rect 497513 385187 497527 385221
rect 497585 385187 497595 385221
rect 497657 385187 497663 385221
rect 497729 385187 497731 385221
rect 497765 385187 497767 385221
rect 497833 385187 497839 385221
rect 497901 385187 497911 385221
rect 497969 385187 497983 385221
rect 498037 385187 498055 385221
rect 498105 385187 498127 385221
rect 498173 385187 498199 385221
rect 498241 385187 498271 385221
rect 498309 385187 498343 385221
rect 498377 385187 498538 385221
rect 497018 384729 497119 384763
rect 497153 384729 497187 384763
rect 497225 384729 497255 384763
rect 497297 384729 497323 384763
rect 497369 384729 497391 384763
rect 497441 384729 497459 384763
rect 497513 384729 497527 384763
rect 497585 384729 497595 384763
rect 497657 384729 497663 384763
rect 497729 384729 497731 384763
rect 497765 384729 497767 384763
rect 497833 384729 497839 384763
rect 497901 384729 497911 384763
rect 497969 384729 497983 384763
rect 498037 384729 498055 384763
rect 498105 384729 498127 384763
rect 498173 384729 498199 384763
rect 498241 384729 498271 384763
rect 498309 384729 498343 384763
rect 498377 384729 498397 384763
rect 496838 384581 496978 384646
rect 496838 384547 496941 384581
rect 496975 384547 496978 384581
rect 496838 384541 496978 384547
rect 496838 384507 496851 384541
rect 496885 384507 496978 384541
rect 496838 384486 496978 384507
rect 496838 384141 496898 384486
rect 496838 384107 496851 384141
rect 496885 384107 496898 384141
rect 496838 383741 496898 384107
rect 496838 383707 496851 383741
rect 496885 383707 496898 383741
rect 496838 383346 496898 383707
rect 497018 383847 497058 384729
rect 498478 384305 498538 385187
rect 497099 384271 497119 384305
rect 497153 384271 497187 384305
rect 497225 384271 497255 384305
rect 497297 384271 497323 384305
rect 497369 384271 497391 384305
rect 497441 384271 497459 384305
rect 497513 384271 497527 384305
rect 497585 384271 497595 384305
rect 497657 384271 497663 384305
rect 497729 384271 497731 384305
rect 497765 384271 497767 384305
rect 497833 384271 497839 384305
rect 497901 384271 497911 384305
rect 497969 384271 497983 384305
rect 498037 384271 498055 384305
rect 498105 384271 498127 384305
rect 498173 384271 498199 384305
rect 498241 384271 498271 384305
rect 498309 384271 498343 384305
rect 498377 384271 498538 384305
rect 497018 383813 497119 383847
rect 497153 383813 497187 383847
rect 497225 383813 497255 383847
rect 497297 383813 497323 383847
rect 497369 383813 497391 383847
rect 497441 383813 497459 383847
rect 497513 383813 497527 383847
rect 497585 383813 497595 383847
rect 497657 383813 497663 383847
rect 497729 383813 497731 383847
rect 497765 383813 497767 383847
rect 497833 383813 497839 383847
rect 497901 383813 497911 383847
rect 497969 383813 497983 383847
rect 498037 383813 498055 383847
rect 498105 383813 498127 383847
rect 498173 383813 498199 383847
rect 498241 383813 498271 383847
rect 498309 383813 498343 383847
rect 498377 383813 498397 383847
rect 496838 383341 496978 383346
rect 496838 383307 496851 383341
rect 496885 383307 496978 383341
rect 496838 383281 496978 383307
rect 496838 383247 496941 383281
rect 496975 383247 496978 383281
rect 496838 383186 496978 383247
rect 496838 382941 496898 383186
rect 496838 382907 496851 382941
rect 496885 382907 496898 382941
rect 496838 382541 496898 382907
rect 496838 382507 496851 382541
rect 496885 382507 496898 382541
rect 496838 382141 496898 382507
rect 496838 382107 496851 382141
rect 496885 382107 496898 382141
rect 496838 382046 496898 382107
rect 497018 382931 497058 383813
rect 498478 383389 498538 384271
rect 497099 383355 497119 383389
rect 497153 383355 497187 383389
rect 497225 383355 497255 383389
rect 497297 383355 497323 383389
rect 497369 383355 497391 383389
rect 497441 383355 497459 383389
rect 497513 383355 497527 383389
rect 497585 383355 497595 383389
rect 497657 383355 497663 383389
rect 497729 383355 497731 383389
rect 497765 383355 497767 383389
rect 497833 383355 497839 383389
rect 497901 383355 497911 383389
rect 497969 383355 497983 383389
rect 498037 383355 498055 383389
rect 498105 383355 498127 383389
rect 498173 383355 498199 383389
rect 498241 383355 498271 383389
rect 498309 383355 498343 383389
rect 498377 383355 498538 383389
rect 497018 382897 497119 382931
rect 497153 382897 497187 382931
rect 497225 382897 497255 382931
rect 497297 382897 497323 382931
rect 497369 382897 497391 382931
rect 497441 382897 497459 382931
rect 497513 382897 497527 382931
rect 497585 382897 497595 382931
rect 497657 382897 497663 382931
rect 497729 382897 497731 382931
rect 497765 382897 497767 382931
rect 497833 382897 497839 382931
rect 497901 382897 497911 382931
rect 497969 382897 497983 382931
rect 498037 382897 498055 382931
rect 498105 382897 498127 382931
rect 498173 382897 498199 382931
rect 498241 382897 498271 382931
rect 498309 382897 498343 382931
rect 498377 382897 498397 382931
rect 496838 381981 496978 382046
rect 496838 381947 496941 381981
rect 496975 381947 496978 381981
rect 496838 381886 496978 381947
rect 497018 382015 497058 382897
rect 498478 382473 498538 383355
rect 497099 382439 497119 382473
rect 497153 382439 497187 382473
rect 497225 382439 497255 382473
rect 497297 382439 497323 382473
rect 497369 382439 497391 382473
rect 497441 382439 497459 382473
rect 497513 382439 497527 382473
rect 497585 382439 497595 382473
rect 497657 382439 497663 382473
rect 497729 382439 497731 382473
rect 497765 382439 497767 382473
rect 497833 382439 497839 382473
rect 497901 382439 497911 382473
rect 497969 382439 497983 382473
rect 498037 382439 498055 382473
rect 498105 382439 498127 382473
rect 498173 382439 498199 382473
rect 498241 382439 498271 382473
rect 498309 382439 498343 382473
rect 498377 382439 498538 382473
rect 497018 381981 497119 382015
rect 497153 381981 497187 382015
rect 497225 381981 497255 382015
rect 497297 381981 497323 382015
rect 497369 381981 497391 382015
rect 497441 381981 497459 382015
rect 497513 381981 497527 382015
rect 497585 381981 497595 382015
rect 497657 381981 497663 382015
rect 497729 381981 497731 382015
rect 497765 381981 497767 382015
rect 497833 381981 497839 382015
rect 497901 381981 497911 382015
rect 497969 381981 497983 382015
rect 498037 381981 498055 382015
rect 498105 381981 498127 382015
rect 498173 381981 498199 382015
rect 498241 381981 498271 382015
rect 498309 381981 498343 382015
rect 498377 381981 498397 382015
rect 496838 381741 496898 381886
rect 496838 381707 496851 381741
rect 496885 381707 496898 381741
rect 496838 381341 496898 381707
rect 496838 381307 496851 381341
rect 496885 381307 496898 381341
rect 496838 380941 496898 381307
rect 496838 380907 496851 380941
rect 496885 380907 496898 380941
rect 496838 380746 496898 380907
rect 497018 381099 497058 381981
rect 498478 381557 498538 382439
rect 497099 381523 497119 381557
rect 497153 381523 497187 381557
rect 497225 381523 497255 381557
rect 497297 381523 497323 381557
rect 497369 381523 497391 381557
rect 497441 381523 497459 381557
rect 497513 381523 497527 381557
rect 497585 381523 497595 381557
rect 497657 381523 497663 381557
rect 497729 381523 497731 381557
rect 497765 381523 497767 381557
rect 497833 381523 497839 381557
rect 497901 381523 497911 381557
rect 497969 381523 497983 381557
rect 498037 381523 498055 381557
rect 498105 381523 498127 381557
rect 498173 381523 498199 381557
rect 498241 381523 498271 381557
rect 498309 381523 498343 381557
rect 498377 381523 498538 381557
rect 497018 381065 497119 381099
rect 497153 381065 497187 381099
rect 497225 381065 497255 381099
rect 497297 381065 497323 381099
rect 497369 381065 497391 381099
rect 497441 381065 497459 381099
rect 497513 381065 497527 381099
rect 497585 381065 497595 381099
rect 497657 381065 497663 381099
rect 497729 381065 497731 381099
rect 497765 381065 497767 381099
rect 497833 381065 497839 381099
rect 497901 381065 497911 381099
rect 497969 381065 497983 381099
rect 498037 381065 498055 381099
rect 498105 381065 498127 381099
rect 498173 381065 498199 381099
rect 498241 381065 498271 381099
rect 498309 381065 498343 381099
rect 498377 381065 498397 381099
rect 496838 380681 496978 380746
rect 496838 380647 496941 380681
rect 496975 380647 496978 380681
rect 496838 380586 496978 380647
rect 496838 380541 496898 380586
rect 496838 380507 496851 380541
rect 496885 380507 496898 380541
rect 496838 380141 496898 380507
rect 496838 380107 496851 380141
rect 496885 380107 496898 380141
rect 496838 379741 496898 380107
rect 496838 379707 496851 379741
rect 496885 379707 496898 379741
rect 496838 379446 496898 379707
rect 497018 380183 497058 381065
rect 498478 380641 498538 381523
rect 497099 380607 497119 380641
rect 497153 380607 497187 380641
rect 497225 380607 497255 380641
rect 497297 380607 497323 380641
rect 497369 380607 497391 380641
rect 497441 380607 497459 380641
rect 497513 380607 497527 380641
rect 497585 380607 497595 380641
rect 497657 380607 497663 380641
rect 497729 380607 497731 380641
rect 497765 380607 497767 380641
rect 497833 380607 497839 380641
rect 497901 380607 497911 380641
rect 497969 380607 497983 380641
rect 498037 380607 498055 380641
rect 498105 380607 498127 380641
rect 498173 380607 498199 380641
rect 498241 380607 498271 380641
rect 498309 380607 498343 380641
rect 498377 380607 498538 380641
rect 497018 380149 497119 380183
rect 497153 380149 497187 380183
rect 497225 380149 497255 380183
rect 497297 380149 497323 380183
rect 497369 380149 497391 380183
rect 497441 380149 497459 380183
rect 497513 380149 497527 380183
rect 497585 380149 497595 380183
rect 497657 380149 497663 380183
rect 497729 380149 497731 380183
rect 497765 380149 497767 380183
rect 497833 380149 497839 380183
rect 497901 380149 497911 380183
rect 497969 380149 497983 380183
rect 498037 380149 498055 380183
rect 498105 380149 498127 380183
rect 498173 380149 498199 380183
rect 498241 380149 498271 380183
rect 498309 380149 498343 380183
rect 498377 380149 498397 380183
rect 496838 379381 496978 379446
rect 496838 379347 496941 379381
rect 496975 379347 496978 379381
rect 496838 379341 496978 379347
rect 496838 379307 496851 379341
rect 496885 379307 496978 379341
rect 496838 379286 496978 379307
rect 496838 378941 496898 379286
rect 496838 378907 496851 378941
rect 496885 378907 496898 378941
rect 496838 378541 496898 378907
rect 496838 378507 496851 378541
rect 496885 378507 496898 378541
rect 496838 378146 496898 378507
rect 497018 379267 497058 380149
rect 498478 379725 498538 380607
rect 497099 379691 497119 379725
rect 497153 379691 497187 379725
rect 497225 379691 497255 379725
rect 497297 379691 497323 379725
rect 497369 379691 497391 379725
rect 497441 379691 497459 379725
rect 497513 379691 497527 379725
rect 497585 379691 497595 379725
rect 497657 379691 497663 379725
rect 497729 379691 497731 379725
rect 497765 379691 497767 379725
rect 497833 379691 497839 379725
rect 497901 379691 497911 379725
rect 497969 379691 497983 379725
rect 498037 379691 498055 379725
rect 498105 379691 498127 379725
rect 498173 379691 498199 379725
rect 498241 379691 498271 379725
rect 498309 379691 498343 379725
rect 498377 379691 498538 379725
rect 497018 379233 497119 379267
rect 497153 379233 497187 379267
rect 497225 379233 497255 379267
rect 497297 379233 497323 379267
rect 497369 379233 497391 379267
rect 497441 379233 497459 379267
rect 497513 379233 497527 379267
rect 497585 379233 497595 379267
rect 497657 379233 497663 379267
rect 497729 379233 497731 379267
rect 497765 379233 497767 379267
rect 497833 379233 497839 379267
rect 497901 379233 497911 379267
rect 497969 379233 497983 379267
rect 498037 379233 498055 379267
rect 498105 379233 498127 379267
rect 498173 379233 498199 379267
rect 498241 379233 498271 379267
rect 498309 379233 498343 379267
rect 498377 379233 498397 379267
rect 497018 378351 497058 379233
rect 498478 378809 498538 379691
rect 497099 378775 497119 378809
rect 497153 378775 497187 378809
rect 497225 378775 497255 378809
rect 497297 378775 497323 378809
rect 497369 378775 497391 378809
rect 497441 378775 497459 378809
rect 497513 378775 497527 378809
rect 497585 378775 497595 378809
rect 497657 378775 497663 378809
rect 497729 378775 497731 378809
rect 497765 378775 497767 378809
rect 497833 378775 497839 378809
rect 497901 378775 497911 378809
rect 497969 378775 497983 378809
rect 498037 378775 498055 378809
rect 498105 378775 498127 378809
rect 498173 378775 498199 378809
rect 498241 378775 498271 378809
rect 498309 378775 498343 378809
rect 498377 378775 498538 378809
rect 497018 378317 497119 378351
rect 497153 378317 497187 378351
rect 497225 378317 497255 378351
rect 497297 378317 497323 378351
rect 497369 378317 497391 378351
rect 497441 378317 497459 378351
rect 497513 378317 497527 378351
rect 497585 378317 497595 378351
rect 497657 378317 497663 378351
rect 497729 378317 497731 378351
rect 497765 378317 497767 378351
rect 497833 378317 497839 378351
rect 497901 378317 497911 378351
rect 497969 378317 497983 378351
rect 498037 378317 498055 378351
rect 498105 378317 498127 378351
rect 498173 378317 498199 378351
rect 498241 378317 498271 378351
rect 498309 378317 498343 378351
rect 498377 378317 498397 378351
rect 496838 378141 496978 378146
rect 496838 378107 496851 378141
rect 496885 378107 496978 378141
rect 496838 378081 496978 378107
rect 496838 378047 496941 378081
rect 496975 378047 496978 378081
rect 496838 377986 496978 378047
rect 496838 377741 496898 377986
rect 496838 377707 496851 377741
rect 496885 377707 496898 377741
rect 496838 377341 496898 377707
rect 496838 377307 496851 377341
rect 496885 377307 496898 377341
rect 496838 376941 496898 377307
rect 496838 376907 496851 376941
rect 496885 376907 496898 376941
rect 496838 376846 496898 376907
rect 497018 377435 497058 378317
rect 498478 377893 498538 378775
rect 497099 377859 497119 377893
rect 497153 377859 497187 377893
rect 497225 377859 497255 377893
rect 497297 377859 497323 377893
rect 497369 377859 497391 377893
rect 497441 377859 497459 377893
rect 497513 377859 497527 377893
rect 497585 377859 497595 377893
rect 497657 377859 497663 377893
rect 497729 377859 497731 377893
rect 497765 377859 497767 377893
rect 497833 377859 497839 377893
rect 497901 377859 497911 377893
rect 497969 377859 497983 377893
rect 498037 377859 498055 377893
rect 498105 377859 498127 377893
rect 498173 377859 498199 377893
rect 498241 377859 498271 377893
rect 498309 377859 498343 377893
rect 498377 377859 498538 377893
rect 497018 377401 497119 377435
rect 497153 377401 497187 377435
rect 497225 377401 497255 377435
rect 497297 377401 497323 377435
rect 497369 377401 497391 377435
rect 497441 377401 497459 377435
rect 497513 377401 497527 377435
rect 497585 377401 497595 377435
rect 497657 377401 497663 377435
rect 497729 377401 497731 377435
rect 497765 377401 497767 377435
rect 497833 377401 497839 377435
rect 497901 377401 497911 377435
rect 497969 377401 497983 377435
rect 498037 377401 498055 377435
rect 498105 377401 498127 377435
rect 498173 377401 498199 377435
rect 498241 377401 498271 377435
rect 498309 377401 498343 377435
rect 498377 377401 498397 377435
rect 496838 376781 496978 376846
rect 496838 376747 496941 376781
rect 496975 376747 496978 376781
rect 496838 376686 496978 376747
rect 496838 376541 496898 376686
rect 496838 376507 496851 376541
rect 496885 376507 496898 376541
rect 496838 376141 496898 376507
rect 496838 376107 496851 376141
rect 496885 376107 496898 376141
rect 496838 375741 496898 376107
rect 496838 375707 496851 375741
rect 496885 375707 496898 375741
rect 496838 375546 496898 375707
rect 497018 376519 497058 377401
rect 498478 376977 498538 377859
rect 497099 376943 497119 376977
rect 497153 376943 497187 376977
rect 497225 376943 497255 376977
rect 497297 376943 497323 376977
rect 497369 376943 497391 376977
rect 497441 376943 497459 376977
rect 497513 376943 497527 376977
rect 497585 376943 497595 376977
rect 497657 376943 497663 376977
rect 497729 376943 497731 376977
rect 497765 376943 497767 376977
rect 497833 376943 497839 376977
rect 497901 376943 497911 376977
rect 497969 376943 497983 376977
rect 498037 376943 498055 376977
rect 498105 376943 498127 376977
rect 498173 376943 498199 376977
rect 498241 376943 498271 376977
rect 498309 376943 498343 376977
rect 498377 376943 498538 376977
rect 497018 376485 497119 376519
rect 497153 376485 497187 376519
rect 497225 376485 497255 376519
rect 497297 376485 497323 376519
rect 497369 376485 497391 376519
rect 497441 376485 497459 376519
rect 497513 376485 497527 376519
rect 497585 376485 497595 376519
rect 497657 376485 497663 376519
rect 497729 376485 497731 376519
rect 497765 376485 497767 376519
rect 497833 376485 497839 376519
rect 497901 376485 497911 376519
rect 497969 376485 497983 376519
rect 498037 376485 498055 376519
rect 498105 376485 498127 376519
rect 498173 376485 498199 376519
rect 498241 376485 498271 376519
rect 498309 376485 498343 376519
rect 498377 376485 498397 376519
rect 497018 375603 497058 376485
rect 498478 376061 498538 376943
rect 497099 376027 497119 376061
rect 497153 376027 497187 376061
rect 497225 376027 497255 376061
rect 497297 376027 497323 376061
rect 497369 376027 497391 376061
rect 497441 376027 497459 376061
rect 497513 376027 497527 376061
rect 497585 376027 497595 376061
rect 497657 376027 497663 376061
rect 497729 376027 497731 376061
rect 497765 376027 497767 376061
rect 497833 376027 497839 376061
rect 497901 376027 497911 376061
rect 497969 376027 497983 376061
rect 498037 376027 498055 376061
rect 498105 376027 498127 376061
rect 498173 376027 498199 376061
rect 498241 376027 498271 376061
rect 498309 376027 498343 376061
rect 498377 376027 498538 376061
rect 497018 375569 497119 375603
rect 497153 375569 497187 375603
rect 497225 375569 497255 375603
rect 497297 375569 497323 375603
rect 497369 375569 497391 375603
rect 497441 375569 497459 375603
rect 497513 375569 497527 375603
rect 497585 375569 497595 375603
rect 497657 375569 497663 375603
rect 497729 375569 497731 375603
rect 497765 375569 497767 375603
rect 497833 375569 497839 375603
rect 497901 375569 497911 375603
rect 497969 375569 497983 375603
rect 498037 375569 498055 375603
rect 498105 375569 498127 375603
rect 498173 375569 498199 375603
rect 498241 375569 498271 375603
rect 498309 375569 498343 375603
rect 498377 375569 498397 375603
rect 496838 375481 496978 375546
rect 496838 375447 496941 375481
rect 496975 375447 496978 375481
rect 496838 375386 496978 375447
rect 496838 375341 496898 375386
rect 496838 375307 496851 375341
rect 496885 375307 496898 375341
rect 496838 374941 496898 375307
rect 496838 374907 496851 374941
rect 496885 374907 496898 374941
rect 496838 374541 496898 374907
rect 496838 374507 496851 374541
rect 496885 374507 496898 374541
rect 496838 374246 496898 374507
rect 497018 374687 497058 375569
rect 498478 375145 498538 376027
rect 497099 375111 497119 375145
rect 497153 375111 497187 375145
rect 497225 375111 497255 375145
rect 497297 375111 497323 375145
rect 497369 375111 497391 375145
rect 497441 375111 497459 375145
rect 497513 375111 497527 375145
rect 497585 375111 497595 375145
rect 497657 375111 497663 375145
rect 497729 375111 497731 375145
rect 497765 375111 497767 375145
rect 497833 375111 497839 375145
rect 497901 375111 497911 375145
rect 497969 375111 497983 375145
rect 498037 375111 498055 375145
rect 498105 375111 498127 375145
rect 498173 375111 498199 375145
rect 498241 375111 498271 375145
rect 498309 375111 498343 375145
rect 498377 375111 498538 375145
rect 497018 374653 497119 374687
rect 497153 374653 497187 374687
rect 497225 374653 497255 374687
rect 497297 374653 497323 374687
rect 497369 374653 497391 374687
rect 497441 374653 497459 374687
rect 497513 374653 497527 374687
rect 497585 374653 497595 374687
rect 497657 374653 497663 374687
rect 497729 374653 497731 374687
rect 497765 374653 497767 374687
rect 497833 374653 497839 374687
rect 497901 374653 497911 374687
rect 497969 374653 497983 374687
rect 498037 374653 498055 374687
rect 498105 374653 498127 374687
rect 498173 374653 498199 374687
rect 498241 374653 498271 374687
rect 498309 374653 498343 374687
rect 498377 374653 498397 374687
rect 496838 374181 496978 374246
rect 496838 374147 496941 374181
rect 496975 374147 496978 374181
rect 496838 374141 496978 374147
rect 496838 374107 496851 374141
rect 496885 374107 496978 374141
rect 496838 374086 496978 374107
rect 496838 373741 496898 374086
rect 496838 373707 496851 373741
rect 496885 373707 496898 373741
rect 496838 373341 496898 373707
rect 496838 373307 496851 373341
rect 496885 373307 496898 373341
rect 496838 372941 496898 373307
rect 496838 372907 496851 372941
rect 496885 372907 496898 372941
rect 496838 372541 496898 372907
rect 496838 372507 496851 372541
rect 496885 372507 496898 372541
rect 496838 372316 496898 372507
rect 497018 373771 497058 374653
rect 498478 374229 498538 375111
rect 497099 374195 497119 374229
rect 497153 374195 497187 374229
rect 497225 374195 497255 374229
rect 497297 374195 497323 374229
rect 497369 374195 497391 374229
rect 497441 374195 497459 374229
rect 497513 374195 497527 374229
rect 497585 374195 497595 374229
rect 497657 374195 497663 374229
rect 497729 374195 497731 374229
rect 497765 374195 497767 374229
rect 497833 374195 497839 374229
rect 497901 374195 497911 374229
rect 497969 374195 497983 374229
rect 498037 374195 498055 374229
rect 498105 374195 498127 374229
rect 498173 374195 498199 374229
rect 498241 374195 498271 374229
rect 498309 374195 498343 374229
rect 498377 374195 498538 374229
rect 497018 373737 497119 373771
rect 497153 373737 497187 373771
rect 497225 373737 497255 373771
rect 497297 373737 497323 373771
rect 497369 373737 497391 373771
rect 497441 373737 497459 373771
rect 497513 373737 497527 373771
rect 497585 373737 497595 373771
rect 497657 373737 497663 373771
rect 497729 373737 497731 373771
rect 497765 373737 497767 373771
rect 497833 373737 497839 373771
rect 497901 373737 497911 373771
rect 497969 373737 497983 373771
rect 498037 373737 498055 373771
rect 498105 373737 498127 373771
rect 498173 373737 498199 373771
rect 498241 373737 498271 373771
rect 498309 373737 498343 373771
rect 498377 373737 498397 373771
rect 497018 372855 497058 373737
rect 498478 373313 498538 374195
rect 497099 373279 497119 373313
rect 497153 373279 497187 373313
rect 497225 373279 497255 373313
rect 497297 373279 497323 373313
rect 497369 373279 497391 373313
rect 497441 373279 497459 373313
rect 497513 373279 497527 373313
rect 497585 373279 497595 373313
rect 497657 373279 497663 373313
rect 497729 373279 497731 373313
rect 497765 373279 497767 373313
rect 497833 373279 497839 373313
rect 497901 373279 497911 373313
rect 497969 373279 497983 373313
rect 498037 373279 498055 373313
rect 498105 373279 498127 373313
rect 498173 373279 498199 373313
rect 498241 373279 498271 373313
rect 498309 373279 498343 373313
rect 498377 373279 498538 373313
rect 497018 372821 497119 372855
rect 497153 372821 497187 372855
rect 497225 372821 497255 372855
rect 497297 372821 497323 372855
rect 497369 372821 497391 372855
rect 497441 372821 497459 372855
rect 497513 372821 497527 372855
rect 497585 372821 497595 372855
rect 497657 372821 497663 372855
rect 497729 372821 497731 372855
rect 497765 372821 497767 372855
rect 497833 372821 497839 372855
rect 497901 372821 497911 372855
rect 497969 372821 497983 372855
rect 498037 372821 498055 372855
rect 498105 372821 498127 372855
rect 498173 372821 498199 372855
rect 498241 372821 498271 372855
rect 498309 372821 498343 372855
rect 498377 372821 498397 372855
rect 497018 372316 497058 372821
rect 498478 372397 498538 373279
rect 497099 372363 497119 372397
rect 497153 372363 497187 372397
rect 497225 372363 497255 372397
rect 497297 372363 497323 372397
rect 497369 372363 497391 372397
rect 497441 372363 497459 372397
rect 497513 372363 497527 372397
rect 497585 372363 497595 372397
rect 497657 372363 497663 372397
rect 497729 372363 497731 372397
rect 497765 372363 497767 372397
rect 497833 372363 497839 372397
rect 497901 372363 497911 372397
rect 497969 372363 497983 372397
rect 498037 372363 498055 372397
rect 498105 372363 498127 372397
rect 498173 372363 498199 372397
rect 498241 372363 498271 372397
rect 498309 372363 498343 372397
rect 498377 372363 498538 372397
rect 498478 372316 498538 372363
rect 498584 399741 498644 399924
rect 498584 399707 498597 399741
rect 498631 399707 498644 399741
rect 498584 399341 498644 399707
rect 498584 399307 498597 399341
rect 498631 399307 498644 399341
rect 498584 398941 498644 399307
rect 498584 398907 498597 398941
rect 498631 398907 498644 398941
rect 498584 398541 498644 398907
rect 498584 398507 498597 398541
rect 498631 398507 498644 398541
rect 498584 398141 498644 398507
rect 498584 398107 498597 398141
rect 498631 398107 498644 398141
rect 498584 397741 498644 398107
rect 498584 397707 498597 397741
rect 498631 397707 498644 397741
rect 498584 397341 498644 397707
rect 498584 397307 498597 397341
rect 498631 397307 498644 397341
rect 498584 396941 498644 397307
rect 498584 396907 498597 396941
rect 498631 396907 498644 396941
rect 498584 396541 498644 396907
rect 498584 396507 498597 396541
rect 498631 396507 498644 396541
rect 498584 396141 498644 396507
rect 498584 396107 498597 396141
rect 498631 396107 498644 396141
rect 498584 395741 498644 396107
rect 498584 395707 498597 395741
rect 498631 395707 498644 395741
rect 498584 395341 498644 395707
rect 498584 395307 498597 395341
rect 498631 395307 498644 395341
rect 498584 394941 498644 395307
rect 498584 394907 498597 394941
rect 498631 394907 498644 394941
rect 498584 394541 498644 394907
rect 498584 394507 498597 394541
rect 498631 394507 498644 394541
rect 498584 394141 498644 394507
rect 498584 394107 498597 394141
rect 498631 394107 498644 394141
rect 498584 393741 498644 394107
rect 498584 393707 498597 393741
rect 498631 393707 498644 393741
rect 498584 393341 498644 393707
rect 498584 393307 498597 393341
rect 498631 393307 498644 393341
rect 498584 392941 498644 393307
rect 498584 392907 498597 392941
rect 498631 392907 498644 392941
rect 498584 392541 498644 392907
rect 498584 392507 498597 392541
rect 498631 392507 498644 392541
rect 498584 392141 498644 392507
rect 498584 392107 498597 392141
rect 498631 392107 498644 392141
rect 498584 391741 498644 392107
rect 498584 391707 498597 391741
rect 498631 391707 498644 391741
rect 498584 391341 498644 391707
rect 498584 391307 498597 391341
rect 498631 391307 498644 391341
rect 498584 390941 498644 391307
rect 498584 390907 498597 390941
rect 498631 390907 498644 390941
rect 498584 390541 498644 390907
rect 498584 390507 498597 390541
rect 498631 390507 498644 390541
rect 498584 390141 498644 390507
rect 498584 390107 498597 390141
rect 498631 390107 498644 390141
rect 498584 389741 498644 390107
rect 498584 389707 498597 389741
rect 498631 389707 498644 389741
rect 498584 389341 498644 389707
rect 498584 389307 498597 389341
rect 498631 389307 498644 389341
rect 498584 388941 498644 389307
rect 498584 388907 498597 388941
rect 498631 388907 498644 388941
rect 498584 388541 498644 388907
rect 498584 388507 498597 388541
rect 498631 388507 498644 388541
rect 498584 388141 498644 388507
rect 498584 388107 498597 388141
rect 498631 388107 498644 388141
rect 498584 387741 498644 388107
rect 498584 387707 498597 387741
rect 498631 387707 498644 387741
rect 498584 387341 498644 387707
rect 498584 387307 498597 387341
rect 498631 387307 498644 387341
rect 498584 386941 498644 387307
rect 498584 386907 498597 386941
rect 498631 386907 498644 386941
rect 498584 386541 498644 386907
rect 498584 386507 498597 386541
rect 498631 386507 498644 386541
rect 498584 386141 498644 386507
rect 498584 386107 498597 386141
rect 498631 386107 498644 386141
rect 498584 385741 498644 386107
rect 498584 385707 498597 385741
rect 498631 385707 498644 385741
rect 498584 385485 498644 385707
rect 498584 385451 498591 385485
rect 498625 385451 498644 385485
rect 498584 385341 498644 385451
rect 498584 385307 498597 385341
rect 498631 385307 498644 385341
rect 498584 384941 498644 385307
rect 498584 384907 498597 384941
rect 498631 384907 498644 384941
rect 498584 384541 498644 384907
rect 498584 384507 498597 384541
rect 498631 384507 498644 384541
rect 498584 384141 498644 384507
rect 498584 384107 498597 384141
rect 498631 384107 498644 384141
rect 498584 383741 498644 384107
rect 498584 383707 498597 383741
rect 498631 383707 498644 383741
rect 498584 383341 498644 383707
rect 498584 383307 498597 383341
rect 498631 383307 498644 383341
rect 498584 382941 498644 383307
rect 498584 382907 498597 382941
rect 498631 382907 498644 382941
rect 498584 382541 498644 382907
rect 498584 382507 498597 382541
rect 498631 382507 498644 382541
rect 498584 382141 498644 382507
rect 498584 382107 498597 382141
rect 498631 382107 498644 382141
rect 498584 381741 498644 382107
rect 498584 381707 498597 381741
rect 498631 381707 498644 381741
rect 498584 381341 498644 381707
rect 498584 381307 498597 381341
rect 498631 381307 498644 381341
rect 498584 380941 498644 381307
rect 498584 380907 498597 380941
rect 498631 380907 498644 380941
rect 498584 380541 498644 380907
rect 498584 380507 498597 380541
rect 498631 380507 498644 380541
rect 498584 380141 498644 380507
rect 498584 380107 498597 380141
rect 498631 380107 498644 380141
rect 498584 379741 498644 380107
rect 498584 379707 498597 379741
rect 498631 379707 498644 379741
rect 498584 379341 498644 379707
rect 498584 379307 498597 379341
rect 498631 379307 498644 379341
rect 498584 378941 498644 379307
rect 498584 378907 498597 378941
rect 498631 378907 498644 378941
rect 498584 378541 498644 378907
rect 498584 378507 498597 378541
rect 498631 378507 498644 378541
rect 498584 378141 498644 378507
rect 498584 378107 498597 378141
rect 498631 378107 498644 378141
rect 498584 377741 498644 378107
rect 498584 377707 498597 377741
rect 498631 377707 498644 377741
rect 498584 377341 498644 377707
rect 498584 377307 498597 377341
rect 498631 377307 498644 377341
rect 498584 376941 498644 377307
rect 498584 376907 498597 376941
rect 498631 376907 498644 376941
rect 498584 376541 498644 376907
rect 498584 376507 498597 376541
rect 498631 376507 498644 376541
rect 498584 376141 498644 376507
rect 498584 376107 498597 376141
rect 498631 376107 498644 376141
rect 498584 375741 498644 376107
rect 498584 375707 498597 375741
rect 498631 375707 498644 375741
rect 498584 375341 498644 375707
rect 498584 375307 498597 375341
rect 498631 375307 498644 375341
rect 498584 374941 498644 375307
rect 498584 374907 498597 374941
rect 498631 374907 498644 374941
rect 498584 374541 498644 374907
rect 498584 374507 498597 374541
rect 498631 374507 498644 374541
rect 498584 374141 498644 374507
rect 498584 374107 498597 374141
rect 498631 374107 498644 374141
rect 498584 373741 498644 374107
rect 498584 373707 498597 373741
rect 498631 373707 498644 373741
rect 498584 373341 498644 373707
rect 498584 373307 498597 373341
rect 498631 373307 498644 373341
rect 498584 372941 498644 373307
rect 498584 372907 498597 372941
rect 498631 372907 498644 372941
rect 498584 372541 498644 372907
rect 498584 372507 498597 372541
rect 498631 372507 498644 372541
rect 498584 372316 498644 372507
rect 498718 399741 498778 400022
rect 504358 399893 504418 400059
rect 504358 399859 504371 399893
rect 504405 399859 504418 399893
rect 498718 399707 498731 399741
rect 498765 399707 498778 399741
rect 498718 399341 498778 399707
rect 498718 399307 498731 399341
rect 498765 399307 498778 399341
rect 498718 398941 498778 399307
rect 498718 398907 498731 398941
rect 498765 398907 498778 398941
rect 498718 398541 498778 398907
rect 498718 398507 498731 398541
rect 498765 398507 498778 398541
rect 498718 398141 498778 398507
rect 498718 398107 498731 398141
rect 498765 398107 498778 398141
rect 498718 397741 498778 398107
rect 498718 397707 498731 397741
rect 498765 397707 498778 397741
rect 498718 397341 498778 397707
rect 498718 397307 498731 397341
rect 498765 397307 498778 397341
rect 498718 396941 498778 397307
rect 498718 396907 498731 396941
rect 498765 396907 498778 396941
rect 498718 396541 498778 396907
rect 498718 396507 498731 396541
rect 498765 396507 498778 396541
rect 498718 396141 498778 396507
rect 498718 396107 498731 396141
rect 498765 396107 498778 396141
rect 498718 395741 498778 396107
rect 498718 395707 498731 395741
rect 498765 395707 498778 395741
rect 498718 395341 498778 395707
rect 498718 395307 498731 395341
rect 498765 395307 498778 395341
rect 498718 394941 498778 395307
rect 498718 394907 498731 394941
rect 498765 394907 498778 394941
rect 498718 394541 498778 394907
rect 498718 394507 498731 394541
rect 498765 394507 498778 394541
rect 498718 394141 498778 394507
rect 498718 394107 498731 394141
rect 498765 394107 498778 394141
rect 498718 393741 498778 394107
rect 498718 393707 498731 393741
rect 498765 393707 498778 393741
rect 498718 393341 498778 393707
rect 498718 393307 498731 393341
rect 498765 393307 498778 393341
rect 498718 392941 498778 393307
rect 498718 392907 498731 392941
rect 498765 392907 498778 392941
rect 498718 392541 498778 392907
rect 500598 399641 500658 399824
rect 500598 399607 500611 399641
rect 500645 399607 500658 399641
rect 500598 399241 500658 399607
rect 500598 399207 500611 399241
rect 500645 399207 500658 399241
rect 500598 398841 500658 399207
rect 500598 398807 500611 398841
rect 500645 398807 500658 398841
rect 500598 398441 500658 398807
rect 500598 398407 500611 398441
rect 500645 398407 500658 398441
rect 500598 398041 500658 398407
rect 500598 398007 500611 398041
rect 500645 398007 500658 398041
rect 500598 397641 500658 398007
rect 500598 397607 500611 397641
rect 500645 397607 500658 397641
rect 500598 397241 500658 397607
rect 500598 397207 500611 397241
rect 500645 397207 500658 397241
rect 500598 396841 500658 397207
rect 500598 396807 500611 396841
rect 500645 396807 500658 396841
rect 500598 396441 500658 396807
rect 500598 396407 500611 396441
rect 500645 396407 500658 396441
rect 500598 396041 500658 396407
rect 500598 396007 500611 396041
rect 500645 396007 500658 396041
rect 500598 395641 500658 396007
rect 500598 395607 500611 395641
rect 500645 395607 500658 395641
rect 500598 395241 500658 395607
rect 500598 395207 500611 395241
rect 500645 395207 500658 395241
rect 500598 394841 500658 395207
rect 500598 394807 500611 394841
rect 500645 394807 500658 394841
rect 500598 394441 500658 394807
rect 500598 394407 500611 394441
rect 500645 394407 500658 394441
rect 500598 394041 500658 394407
rect 500598 394007 500611 394041
rect 500645 394007 500658 394041
rect 500598 393641 500658 394007
rect 500598 393607 500611 393641
rect 500645 393607 500658 393641
rect 500598 393241 500658 393607
rect 500598 393207 500611 393241
rect 500645 393207 500658 393241
rect 500598 392841 500658 393207
rect 500598 392807 500611 392841
rect 500645 392807 500658 392841
rect 500598 392656 500658 392807
rect 502478 399641 502538 399824
rect 502478 399607 502491 399641
rect 502525 399607 502538 399641
rect 502478 399241 502538 399607
rect 502478 399207 502491 399241
rect 502525 399207 502538 399241
rect 502478 398841 502538 399207
rect 502478 398807 502491 398841
rect 502525 398807 502538 398841
rect 504358 399693 504418 399859
rect 505298 400293 506298 400364
rect 505298 400277 506251 400293
rect 505298 399835 505337 400277
rect 505439 400259 506251 400277
rect 506285 400259 506298 400293
rect 505439 400093 506298 400259
rect 505439 400059 506251 400093
rect 506285 400059 506298 400093
rect 505439 399893 506298 400059
rect 505439 399859 506251 399893
rect 506285 399859 506298 399893
rect 505439 399835 506298 399859
rect 505298 399748 506298 399835
rect 504358 399659 504371 399693
rect 504405 399659 504418 399693
rect 504358 399493 504418 399659
rect 504358 399459 504371 399493
rect 504405 399459 504418 399493
rect 504358 399293 504418 399459
rect 504358 399259 504371 399293
rect 504405 399259 504418 399293
rect 506238 399693 506298 399748
rect 506238 399659 506251 399693
rect 506285 399659 506298 399693
rect 506238 399493 506298 399659
rect 506238 399459 506251 399493
rect 506285 399459 506298 399493
rect 506238 399293 506298 399459
rect 504358 399093 504418 399259
rect 504358 399059 504371 399093
rect 504405 399059 504418 399093
rect 504358 398836 504418 399059
rect 505193 398836 505583 399268
rect 506238 399259 506251 399293
rect 506285 399259 506298 399293
rect 506238 399093 506298 399259
rect 506238 399059 506251 399093
rect 506285 399059 506298 399093
rect 506238 398836 506298 399059
rect 502478 398441 502538 398807
rect 502478 398407 502491 398441
rect 502525 398407 502538 398441
rect 502478 398041 502538 398407
rect 502478 398007 502491 398041
rect 502525 398007 502538 398041
rect 502478 397641 502538 398007
rect 502478 397607 502491 397641
rect 502525 397607 502538 397641
rect 502478 397241 502538 397607
rect 502478 397207 502491 397241
rect 502525 397207 502538 397241
rect 502478 396841 502538 397207
rect 502478 396807 502491 396841
rect 502525 396807 502538 396841
rect 502478 396441 502538 396807
rect 502478 396407 502491 396441
rect 502525 396407 502538 396441
rect 502478 396041 502538 396407
rect 504358 398349 504418 398532
rect 504358 398315 504371 398349
rect 504405 398315 504418 398349
rect 504358 398149 504418 398315
rect 504358 398115 504371 398149
rect 504405 398115 504418 398149
rect 504358 397949 504418 398115
rect 506238 398349 506298 398532
rect 506238 398315 506251 398349
rect 506285 398315 506298 398349
rect 506238 398149 506298 398315
rect 506238 398115 506251 398149
rect 506285 398115 506298 398149
rect 504358 397915 504371 397949
rect 504405 397915 504418 397949
rect 504358 397749 504418 397915
rect 504358 397715 504371 397749
rect 504405 397715 504418 397749
rect 504358 397549 504418 397715
rect 506238 397949 506298 398115
rect 506238 397915 506251 397949
rect 506285 397915 506298 397949
rect 506238 397749 506298 397915
rect 506238 397715 506251 397749
rect 506285 397715 506298 397749
rect 506238 397620 506298 397715
rect 504358 397515 504371 397549
rect 504405 397515 504418 397549
rect 504358 397349 504418 397515
rect 504358 397315 504371 397349
rect 504405 397315 504418 397349
rect 504358 397149 504418 397315
rect 504358 397115 504371 397149
rect 504405 397115 504418 397149
rect 504358 396949 504418 397115
rect 505298 397549 506298 397620
rect 505298 397533 506251 397549
rect 505298 397091 505337 397533
rect 505439 397515 506251 397533
rect 506285 397515 506298 397549
rect 505439 397349 506298 397515
rect 505439 397315 506251 397349
rect 506285 397315 506298 397349
rect 505439 397149 506298 397315
rect 505439 397115 506251 397149
rect 506285 397115 506298 397149
rect 505439 397091 506298 397115
rect 505298 397004 506298 397091
rect 504358 396915 504371 396949
rect 504405 396915 504418 396949
rect 504358 396749 504418 396915
rect 504358 396715 504371 396749
rect 504405 396715 504418 396749
rect 504358 396549 504418 396715
rect 504358 396515 504371 396549
rect 504405 396515 504418 396549
rect 506238 396949 506298 397004
rect 506238 396915 506251 396949
rect 506285 396915 506298 396949
rect 506238 396749 506298 396915
rect 506238 396715 506251 396749
rect 506285 396715 506298 396749
rect 506238 396549 506298 396715
rect 504358 396349 504418 396515
rect 504358 396315 504371 396349
rect 504405 396315 504418 396349
rect 504358 396092 504418 396315
rect 505193 396092 505583 396524
rect 506238 396515 506251 396549
rect 506285 396515 506298 396549
rect 506238 396349 506298 396515
rect 506238 396315 506251 396349
rect 506285 396315 506298 396349
rect 506238 396092 506298 396315
rect 511878 398251 511938 398434
rect 511878 398217 511891 398251
rect 511925 398217 511938 398251
rect 511878 398051 511938 398217
rect 511878 398017 511891 398051
rect 511925 398017 511938 398051
rect 511878 397851 511938 398017
rect 513758 398251 513818 398434
rect 513758 398217 513771 398251
rect 513805 398217 513818 398251
rect 513758 398051 513818 398217
rect 513758 398017 513771 398051
rect 513805 398017 513818 398051
rect 511878 397817 511891 397851
rect 511925 397817 511938 397851
rect 511878 397651 511938 397817
rect 511878 397617 511891 397651
rect 511925 397617 511938 397651
rect 511878 397451 511938 397617
rect 513758 397851 513818 398017
rect 513758 397817 513771 397851
rect 513805 397817 513818 397851
rect 513758 397651 513818 397817
rect 513758 397617 513771 397651
rect 513805 397617 513818 397651
rect 513758 397522 513818 397617
rect 511878 397417 511891 397451
rect 511925 397417 511938 397451
rect 511878 397251 511938 397417
rect 511878 397217 511891 397251
rect 511925 397217 511938 397251
rect 511878 397051 511938 397217
rect 511878 397017 511891 397051
rect 511925 397017 511938 397051
rect 511878 396851 511938 397017
rect 512818 397451 513818 397522
rect 512818 397435 513771 397451
rect 512818 396993 512857 397435
rect 512959 397417 513771 397435
rect 513805 397417 513818 397451
rect 512959 397251 513818 397417
rect 512959 397217 513771 397251
rect 513805 397217 513818 397251
rect 512959 397051 513818 397217
rect 512959 397017 513771 397051
rect 513805 397017 513818 397051
rect 512959 396993 513818 397017
rect 512818 396906 513818 396993
rect 511878 396817 511891 396851
rect 511925 396817 511938 396851
rect 511878 396651 511938 396817
rect 511878 396617 511891 396651
rect 511925 396617 511938 396651
rect 511878 396451 511938 396617
rect 511878 396417 511891 396451
rect 511925 396417 511938 396451
rect 513758 396851 513818 396906
rect 513758 396817 513771 396851
rect 513805 396817 513818 396851
rect 513758 396651 513818 396817
rect 513758 396617 513771 396651
rect 513805 396617 513818 396651
rect 513758 396451 513818 396617
rect 511878 396251 511938 396417
rect 511878 396217 511891 396251
rect 511925 396217 511938 396251
rect 502478 396007 502491 396041
rect 502525 396007 502538 396041
rect 502478 395641 502538 396007
rect 511878 395994 511938 396217
rect 512713 395994 513103 396426
rect 513758 396417 513771 396451
rect 513805 396417 513818 396451
rect 513758 396251 513818 396417
rect 513758 396217 513771 396251
rect 513805 396217 513818 396251
rect 513758 395994 513818 396217
rect 502478 395607 502491 395641
rect 502525 395607 502538 395641
rect 502478 395241 502538 395607
rect 502478 395207 502491 395241
rect 502525 395207 502538 395241
rect 502478 394841 502538 395207
rect 502478 394807 502491 394841
rect 502525 394807 502538 394841
rect 502478 394441 502538 394807
rect 502478 394407 502491 394441
rect 502525 394407 502538 394441
rect 502478 394041 502538 394407
rect 502478 394007 502491 394041
rect 502525 394007 502538 394041
rect 502478 393641 502538 394007
rect 502478 393607 502491 393641
rect 502525 393607 502538 393641
rect 502478 393241 502538 393607
rect 502478 393207 502491 393241
rect 502525 393207 502538 393241
rect 502478 392841 502538 393207
rect 502478 392807 502491 392841
rect 502525 392807 502538 392841
rect 502478 392656 502538 392807
rect 504358 395603 504418 395786
rect 504358 395569 504371 395603
rect 504405 395569 504418 395603
rect 504358 395403 504418 395569
rect 504358 395369 504371 395403
rect 504405 395369 504418 395403
rect 504358 395203 504418 395369
rect 506238 395603 506298 395786
rect 506238 395569 506251 395603
rect 506285 395569 506298 395603
rect 506238 395403 506298 395569
rect 506238 395369 506251 395403
rect 506285 395369 506298 395403
rect 504358 395169 504371 395203
rect 504405 395169 504418 395203
rect 504358 395003 504418 395169
rect 504358 394969 504371 395003
rect 504405 394969 504418 395003
rect 504358 394803 504418 394969
rect 504358 394769 504371 394803
rect 504405 394769 504418 394803
rect 504358 394603 504418 394769
rect 504358 394569 504371 394603
rect 504405 394569 504418 394603
rect 506238 395203 506298 395369
rect 506238 395169 506251 395203
rect 506285 395169 506298 395203
rect 506238 395003 506298 395169
rect 506238 394969 506251 395003
rect 506285 394969 506298 395003
rect 506238 394803 506298 394969
rect 506238 394769 506251 394803
rect 506285 394769 506298 394803
rect 506238 394603 506298 394769
rect 506238 394588 506251 394603
rect 504358 394403 504418 394569
rect 504358 394369 504371 394403
rect 504405 394369 504418 394403
rect 504358 394203 504418 394369
rect 504358 394169 504371 394203
rect 504405 394169 504418 394203
rect 504358 394003 504418 394169
rect 504358 393969 504371 394003
rect 504405 393969 504418 394003
rect 505298 394569 506251 394588
rect 506285 394569 506298 394603
rect 505298 394501 506298 394569
rect 505298 394059 505337 394501
rect 505439 394403 506298 394501
rect 505439 394369 506251 394403
rect 506285 394369 506298 394403
rect 505439 394203 506298 394369
rect 505439 394169 506251 394203
rect 506285 394169 506298 394203
rect 505439 394059 506298 394169
rect 505298 394003 506298 394059
rect 505298 393972 506251 394003
rect 504358 393803 504418 393969
rect 504358 393769 504371 393803
rect 504405 393769 504418 393803
rect 504358 393603 504418 393769
rect 504358 393569 504371 393603
rect 504405 393569 504418 393603
rect 504358 393403 504418 393569
rect 504358 393369 504371 393403
rect 504405 393369 504418 393403
rect 504358 393203 504418 393369
rect 506238 393969 506251 393972
rect 506285 393969 506298 394003
rect 506238 393803 506298 393969
rect 506238 393769 506251 393803
rect 506285 393769 506298 393803
rect 506238 393603 506298 393769
rect 506238 393569 506251 393603
rect 506285 393569 506298 393603
rect 506238 393403 506298 393569
rect 506238 393369 506251 393403
rect 506285 393369 506298 393403
rect 504358 393169 504371 393203
rect 504405 393169 504418 393203
rect 504358 393003 504418 393169
rect 504358 392969 504371 393003
rect 504405 392969 504418 393003
rect 504358 392774 504418 392969
rect 505193 392773 505583 393205
rect 506238 393203 506298 393369
rect 508118 395507 508178 395690
rect 508118 395473 508131 395507
rect 508165 395473 508178 395507
rect 508118 395307 508178 395473
rect 508118 395273 508131 395307
rect 508165 395273 508178 395307
rect 508118 395107 508178 395273
rect 509998 395507 510058 395690
rect 509998 395473 510011 395507
rect 510045 395473 510058 395507
rect 509998 395307 510058 395473
rect 509998 395273 510011 395307
rect 510045 395273 510058 395307
rect 508118 395073 508131 395107
rect 508165 395073 508178 395107
rect 508118 394907 508178 395073
rect 508118 394873 508131 394907
rect 508165 394873 508178 394907
rect 508118 394707 508178 394873
rect 509998 395107 510058 395273
rect 509998 395073 510011 395107
rect 510045 395073 510058 395107
rect 509998 394907 510058 395073
rect 509998 394873 510011 394907
rect 510045 394873 510058 394907
rect 509998 394778 510058 394873
rect 508118 394673 508131 394707
rect 508165 394673 508178 394707
rect 508118 394507 508178 394673
rect 508118 394473 508131 394507
rect 508165 394473 508178 394507
rect 508118 394307 508178 394473
rect 508118 394273 508131 394307
rect 508165 394273 508178 394307
rect 508118 394107 508178 394273
rect 509058 394707 510058 394778
rect 509058 394691 510011 394707
rect 509058 394249 509097 394691
rect 509199 394673 510011 394691
rect 510045 394673 510058 394707
rect 509199 394507 510058 394673
rect 509199 394473 510011 394507
rect 510045 394473 510058 394507
rect 509199 394307 510058 394473
rect 509199 394273 510011 394307
rect 510045 394273 510058 394307
rect 509199 394249 510058 394273
rect 509058 394162 510058 394249
rect 508118 394073 508131 394107
rect 508165 394073 508178 394107
rect 508118 393907 508178 394073
rect 508118 393873 508131 393907
rect 508165 393873 508178 393907
rect 508118 393707 508178 393873
rect 508118 393673 508131 393707
rect 508165 393673 508178 393707
rect 509998 394107 510058 394162
rect 509998 394073 510011 394107
rect 510045 394073 510058 394107
rect 509998 393907 510058 394073
rect 509998 393873 510011 393907
rect 510045 393873 510058 393907
rect 509998 393707 510058 393873
rect 508118 393507 508178 393673
rect 508118 393473 508131 393507
rect 508165 393473 508178 393507
rect 508118 393250 508178 393473
rect 508953 393250 509343 393682
rect 509998 393673 510011 393707
rect 510045 393673 510058 393707
rect 509998 393507 510058 393673
rect 509998 393473 510011 393507
rect 510045 393473 510058 393507
rect 509998 393250 510058 393473
rect 511878 395507 511938 395690
rect 511878 395473 511891 395507
rect 511925 395473 511938 395507
rect 511878 395307 511938 395473
rect 511878 395273 511891 395307
rect 511925 395273 511938 395307
rect 511878 395107 511938 395273
rect 513758 395507 513818 395690
rect 513758 395473 513771 395507
rect 513805 395473 513818 395507
rect 513758 395307 513818 395473
rect 513758 395273 513771 395307
rect 513805 395273 513818 395307
rect 511878 395073 511891 395107
rect 511925 395073 511938 395107
rect 511878 394907 511938 395073
rect 511878 394873 511891 394907
rect 511925 394873 511938 394907
rect 511878 394707 511938 394873
rect 513758 395107 513818 395273
rect 513758 395073 513771 395107
rect 513805 395073 513818 395107
rect 513758 394907 513818 395073
rect 513758 394873 513771 394907
rect 513805 394873 513818 394907
rect 513758 394778 513818 394873
rect 511878 394673 511891 394707
rect 511925 394673 511938 394707
rect 511878 394507 511938 394673
rect 511878 394473 511891 394507
rect 511925 394473 511938 394507
rect 511878 394307 511938 394473
rect 511878 394273 511891 394307
rect 511925 394273 511938 394307
rect 511878 394107 511938 394273
rect 512818 394707 513818 394778
rect 512818 394691 513771 394707
rect 512818 394249 512857 394691
rect 512959 394673 513771 394691
rect 513805 394673 513818 394707
rect 512959 394507 513818 394673
rect 512959 394473 513771 394507
rect 513805 394473 513818 394507
rect 512959 394307 513818 394473
rect 512959 394273 513771 394307
rect 513805 394273 513818 394307
rect 512959 394249 513818 394273
rect 512818 394162 513818 394249
rect 511878 394073 511891 394107
rect 511925 394073 511938 394107
rect 511878 393907 511938 394073
rect 511878 393873 511891 393907
rect 511925 393873 511938 393907
rect 511878 393707 511938 393873
rect 511878 393673 511891 393707
rect 511925 393673 511938 393707
rect 513758 394107 513818 394162
rect 513758 394073 513771 394107
rect 513805 394073 513818 394107
rect 513758 393907 513818 394073
rect 513758 393873 513771 393907
rect 513805 393873 513818 393907
rect 513758 393707 513818 393873
rect 511878 393507 511938 393673
rect 511878 393473 511891 393507
rect 511925 393473 511938 393507
rect 511878 393250 511938 393473
rect 512713 393250 513103 393682
rect 513758 393673 513771 393707
rect 513805 393673 513818 393707
rect 513758 393507 513818 393673
rect 513758 393473 513771 393507
rect 513805 393473 513818 393507
rect 513758 393250 513818 393473
rect 506238 393169 506251 393203
rect 506285 393169 506298 393203
rect 506238 393003 506298 393169
rect 506238 392969 506251 393003
rect 506285 392969 506298 393003
rect 506238 392774 506298 392969
rect 508118 392761 508178 392944
rect 508118 392727 508131 392761
rect 508165 392727 508178 392761
rect 498718 392507 498731 392541
rect 498765 392507 498778 392541
rect 498718 392141 498778 392507
rect 508118 392561 508178 392727
rect 508118 392527 508131 392561
rect 508165 392527 508178 392561
rect 498718 392107 498731 392141
rect 498765 392107 498778 392141
rect 498718 391741 498778 392107
rect 498718 391707 498731 391741
rect 498765 391707 498778 391741
rect 498718 391341 498778 391707
rect 498718 391307 498731 391341
rect 498765 391307 498778 391341
rect 498718 390941 498778 391307
rect 498718 390907 498731 390941
rect 498765 390907 498778 390941
rect 498718 390541 498778 390907
rect 498718 390507 498731 390541
rect 498765 390507 498778 390541
rect 498718 390141 498778 390507
rect 498718 390107 498731 390141
rect 498765 390107 498778 390141
rect 498718 389741 498778 390107
rect 498718 389707 498731 389741
rect 498765 389707 498778 389741
rect 498718 389341 498778 389707
rect 498718 389307 498731 389341
rect 498765 389307 498778 389341
rect 498718 388941 498778 389307
rect 498718 388907 498731 388941
rect 498765 388907 498778 388941
rect 498718 388541 498778 388907
rect 498718 388507 498731 388541
rect 498765 388507 498778 388541
rect 498718 388141 498778 388507
rect 498718 388107 498731 388141
rect 498765 388107 498778 388141
rect 498718 387741 498778 388107
rect 498718 387707 498731 387741
rect 498765 387707 498778 387741
rect 498718 387341 498778 387707
rect 498718 387307 498731 387341
rect 498765 387307 498778 387341
rect 498718 386941 498778 387307
rect 498718 386907 498731 386941
rect 498765 386907 498778 386941
rect 498718 386541 498778 386907
rect 500598 392350 500658 392378
rect 500598 392337 500868 392350
rect 500598 392303 500751 392337
rect 500785 392303 500868 392337
rect 500598 392290 500868 392303
rect 500598 392097 500658 392290
rect 502238 392233 502298 392280
rect 500598 392063 500611 392097
rect 500645 392063 500658 392097
rect 500598 391697 500658 392063
rect 500598 391663 500611 391697
rect 500645 391663 500658 391697
rect 500598 391302 500658 391663
rect 500778 391775 500818 392220
rect 500859 392199 500879 392233
rect 500913 392199 500947 392233
rect 500985 392199 501015 392233
rect 501057 392199 501083 392233
rect 501129 392199 501151 392233
rect 501201 392199 501219 392233
rect 501273 392199 501287 392233
rect 501345 392199 501355 392233
rect 501417 392199 501423 392233
rect 501489 392199 501491 392233
rect 501525 392199 501527 392233
rect 501593 392199 501599 392233
rect 501661 392199 501671 392233
rect 501729 392199 501743 392233
rect 501797 392199 501815 392233
rect 501865 392199 501887 392233
rect 501933 392199 501959 392233
rect 502001 392199 502031 392233
rect 502069 392199 502103 392233
rect 502137 392201 502298 392233
rect 502137 392199 502229 392201
rect 502263 392167 502298 392201
rect 500778 391741 500879 391775
rect 500913 391741 500947 391775
rect 500985 391741 501015 391775
rect 501057 391741 501083 391775
rect 501129 391741 501151 391775
rect 501201 391741 501219 391775
rect 501273 391741 501287 391775
rect 501345 391741 501355 391775
rect 501417 391741 501423 391775
rect 501489 391741 501491 391775
rect 501525 391741 501527 391775
rect 501593 391741 501599 391775
rect 501661 391741 501671 391775
rect 501729 391741 501743 391775
rect 501797 391741 501815 391775
rect 501865 391741 501887 391775
rect 501933 391741 501959 391775
rect 502001 391741 502031 391775
rect 502069 391741 502103 391775
rect 502137 391741 502157 391775
rect 500598 391297 500738 391302
rect 500598 391263 500611 391297
rect 500645 391263 500738 391297
rect 500598 391237 500738 391263
rect 500598 391203 500701 391237
rect 500735 391203 500738 391237
rect 500598 391142 500738 391203
rect 500598 390897 500658 391142
rect 500598 390863 500611 390897
rect 500645 390863 500658 390897
rect 500598 390497 500658 390863
rect 500598 390463 500611 390497
rect 500645 390463 500658 390497
rect 500598 390097 500658 390463
rect 500598 390063 500611 390097
rect 500645 390063 500658 390097
rect 500598 390002 500658 390063
rect 500778 390859 500818 391741
rect 502238 391317 502298 392167
rect 500859 391283 500879 391317
rect 500913 391283 500947 391317
rect 500985 391283 501015 391317
rect 501057 391283 501083 391317
rect 501129 391283 501151 391317
rect 501201 391283 501219 391317
rect 501273 391283 501287 391317
rect 501345 391283 501355 391317
rect 501417 391283 501423 391317
rect 501489 391283 501491 391317
rect 501525 391283 501527 391317
rect 501593 391283 501599 391317
rect 501661 391283 501671 391317
rect 501729 391283 501743 391317
rect 501797 391283 501815 391317
rect 501865 391283 501887 391317
rect 501933 391283 501959 391317
rect 502001 391283 502031 391317
rect 502069 391283 502103 391317
rect 502137 391283 502298 391317
rect 500778 390825 500879 390859
rect 500913 390825 500947 390859
rect 500985 390825 501015 390859
rect 501057 390825 501083 390859
rect 501129 390825 501151 390859
rect 501201 390825 501219 390859
rect 501273 390825 501287 390859
rect 501345 390825 501355 390859
rect 501417 390825 501423 390859
rect 501489 390825 501491 390859
rect 501525 390825 501527 390859
rect 501593 390825 501599 390859
rect 501661 390825 501671 390859
rect 501729 390825 501743 390859
rect 501797 390825 501815 390859
rect 501865 390825 501887 390859
rect 501933 390825 501959 390859
rect 502001 390825 502031 390859
rect 502069 390825 502103 390859
rect 502137 390825 502157 390859
rect 500778 390085 500818 390825
rect 502238 390401 502298 391283
rect 500859 390367 500879 390401
rect 500913 390367 500947 390401
rect 500985 390367 501015 390401
rect 501057 390367 501083 390401
rect 501129 390367 501151 390401
rect 501201 390367 501219 390401
rect 501273 390367 501287 390401
rect 501345 390367 501355 390401
rect 501417 390367 501423 390401
rect 501489 390367 501491 390401
rect 501525 390367 501527 390401
rect 501593 390367 501599 390401
rect 501661 390367 501671 390401
rect 501729 390367 501743 390401
rect 501797 390367 501815 390401
rect 501865 390367 501887 390401
rect 501933 390367 501959 390401
rect 502001 390367 502031 390401
rect 502069 390367 502103 390401
rect 502137 390367 502298 390401
rect 500778 390051 500801 390085
rect 500598 389937 500738 390002
rect 500598 389903 500701 389937
rect 500735 389903 500738 389937
rect 500598 389842 500738 389903
rect 500778 389943 500818 390051
rect 500778 389909 500879 389943
rect 500913 389909 500947 389943
rect 500985 389909 501015 389943
rect 501057 389909 501083 389943
rect 501129 389909 501151 389943
rect 501201 389909 501219 389943
rect 501273 389909 501287 389943
rect 501345 389909 501355 389943
rect 501417 389909 501423 389943
rect 501489 389909 501491 389943
rect 501525 389909 501527 389943
rect 501593 389909 501599 389943
rect 501661 389909 501671 389943
rect 501729 389909 501743 389943
rect 501797 389909 501815 389943
rect 501865 389909 501887 389943
rect 501933 389909 501959 389943
rect 502001 389909 502031 389943
rect 502069 389909 502103 389943
rect 502137 389909 502157 389943
rect 500598 389697 500658 389842
rect 500598 389663 500611 389697
rect 500645 389663 500658 389697
rect 500598 389297 500658 389663
rect 500598 389263 500611 389297
rect 500645 389263 500658 389297
rect 500598 388897 500658 389263
rect 500598 388863 500611 388897
rect 500645 388863 500658 388897
rect 500598 388702 500658 388863
rect 500778 389027 500818 389909
rect 502238 389485 502298 390367
rect 500859 389451 500879 389485
rect 500913 389451 500947 389485
rect 500985 389451 501015 389485
rect 501057 389451 501083 389485
rect 501129 389451 501151 389485
rect 501201 389451 501219 389485
rect 501273 389451 501287 389485
rect 501345 389451 501355 389485
rect 501417 389451 501423 389485
rect 501489 389451 501491 389485
rect 501525 389451 501527 389485
rect 501593 389451 501599 389485
rect 501661 389451 501671 389485
rect 501729 389451 501743 389485
rect 501797 389451 501815 389485
rect 501865 389451 501887 389485
rect 501933 389451 501959 389485
rect 502001 389451 502031 389485
rect 502069 389451 502103 389485
rect 502137 389451 502298 389485
rect 500778 388993 500879 389027
rect 500913 388993 500947 389027
rect 500985 388993 501015 389027
rect 501057 388993 501083 389027
rect 501129 388993 501151 389027
rect 501201 388993 501219 389027
rect 501273 388993 501287 389027
rect 501345 388993 501355 389027
rect 501417 388993 501423 389027
rect 501489 388993 501491 389027
rect 501525 388993 501527 389027
rect 501593 388993 501599 389027
rect 501661 388993 501671 389027
rect 501729 388993 501743 389027
rect 501797 388993 501815 389027
rect 501865 388993 501887 389027
rect 501933 388993 501959 389027
rect 502001 388993 502031 389027
rect 502069 388993 502103 389027
rect 502137 388993 502157 389027
rect 500598 388637 500738 388702
rect 500598 388603 500701 388637
rect 500735 388603 500738 388637
rect 500598 388542 500738 388603
rect 500598 388497 500658 388542
rect 500598 388463 500611 388497
rect 500645 388463 500658 388497
rect 500598 388097 500658 388463
rect 500598 388063 500611 388097
rect 500645 388063 500658 388097
rect 500598 387697 500658 388063
rect 500598 387663 500611 387697
rect 500645 387663 500658 387697
rect 500598 387297 500658 387663
rect 500598 387263 500611 387297
rect 500645 387263 500658 387297
rect 500598 386897 500658 387263
rect 500598 386863 500611 386897
rect 500645 386863 500658 386897
rect 500598 386656 500658 386863
rect 500778 388111 500818 388993
rect 502238 388569 502298 389451
rect 500859 388535 500879 388569
rect 500913 388535 500947 388569
rect 500985 388535 501015 388569
rect 501057 388535 501083 388569
rect 501129 388535 501151 388569
rect 501201 388535 501219 388569
rect 501273 388535 501287 388569
rect 501345 388535 501355 388569
rect 501417 388535 501423 388569
rect 501489 388535 501491 388569
rect 501525 388535 501527 388569
rect 501593 388535 501599 388569
rect 501661 388535 501671 388569
rect 501729 388535 501743 388569
rect 501797 388535 501815 388569
rect 501865 388535 501887 388569
rect 501933 388535 501959 388569
rect 502001 388535 502031 388569
rect 502069 388535 502103 388569
rect 502137 388535 502298 388569
rect 500778 388077 500879 388111
rect 500913 388077 500947 388111
rect 500985 388077 501015 388111
rect 501057 388077 501083 388111
rect 501129 388077 501151 388111
rect 501201 388077 501219 388111
rect 501273 388077 501287 388111
rect 501345 388077 501355 388111
rect 501417 388077 501423 388111
rect 501489 388077 501491 388111
rect 501525 388077 501527 388111
rect 501593 388077 501599 388111
rect 501661 388077 501671 388111
rect 501729 388077 501743 388111
rect 501797 388077 501815 388111
rect 501865 388077 501887 388111
rect 501933 388077 501959 388111
rect 502001 388077 502031 388111
rect 502069 388077 502103 388111
rect 502137 388077 502157 388111
rect 500778 387195 500818 388077
rect 502238 387653 502298 388535
rect 500859 387619 500879 387653
rect 500913 387619 500947 387653
rect 500985 387619 501015 387653
rect 501057 387619 501083 387653
rect 501129 387619 501151 387653
rect 501201 387619 501219 387653
rect 501273 387619 501287 387653
rect 501345 387619 501355 387653
rect 501417 387619 501423 387653
rect 501489 387619 501491 387653
rect 501525 387619 501527 387653
rect 501593 387619 501599 387653
rect 501661 387619 501671 387653
rect 501729 387619 501743 387653
rect 501797 387619 501815 387653
rect 501865 387619 501887 387653
rect 501933 387619 501959 387653
rect 502001 387619 502031 387653
rect 502069 387619 502103 387653
rect 502137 387619 502298 387653
rect 500778 387161 500879 387195
rect 500913 387161 500947 387195
rect 500985 387161 501015 387195
rect 501057 387161 501083 387195
rect 501129 387161 501151 387195
rect 501201 387161 501219 387195
rect 501273 387161 501287 387195
rect 501345 387161 501355 387195
rect 501417 387161 501423 387195
rect 501489 387161 501491 387195
rect 501525 387161 501527 387195
rect 501593 387161 501599 387195
rect 501661 387161 501671 387195
rect 501729 387161 501743 387195
rect 501797 387161 501815 387195
rect 501865 387161 501887 387195
rect 501933 387161 501959 387195
rect 502001 387161 502031 387195
rect 502069 387161 502103 387195
rect 502137 387161 502157 387195
rect 500778 386656 500818 387161
rect 502238 386865 502298 387619
rect 502263 386831 502298 386865
rect 502238 386737 502298 386831
rect 500859 386703 500879 386737
rect 500913 386703 500947 386737
rect 500985 386703 501015 386737
rect 501057 386703 501083 386737
rect 501129 386703 501151 386737
rect 501201 386703 501219 386737
rect 501273 386703 501287 386737
rect 501345 386703 501355 386737
rect 501417 386703 501423 386737
rect 501489 386703 501491 386737
rect 501525 386703 501527 386737
rect 501593 386703 501599 386737
rect 501661 386703 501671 386737
rect 501729 386703 501743 386737
rect 501797 386703 501815 386737
rect 501865 386703 501887 386737
rect 501933 386703 501959 386737
rect 502001 386703 502031 386737
rect 502069 386703 502103 386737
rect 502137 386703 502298 386737
rect 502238 386656 502298 386703
rect 502344 392097 502404 392280
rect 502344 392063 502357 392097
rect 502391 392063 502404 392097
rect 502344 391697 502404 392063
rect 502344 391663 502357 391697
rect 502391 391663 502404 391697
rect 502344 391297 502404 391663
rect 502344 391263 502357 391297
rect 502391 391263 502404 391297
rect 502344 390897 502404 391263
rect 502344 390863 502357 390897
rect 502391 390863 502404 390897
rect 502344 390497 502404 390863
rect 502344 390463 502357 390497
rect 502391 390463 502404 390497
rect 502344 390097 502404 390463
rect 502344 390063 502357 390097
rect 502391 390063 502404 390097
rect 502344 389697 502404 390063
rect 502344 389663 502357 389697
rect 502391 389663 502404 389697
rect 502344 389297 502404 389663
rect 502344 389263 502357 389297
rect 502391 389263 502404 389297
rect 502344 388897 502404 389263
rect 502344 388863 502357 388897
rect 502391 388863 502404 388897
rect 502344 388497 502404 388863
rect 502344 388463 502357 388497
rect 502391 388463 502404 388497
rect 502344 388097 502404 388463
rect 502344 388063 502357 388097
rect 502391 388063 502404 388097
rect 502344 387697 502404 388063
rect 502344 387663 502357 387697
rect 502391 387663 502404 387697
rect 502344 387297 502404 387663
rect 502344 387263 502357 387297
rect 502391 387263 502404 387297
rect 502344 386897 502404 387263
rect 502344 386863 502357 386897
rect 502391 386863 502404 386897
rect 502344 386681 502404 386863
rect 502344 386656 502365 386681
rect 502399 386656 502404 386681
rect 502478 392097 502538 392378
rect 502478 392063 502491 392097
rect 502525 392063 502538 392097
rect 502478 391697 502538 392063
rect 502478 391663 502491 391697
rect 502525 391663 502538 391697
rect 502478 391297 502538 391663
rect 502478 391263 502491 391297
rect 502525 391263 502538 391297
rect 502478 390897 502538 391263
rect 502478 390863 502491 390897
rect 502525 390863 502538 390897
rect 502478 390497 502538 390863
rect 502478 390463 502491 390497
rect 502525 390463 502538 390497
rect 502478 390097 502538 390463
rect 502478 390063 502491 390097
rect 502525 390063 502538 390097
rect 502478 389697 502538 390063
rect 504358 392273 504418 392456
rect 504358 392239 504371 392273
rect 504405 392239 504418 392273
rect 504358 392073 504418 392239
rect 504358 392039 504371 392073
rect 504405 392039 504418 392073
rect 504358 391873 504418 392039
rect 506238 392273 506298 392456
rect 506238 392239 506251 392273
rect 506285 392239 506298 392273
rect 506238 392073 506298 392239
rect 506238 392039 506251 392073
rect 506285 392039 506298 392073
rect 504358 391839 504371 391873
rect 504405 391839 504418 391873
rect 504358 391673 504418 391839
rect 504358 391639 504371 391673
rect 504405 391639 504418 391673
rect 504358 391473 504418 391639
rect 506238 391873 506298 392039
rect 506238 391839 506251 391873
rect 506285 391839 506298 391873
rect 506238 391673 506298 391839
rect 506238 391639 506251 391673
rect 506285 391639 506298 391673
rect 506238 391544 506298 391639
rect 504358 391439 504371 391473
rect 504405 391439 504418 391473
rect 504358 391273 504418 391439
rect 504358 391239 504371 391273
rect 504405 391239 504418 391273
rect 504358 391073 504418 391239
rect 504358 391039 504371 391073
rect 504405 391039 504418 391073
rect 504358 390873 504418 391039
rect 505298 391473 506298 391544
rect 505298 391457 506251 391473
rect 505298 391015 505337 391457
rect 505439 391439 506251 391457
rect 506285 391439 506298 391473
rect 505439 391273 506298 391439
rect 505439 391239 506251 391273
rect 506285 391239 506298 391273
rect 505439 391073 506298 391239
rect 505439 391039 506251 391073
rect 506285 391039 506298 391073
rect 505439 391015 506298 391039
rect 505298 390928 506298 391015
rect 504358 390839 504371 390873
rect 504405 390839 504418 390873
rect 504358 390673 504418 390839
rect 504358 390639 504371 390673
rect 504405 390639 504418 390673
rect 504358 390473 504418 390639
rect 504358 390439 504371 390473
rect 504405 390439 504418 390473
rect 506238 390873 506298 390928
rect 506238 390839 506251 390873
rect 506285 390839 506298 390873
rect 506238 390673 506298 390839
rect 506238 390639 506251 390673
rect 506285 390639 506298 390673
rect 506238 390473 506298 390639
rect 504358 390273 504418 390439
rect 504358 390239 504371 390273
rect 504405 390239 504418 390273
rect 504358 390016 504418 390239
rect 505193 390016 505583 390448
rect 506238 390439 506251 390473
rect 506285 390439 506298 390473
rect 506238 390273 506298 390439
rect 506238 390239 506251 390273
rect 506285 390239 506298 390273
rect 506238 390016 506298 390239
rect 508118 392361 508178 392527
rect 509998 392761 510058 392944
rect 509998 392727 510011 392761
rect 510045 392727 510058 392761
rect 509998 392561 510058 392727
rect 509998 392527 510011 392561
rect 510045 392527 510058 392561
rect 508118 392327 508131 392361
rect 508165 392327 508178 392361
rect 508118 392161 508178 392327
rect 508118 392127 508131 392161
rect 508165 392127 508178 392161
rect 508118 391961 508178 392127
rect 508118 391927 508131 391961
rect 508165 391927 508178 391961
rect 508118 391761 508178 391927
rect 508118 391727 508131 391761
rect 508165 391727 508178 391761
rect 509998 392361 510058 392527
rect 509998 392327 510011 392361
rect 510045 392327 510058 392361
rect 509998 392161 510058 392327
rect 509998 392127 510011 392161
rect 510045 392127 510058 392161
rect 509998 391961 510058 392127
rect 509998 391927 510011 391961
rect 510045 391927 510058 391961
rect 509998 391761 510058 391927
rect 509998 391746 510011 391761
rect 508118 391561 508178 391727
rect 508118 391527 508131 391561
rect 508165 391527 508178 391561
rect 508118 391361 508178 391527
rect 508118 391327 508131 391361
rect 508165 391327 508178 391361
rect 508118 391161 508178 391327
rect 508118 391127 508131 391161
rect 508165 391127 508178 391161
rect 509058 391727 510011 391746
rect 510045 391727 510058 391761
rect 509058 391659 510058 391727
rect 509058 391217 509097 391659
rect 509199 391561 510058 391659
rect 509199 391527 510011 391561
rect 510045 391527 510058 391561
rect 509199 391361 510058 391527
rect 509199 391327 510011 391361
rect 510045 391327 510058 391361
rect 509199 391217 510058 391327
rect 509058 391161 510058 391217
rect 509058 391130 510011 391161
rect 508118 390961 508178 391127
rect 508118 390927 508131 390961
rect 508165 390927 508178 390961
rect 508118 390761 508178 390927
rect 508118 390727 508131 390761
rect 508165 390727 508178 390761
rect 508118 390561 508178 390727
rect 508118 390527 508131 390561
rect 508165 390527 508178 390561
rect 508118 390361 508178 390527
rect 509998 391127 510011 391130
rect 510045 391127 510058 391161
rect 509998 390961 510058 391127
rect 509998 390927 510011 390961
rect 510045 390927 510058 390961
rect 509998 390761 510058 390927
rect 509998 390727 510011 390761
rect 510045 390727 510058 390761
rect 509998 390561 510058 390727
rect 509998 390527 510011 390561
rect 510045 390527 510058 390561
rect 508118 390327 508131 390361
rect 508165 390327 508178 390361
rect 508118 390161 508178 390327
rect 508118 390127 508131 390161
rect 508165 390127 508178 390161
rect 508118 389932 508178 390127
rect 508953 389931 509343 390363
rect 509998 390361 510058 390527
rect 511878 392763 511938 392946
rect 511878 392729 511891 392763
rect 511925 392729 511938 392763
rect 511878 392563 511938 392729
rect 511878 392529 511891 392563
rect 511925 392529 511938 392563
rect 511878 392363 511938 392529
rect 513758 392763 513818 392946
rect 513758 392729 513771 392763
rect 513805 392729 513818 392763
rect 513758 392563 513818 392729
rect 513758 392529 513771 392563
rect 513805 392529 513818 392563
rect 511878 392329 511891 392363
rect 511925 392329 511938 392363
rect 511878 392163 511938 392329
rect 511878 392129 511891 392163
rect 511925 392129 511938 392163
rect 511878 391963 511938 392129
rect 513758 392363 513818 392529
rect 513758 392329 513771 392363
rect 513805 392329 513818 392363
rect 513758 392163 513818 392329
rect 513758 392129 513771 392163
rect 513805 392129 513818 392163
rect 513758 392034 513818 392129
rect 511878 391929 511891 391963
rect 511925 391929 511938 391963
rect 511878 391763 511938 391929
rect 511878 391729 511891 391763
rect 511925 391729 511938 391763
rect 511878 391563 511938 391729
rect 511878 391529 511891 391563
rect 511925 391529 511938 391563
rect 511878 391363 511938 391529
rect 512818 391963 513818 392034
rect 512818 391947 513771 391963
rect 512818 391505 512857 391947
rect 512959 391929 513771 391947
rect 513805 391929 513818 391963
rect 512959 391763 513818 391929
rect 512959 391729 513771 391763
rect 513805 391729 513818 391763
rect 512959 391563 513818 391729
rect 512959 391529 513771 391563
rect 513805 391529 513818 391563
rect 512959 391505 513818 391529
rect 512818 391418 513818 391505
rect 511878 391329 511891 391363
rect 511925 391329 511938 391363
rect 511878 391163 511938 391329
rect 511878 391129 511891 391163
rect 511925 391129 511938 391163
rect 511878 390963 511938 391129
rect 511878 390929 511891 390963
rect 511925 390929 511938 390963
rect 513758 391363 513818 391418
rect 513758 391329 513771 391363
rect 513805 391329 513818 391363
rect 513758 391163 513818 391329
rect 513758 391129 513771 391163
rect 513805 391129 513818 391163
rect 513758 390963 513818 391129
rect 511878 390763 511938 390929
rect 511878 390729 511891 390763
rect 511925 390729 511938 390763
rect 511878 390506 511938 390729
rect 512713 390506 513103 390938
rect 513758 390929 513771 390963
rect 513805 390929 513818 390963
rect 513758 390763 513818 390929
rect 513758 390729 513771 390763
rect 513805 390729 513818 390763
rect 513758 390506 513818 390729
rect 515638 392371 515698 392554
rect 515638 392337 515651 392371
rect 515685 392337 515698 392371
rect 515638 392171 515698 392337
rect 515638 392137 515651 392171
rect 515685 392137 515698 392171
rect 515638 391971 515698 392137
rect 517518 392371 517578 392554
rect 517518 392337 517531 392371
rect 517565 392337 517578 392371
rect 517518 392171 517578 392337
rect 517518 392137 517531 392171
rect 517565 392137 517578 392171
rect 515638 391937 515651 391971
rect 515685 391937 515698 391971
rect 515638 391771 515698 391937
rect 515638 391737 515651 391771
rect 515685 391737 515698 391771
rect 515638 391571 515698 391737
rect 517518 391971 517578 392137
rect 517518 391937 517531 391971
rect 517565 391937 517578 391971
rect 517518 391771 517578 391937
rect 517518 391737 517531 391771
rect 517565 391737 517578 391771
rect 517518 391642 517578 391737
rect 515638 391537 515651 391571
rect 515685 391537 515698 391571
rect 515638 391371 515698 391537
rect 515638 391337 515651 391371
rect 515685 391337 515698 391371
rect 515638 391171 515698 391337
rect 515638 391137 515651 391171
rect 515685 391137 515698 391171
rect 515638 390971 515698 391137
rect 516578 391571 517578 391642
rect 516578 391555 517531 391571
rect 516578 391113 516617 391555
rect 516719 391537 517531 391555
rect 517565 391537 517578 391571
rect 516719 391371 517578 391537
rect 516719 391337 517531 391371
rect 517565 391337 517578 391371
rect 516719 391171 517578 391337
rect 516719 391137 517531 391171
rect 517565 391137 517578 391171
rect 516719 391113 517578 391137
rect 516578 391026 517578 391113
rect 515638 390937 515651 390971
rect 515685 390937 515698 390971
rect 515638 390771 515698 390937
rect 515638 390737 515651 390771
rect 515685 390737 515698 390771
rect 515638 390571 515698 390737
rect 515638 390537 515651 390571
rect 515685 390537 515698 390571
rect 517518 390971 517578 391026
rect 517518 390937 517531 390971
rect 517565 390937 517578 390971
rect 517518 390771 517578 390937
rect 517518 390737 517531 390771
rect 517565 390737 517578 390771
rect 517518 390571 517578 390737
rect 509998 390327 510011 390361
rect 510045 390327 510058 390361
rect 509998 390161 510058 390327
rect 509998 390127 510011 390161
rect 510045 390127 510058 390161
rect 509998 389932 510058 390127
rect 515638 390371 515698 390537
rect 515638 390337 515651 390371
rect 515685 390337 515698 390371
rect 515638 390114 515698 390337
rect 516473 390114 516863 390546
rect 517518 390537 517531 390571
rect 517565 390537 517578 390571
rect 517518 390371 517578 390537
rect 517518 390337 517531 390371
rect 517565 390337 517578 390371
rect 517518 390114 517578 390337
rect 519398 390901 519458 391084
rect 519398 390867 519411 390901
rect 519445 390867 519458 390901
rect 519398 390701 519458 390867
rect 519398 390667 519411 390701
rect 519445 390667 519458 390701
rect 519398 390501 519458 390667
rect 521278 390901 521338 391084
rect 521278 390867 521291 390901
rect 521325 390867 521338 390901
rect 521278 390701 521338 390867
rect 521278 390667 521291 390701
rect 521325 390667 521338 390701
rect 519398 390467 519411 390501
rect 519445 390467 519458 390501
rect 519398 390301 519458 390467
rect 519398 390267 519411 390301
rect 519445 390267 519458 390301
rect 519398 390101 519458 390267
rect 521278 390501 521338 390667
rect 521278 390467 521291 390501
rect 521325 390467 521338 390501
rect 521278 390301 521338 390467
rect 521278 390267 521291 390301
rect 521325 390267 521338 390301
rect 521278 390172 521338 390267
rect 519398 390067 519411 390101
rect 519445 390067 519458 390101
rect 502478 389663 502491 389697
rect 502525 389663 502538 389697
rect 502478 389297 502538 389663
rect 519398 389901 519458 390067
rect 519398 389867 519411 389901
rect 519445 389867 519458 389901
rect 519398 389701 519458 389867
rect 519398 389667 519411 389701
rect 519445 389667 519458 389701
rect 502478 389263 502491 389297
rect 502525 389263 502538 389297
rect 502478 388897 502538 389263
rect 502478 388863 502491 388897
rect 502525 388863 502538 388897
rect 502478 388497 502538 388863
rect 502478 388463 502491 388497
rect 502525 388463 502538 388497
rect 502478 388097 502538 388463
rect 502478 388063 502491 388097
rect 502525 388063 502538 388097
rect 502478 387697 502538 388063
rect 502478 387663 502491 387697
rect 502525 387663 502538 387697
rect 502478 387297 502538 387663
rect 502478 387263 502491 387297
rect 502525 387263 502538 387297
rect 502478 386897 502538 387263
rect 502478 386863 502491 386897
rect 502525 386863 502538 386897
rect 502478 386656 502538 386863
rect 504358 389353 504418 389634
rect 506238 389606 506298 389634
rect 506028 389593 506298 389606
rect 506028 389559 506111 389593
rect 506145 389559 506298 389593
rect 506028 389546 506298 389559
rect 504358 389319 504371 389353
rect 504405 389319 504418 389353
rect 504358 388953 504418 389319
rect 504358 388919 504371 388953
rect 504405 388919 504418 388953
rect 504358 388553 504418 388919
rect 504358 388519 504371 388553
rect 504405 388519 504418 388553
rect 504358 388153 504418 388519
rect 504358 388119 504371 388153
rect 504405 388119 504418 388153
rect 504358 387753 504418 388119
rect 504358 387719 504371 387753
rect 504405 387719 504418 387753
rect 504358 387353 504418 387719
rect 504358 387319 504371 387353
rect 504405 387319 504418 387353
rect 504358 386953 504418 387319
rect 504358 386919 504371 386953
rect 504405 386919 504418 386953
rect 498718 386507 498731 386541
rect 498765 386507 498778 386541
rect 498718 386141 498778 386507
rect 498718 386107 498731 386141
rect 498765 386107 498778 386141
rect 498718 385741 498778 386107
rect 498718 385707 498731 385741
rect 498765 385707 498778 385741
rect 504358 386553 504418 386919
rect 504358 386519 504371 386553
rect 504405 386519 504418 386553
rect 504358 386153 504418 386519
rect 504358 386119 504371 386153
rect 504405 386119 504418 386153
rect 504358 385753 504418 386119
rect 504358 385719 504371 385753
rect 504405 385719 504418 385753
rect 498718 385341 498778 385707
rect 498718 385307 498731 385341
rect 498765 385307 498778 385341
rect 498718 384941 498778 385307
rect 498718 384907 498731 384941
rect 498765 384907 498778 384941
rect 498718 384541 498778 384907
rect 498718 384507 498731 384541
rect 498765 384507 498778 384541
rect 498718 384141 498778 384507
rect 498718 384107 498731 384141
rect 498765 384107 498778 384141
rect 498718 383741 498778 384107
rect 498718 383707 498731 383741
rect 498765 383707 498778 383741
rect 498718 383341 498778 383707
rect 498718 383307 498731 383341
rect 498765 383307 498778 383341
rect 498718 382941 498778 383307
rect 498718 382907 498731 382941
rect 498765 382907 498778 382941
rect 498718 382541 498778 382907
rect 498718 382507 498731 382541
rect 498765 382507 498778 382541
rect 498718 382141 498778 382507
rect 498718 382107 498731 382141
rect 498765 382107 498778 382141
rect 498718 381741 498778 382107
rect 498718 381707 498731 381741
rect 498765 381707 498778 381741
rect 498718 381341 498778 381707
rect 498718 381307 498731 381341
rect 498765 381307 498778 381341
rect 498718 380941 498778 381307
rect 498718 380907 498731 380941
rect 498765 380907 498778 380941
rect 498718 380541 498778 380907
rect 498718 380507 498731 380541
rect 498765 380507 498778 380541
rect 498718 380141 498778 380507
rect 498718 380107 498731 380141
rect 498765 380107 498778 380141
rect 498718 379741 498778 380107
rect 500598 385686 500658 385714
rect 500598 385673 500868 385686
rect 500598 385639 500751 385673
rect 500785 385639 500868 385673
rect 500598 385626 500868 385639
rect 500598 385433 500658 385626
rect 502238 385569 502298 385616
rect 500598 385399 500611 385433
rect 500645 385399 500658 385433
rect 500598 385033 500658 385399
rect 500598 384999 500611 385033
rect 500645 384999 500658 385033
rect 500598 384638 500658 384999
rect 500778 385111 500818 385556
rect 500859 385535 500879 385569
rect 500913 385535 500947 385569
rect 500985 385535 501015 385569
rect 501057 385535 501083 385569
rect 501129 385535 501151 385569
rect 501201 385535 501219 385569
rect 501273 385535 501287 385569
rect 501345 385535 501355 385569
rect 501417 385535 501423 385569
rect 501489 385535 501491 385569
rect 501525 385535 501527 385569
rect 501593 385535 501599 385569
rect 501661 385535 501671 385569
rect 501729 385535 501743 385569
rect 501797 385535 501815 385569
rect 501865 385535 501887 385569
rect 501933 385535 501959 385569
rect 502001 385535 502031 385569
rect 502069 385535 502103 385569
rect 502137 385535 502298 385569
rect 500778 385077 500879 385111
rect 500913 385077 500947 385111
rect 500985 385077 501015 385111
rect 501057 385077 501083 385111
rect 501129 385077 501151 385111
rect 501201 385077 501219 385111
rect 501273 385077 501287 385111
rect 501345 385077 501355 385111
rect 501417 385077 501423 385111
rect 501489 385077 501491 385111
rect 501525 385077 501527 385111
rect 501593 385077 501599 385111
rect 501661 385077 501671 385111
rect 501729 385077 501743 385111
rect 501797 385077 501815 385111
rect 501865 385077 501887 385111
rect 501933 385077 501959 385111
rect 502001 385077 502031 385111
rect 502069 385077 502103 385111
rect 502137 385077 502157 385111
rect 500598 384633 500738 384638
rect 500598 384599 500611 384633
rect 500645 384599 500738 384633
rect 500598 384573 500738 384599
rect 500598 384539 500701 384573
rect 500735 384539 500738 384573
rect 500598 384478 500738 384539
rect 500598 384233 500658 384478
rect 500598 384199 500611 384233
rect 500645 384199 500658 384233
rect 500598 383833 500658 384199
rect 500598 383799 500611 383833
rect 500645 383799 500658 383833
rect 500598 383433 500658 383799
rect 500598 383399 500611 383433
rect 500645 383399 500658 383433
rect 500598 383338 500658 383399
rect 500778 384195 500818 385077
rect 502238 384653 502298 385535
rect 500859 384619 500879 384653
rect 500913 384619 500947 384653
rect 500985 384619 501015 384653
rect 501057 384619 501083 384653
rect 501129 384619 501151 384653
rect 501201 384619 501219 384653
rect 501273 384619 501287 384653
rect 501345 384619 501355 384653
rect 501417 384619 501423 384653
rect 501489 384619 501491 384653
rect 501525 384619 501527 384653
rect 501593 384619 501599 384653
rect 501661 384619 501671 384653
rect 501729 384619 501743 384653
rect 501797 384619 501815 384653
rect 501865 384619 501887 384653
rect 501933 384619 501959 384653
rect 502001 384619 502031 384653
rect 502069 384619 502103 384653
rect 502137 384619 502298 384653
rect 500778 384161 500879 384195
rect 500913 384161 500947 384195
rect 500985 384161 501015 384195
rect 501057 384161 501083 384195
rect 501129 384161 501151 384195
rect 501201 384161 501219 384195
rect 501273 384161 501287 384195
rect 501345 384161 501355 384195
rect 501417 384161 501423 384195
rect 501489 384161 501491 384195
rect 501525 384161 501527 384195
rect 501593 384161 501599 384195
rect 501661 384161 501671 384195
rect 501729 384161 501743 384195
rect 501797 384161 501815 384195
rect 501865 384161 501887 384195
rect 501933 384161 501959 384195
rect 502001 384161 502031 384195
rect 502069 384161 502103 384195
rect 502137 384161 502157 384195
rect 500598 383273 500738 383338
rect 500598 383239 500701 383273
rect 500735 383239 500738 383273
rect 500598 383178 500738 383239
rect 500778 383279 500818 384161
rect 502238 383737 502298 384619
rect 500859 383703 500879 383737
rect 500913 383703 500947 383737
rect 500985 383703 501015 383737
rect 501057 383703 501083 383737
rect 501129 383703 501151 383737
rect 501201 383703 501219 383737
rect 501273 383703 501287 383737
rect 501345 383703 501355 383737
rect 501417 383703 501423 383737
rect 501489 383703 501491 383737
rect 501525 383703 501527 383737
rect 501593 383703 501599 383737
rect 501661 383703 501671 383737
rect 501729 383703 501743 383737
rect 501797 383703 501815 383737
rect 501865 383703 501887 383737
rect 501933 383703 501959 383737
rect 502001 383703 502031 383737
rect 502069 383703 502103 383737
rect 502137 383703 502298 383737
rect 500778 383245 500879 383279
rect 500913 383245 500947 383279
rect 500985 383245 501015 383279
rect 501057 383245 501083 383279
rect 501129 383245 501151 383279
rect 501201 383245 501219 383279
rect 501273 383245 501287 383279
rect 501345 383245 501355 383279
rect 501417 383245 501423 383279
rect 501489 383245 501491 383279
rect 501525 383245 501527 383279
rect 501593 383245 501599 383279
rect 501661 383245 501671 383279
rect 501729 383245 501743 383279
rect 501797 383245 501815 383279
rect 501865 383245 501887 383279
rect 501933 383245 501959 383279
rect 502001 383245 502031 383279
rect 502069 383245 502103 383279
rect 502137 383245 502157 383279
rect 500598 383033 500658 383178
rect 500598 382999 500611 383033
rect 500645 382999 500658 383033
rect 500598 382633 500658 382999
rect 500598 382599 500611 382633
rect 500645 382599 500658 382633
rect 500598 382233 500658 382599
rect 500598 382199 500611 382233
rect 500645 382199 500658 382233
rect 500598 382038 500658 382199
rect 500778 382363 500818 383245
rect 502238 382821 502298 383703
rect 500859 382787 500879 382821
rect 500913 382787 500947 382821
rect 500985 382787 501015 382821
rect 501057 382787 501083 382821
rect 501129 382787 501151 382821
rect 501201 382787 501219 382821
rect 501273 382787 501287 382821
rect 501345 382787 501355 382821
rect 501417 382787 501423 382821
rect 501489 382787 501491 382821
rect 501525 382787 501527 382821
rect 501593 382787 501599 382821
rect 501661 382787 501671 382821
rect 501729 382787 501743 382821
rect 501797 382787 501815 382821
rect 501865 382787 501887 382821
rect 501933 382787 501959 382821
rect 502001 382787 502031 382821
rect 502069 382787 502103 382821
rect 502137 382787 502298 382821
rect 500778 382329 500879 382363
rect 500913 382329 500947 382363
rect 500985 382329 501015 382363
rect 501057 382329 501083 382363
rect 501129 382329 501151 382363
rect 501201 382329 501219 382363
rect 501273 382329 501287 382363
rect 501345 382329 501355 382363
rect 501417 382329 501423 382363
rect 501489 382329 501491 382363
rect 501525 382329 501527 382363
rect 501593 382329 501599 382363
rect 501661 382329 501671 382363
rect 501729 382329 501743 382363
rect 501797 382329 501815 382363
rect 501865 382329 501887 382363
rect 501933 382329 501959 382363
rect 502001 382329 502031 382363
rect 502069 382329 502103 382363
rect 502137 382329 502157 382363
rect 500598 381973 500738 382038
rect 500598 381939 500701 381973
rect 500735 381939 500738 381973
rect 500598 381878 500738 381939
rect 500598 381833 500658 381878
rect 500598 381799 500611 381833
rect 500645 381799 500658 381833
rect 500598 381433 500658 381799
rect 500598 381399 500611 381433
rect 500645 381399 500658 381433
rect 500598 381033 500658 381399
rect 500598 380999 500611 381033
rect 500645 380999 500658 381033
rect 500598 380633 500658 380999
rect 500598 380599 500611 380633
rect 500645 380599 500658 380633
rect 500598 380233 500658 380599
rect 500598 380199 500611 380233
rect 500645 380199 500658 380233
rect 500598 379992 500658 380199
rect 500778 381447 500818 382329
rect 502238 381905 502298 382787
rect 500859 381871 500879 381905
rect 500913 381871 500947 381905
rect 500985 381871 501015 381905
rect 501057 381871 501083 381905
rect 501129 381871 501151 381905
rect 501201 381871 501219 381905
rect 501273 381871 501287 381905
rect 501345 381871 501355 381905
rect 501417 381871 501423 381905
rect 501489 381871 501491 381905
rect 501525 381871 501527 381905
rect 501593 381871 501599 381905
rect 501661 381871 501671 381905
rect 501729 381871 501743 381905
rect 501797 381871 501815 381905
rect 501865 381871 501887 381905
rect 501933 381871 501959 381905
rect 502001 381871 502031 381905
rect 502069 381871 502103 381905
rect 502137 381871 502298 381905
rect 500778 381413 500879 381447
rect 500913 381413 500947 381447
rect 500985 381413 501015 381447
rect 501057 381413 501083 381447
rect 501129 381413 501151 381447
rect 501201 381413 501219 381447
rect 501273 381413 501287 381447
rect 501345 381413 501355 381447
rect 501417 381413 501423 381447
rect 501489 381413 501491 381447
rect 501525 381413 501527 381447
rect 501593 381413 501599 381447
rect 501661 381413 501671 381447
rect 501729 381413 501743 381447
rect 501797 381413 501815 381447
rect 501865 381413 501887 381447
rect 501933 381413 501959 381447
rect 502001 381413 502031 381447
rect 502069 381413 502103 381447
rect 502137 381413 502157 381447
rect 500778 380531 500818 381413
rect 502238 380989 502298 381871
rect 500859 380955 500879 380989
rect 500913 380955 500947 380989
rect 500985 380955 501015 380989
rect 501057 380955 501083 380989
rect 501129 380955 501151 380989
rect 501201 380955 501219 380989
rect 501273 380955 501287 380989
rect 501345 380955 501355 380989
rect 501417 380955 501423 380989
rect 501489 380955 501491 380989
rect 501525 380955 501527 380989
rect 501593 380955 501599 380989
rect 501661 380955 501671 380989
rect 501729 380955 501743 380989
rect 501797 380955 501815 380989
rect 501865 380955 501887 380989
rect 501933 380955 501959 380989
rect 502001 380955 502031 380989
rect 502069 380955 502103 380989
rect 502137 380955 502298 380989
rect 500778 380497 500879 380531
rect 500913 380497 500947 380531
rect 500985 380497 501015 380531
rect 501057 380497 501083 380531
rect 501129 380497 501151 380531
rect 501201 380497 501219 380531
rect 501273 380497 501287 380531
rect 501345 380497 501355 380531
rect 501417 380497 501423 380531
rect 501489 380497 501491 380531
rect 501525 380497 501527 380531
rect 501593 380497 501599 380531
rect 501661 380497 501671 380531
rect 501729 380497 501743 380531
rect 501797 380497 501815 380531
rect 501865 380497 501887 380531
rect 501933 380497 501959 380531
rect 502001 380497 502031 380531
rect 502069 380497 502103 380531
rect 502137 380497 502157 380531
rect 500778 379992 500818 380497
rect 502238 380073 502298 380955
rect 500859 380039 500879 380073
rect 500913 380039 500947 380073
rect 500985 380039 501015 380073
rect 501057 380039 501083 380073
rect 501129 380039 501151 380073
rect 501201 380039 501219 380073
rect 501273 380039 501287 380073
rect 501345 380039 501355 380073
rect 501417 380039 501423 380073
rect 501489 380039 501491 380073
rect 501525 380039 501527 380073
rect 501593 380039 501599 380073
rect 501661 380039 501671 380073
rect 501729 380039 501743 380073
rect 501797 380039 501815 380073
rect 501865 380039 501887 380073
rect 501933 380039 501959 380073
rect 502001 380039 502031 380073
rect 502069 380039 502103 380073
rect 502137 380039 502298 380073
rect 502238 379992 502298 380039
rect 502344 385485 502404 385616
rect 502344 385451 502365 385485
rect 502399 385451 502404 385485
rect 502344 385433 502404 385451
rect 502344 385399 502357 385433
rect 502391 385399 502404 385433
rect 502344 385033 502404 385399
rect 502344 384999 502357 385033
rect 502391 384999 502404 385033
rect 502344 384633 502404 384999
rect 502344 384599 502357 384633
rect 502391 384599 502404 384633
rect 502344 384233 502404 384599
rect 502344 384199 502357 384233
rect 502391 384199 502404 384233
rect 502344 383833 502404 384199
rect 502344 383799 502357 383833
rect 502391 383799 502404 383833
rect 502344 383433 502404 383799
rect 502344 383399 502357 383433
rect 502391 383399 502404 383433
rect 502344 383033 502404 383399
rect 502344 382999 502357 383033
rect 502391 382999 502404 383033
rect 502344 382633 502404 382999
rect 502344 382599 502357 382633
rect 502391 382599 502404 382633
rect 502344 382233 502404 382599
rect 502344 382199 502357 382233
rect 502391 382199 502404 382233
rect 502344 381833 502404 382199
rect 502344 381799 502357 381833
rect 502391 381799 502404 381833
rect 502344 381433 502404 381799
rect 502344 381399 502357 381433
rect 502391 381399 502404 381433
rect 502344 381033 502404 381399
rect 502344 380999 502357 381033
rect 502391 380999 502404 381033
rect 502344 380633 502404 380999
rect 502344 380599 502357 380633
rect 502391 380599 502404 380633
rect 502344 380233 502404 380599
rect 502344 380199 502357 380233
rect 502391 380199 502404 380233
rect 502344 379992 502404 380199
rect 502478 385433 502538 385714
rect 502478 385399 502491 385433
rect 502525 385399 502538 385433
rect 502478 385033 502538 385399
rect 504358 385356 504418 385719
rect 504518 389067 504578 389536
rect 505738 389525 505798 389536
rect 505614 389524 505798 389525
rect 504864 389490 504891 389524
rect 504945 389490 504963 389524
rect 505013 389490 505035 389524
rect 505081 389490 505107 389524
rect 505149 389490 505179 389524
rect 505217 389490 505251 389524
rect 505285 389490 505319 389524
rect 505357 389490 505387 389524
rect 505429 389490 505455 389524
rect 505501 389490 505523 389524
rect 505573 389490 505591 389524
rect 505645 389491 505798 389524
rect 505645 389490 505672 389491
rect 504518 389066 504882 389067
rect 504518 389033 504891 389066
rect 504518 388151 504578 389033
rect 504864 389032 504891 389033
rect 504945 389032 504963 389066
rect 505013 389032 505035 389066
rect 505081 389032 505107 389066
rect 505149 389032 505179 389066
rect 505217 389032 505251 389066
rect 505285 389032 505319 389066
rect 505357 389032 505387 389066
rect 505429 389032 505455 389066
rect 505501 389032 505523 389066
rect 505573 389032 505591 389066
rect 505645 389032 505672 389066
rect 505738 388609 505798 389491
rect 505614 388608 505798 388609
rect 504864 388574 504891 388608
rect 504945 388574 504963 388608
rect 505013 388574 505035 388608
rect 505081 388574 505107 388608
rect 505149 388574 505179 388608
rect 505217 388574 505251 388608
rect 505285 388574 505319 388608
rect 505357 388574 505387 388608
rect 505429 388574 505455 388608
rect 505501 388574 505523 388608
rect 505573 388574 505591 388608
rect 505645 388575 505798 388608
rect 505645 388574 505672 388575
rect 504518 388150 504882 388151
rect 504518 388117 504891 388150
rect 504518 387235 504578 388117
rect 504864 388116 504891 388117
rect 504945 388116 504963 388150
rect 505013 388116 505035 388150
rect 505081 388116 505107 388150
rect 505149 388116 505179 388150
rect 505217 388116 505251 388150
rect 505285 388116 505319 388150
rect 505357 388116 505387 388150
rect 505429 388116 505455 388150
rect 505501 388116 505523 388150
rect 505573 388116 505591 388150
rect 505645 388116 505672 388150
rect 505738 387693 505798 388575
rect 505614 387692 505798 387693
rect 504864 387658 504891 387692
rect 504945 387658 504963 387692
rect 505013 387658 505035 387692
rect 505081 387658 505107 387692
rect 505149 387658 505179 387692
rect 505217 387658 505251 387692
rect 505285 387658 505319 387692
rect 505357 387658 505387 387692
rect 505429 387658 505455 387692
rect 505501 387658 505523 387692
rect 505573 387658 505591 387692
rect 505645 387659 505798 387692
rect 505645 387658 505672 387659
rect 504518 387234 504882 387235
rect 504518 387201 504891 387234
rect 504518 386319 504578 387201
rect 504864 387200 504891 387201
rect 504945 387200 504963 387234
rect 505013 387200 505035 387234
rect 505081 387200 505107 387234
rect 505149 387200 505179 387234
rect 505217 387200 505251 387234
rect 505285 387200 505319 387234
rect 505357 387200 505387 387234
rect 505429 387200 505455 387234
rect 505501 387200 505523 387234
rect 505573 387200 505591 387234
rect 505645 387200 505672 387234
rect 505738 386777 505798 387659
rect 505904 389353 505964 389456
rect 505904 389319 505917 389353
rect 505951 389319 505964 389353
rect 505904 388953 505964 389319
rect 505904 388919 505917 388953
rect 505951 388919 505964 388953
rect 505904 388553 505964 388919
rect 506238 389353 506298 389546
rect 506238 389319 506251 389353
rect 506285 389319 506298 389353
rect 506238 388953 506298 389319
rect 506238 388919 506251 388953
rect 506285 388919 506298 388953
rect 506238 388556 506298 388919
rect 515638 389353 515698 389634
rect 517518 389606 517578 389634
rect 517308 389593 517578 389606
rect 517308 389559 517391 389593
rect 517425 389559 517578 389593
rect 517308 389546 517578 389559
rect 515638 389319 515651 389353
rect 515685 389319 515698 389353
rect 515638 388953 515698 389319
rect 515638 388919 515651 388953
rect 515685 388919 515698 388953
rect 505904 388519 505917 388553
rect 505951 388519 505964 388553
rect 505904 388153 505964 388519
rect 506118 388553 506298 388556
rect 506118 388519 506251 388553
rect 506285 388519 506298 388553
rect 506118 388491 506298 388519
rect 506118 388457 506141 388491
rect 506175 388457 506298 388491
rect 506118 388396 506298 388457
rect 505904 388119 505917 388153
rect 505951 388119 505964 388153
rect 505904 387753 505964 388119
rect 505904 387719 505917 387753
rect 505951 387719 505964 387753
rect 505904 387353 505964 387719
rect 505904 387319 505917 387353
rect 505951 387319 505964 387353
rect 505904 386953 505964 387319
rect 506238 388153 506298 388396
rect 506238 388119 506251 388153
rect 506285 388119 506298 388153
rect 506238 387753 506298 388119
rect 506238 387719 506251 387753
rect 506285 387719 506298 387753
rect 506238 387353 506298 387719
rect 506238 387319 506251 387353
rect 506285 387319 506298 387353
rect 506238 387256 506298 387319
rect 506118 387191 506298 387256
rect 506118 387157 506141 387191
rect 506175 387157 506298 387191
rect 506118 387096 506298 387157
rect 505904 386919 505917 386953
rect 505951 386919 505964 386953
rect 505904 386865 505964 386919
rect 505935 386831 505964 386865
rect 505614 386776 505798 386777
rect 504864 386742 504891 386776
rect 504945 386742 504963 386776
rect 505013 386742 505035 386776
rect 505081 386742 505107 386776
rect 505149 386742 505179 386776
rect 505217 386742 505251 386776
rect 505285 386742 505319 386776
rect 505357 386742 505387 386776
rect 505429 386742 505455 386776
rect 505501 386742 505523 386776
rect 505573 386742 505591 386776
rect 505645 386743 505798 386776
rect 505645 386742 505672 386743
rect 504518 386318 504882 386319
rect 504518 386285 504891 386318
rect 504518 385403 504578 386285
rect 504864 386284 504891 386285
rect 504945 386284 504963 386318
rect 505013 386284 505035 386318
rect 505081 386284 505107 386318
rect 505149 386284 505179 386318
rect 505217 386284 505251 386318
rect 505285 386284 505319 386318
rect 505357 386284 505387 386318
rect 505429 386284 505455 386318
rect 505501 386284 505523 386318
rect 505573 386284 505591 386318
rect 505645 386284 505672 386318
rect 505738 385861 505798 386743
rect 505614 385860 505798 385861
rect 504864 385826 504891 385860
rect 504945 385826 504963 385860
rect 505013 385826 505035 385860
rect 505081 385826 505107 385860
rect 505149 385826 505179 385860
rect 505217 385826 505251 385860
rect 505285 385826 505319 385860
rect 505357 385826 505387 385860
rect 505429 385826 505455 385860
rect 505501 385826 505523 385860
rect 505573 385826 505591 385860
rect 505645 385827 505798 385860
rect 505645 385826 505672 385827
rect 504518 385402 504882 385403
rect 504518 385369 504891 385402
rect 504518 385356 504578 385369
rect 504864 385368 504891 385369
rect 504945 385368 504963 385402
rect 505013 385368 505035 385402
rect 505081 385368 505107 385402
rect 505149 385368 505179 385402
rect 505217 385368 505251 385402
rect 505285 385368 505319 385402
rect 505357 385368 505387 385402
rect 505429 385368 505455 385402
rect 505501 385368 505523 385402
rect 505573 385368 505591 385402
rect 505645 385368 505672 385402
rect 505738 385356 505798 385827
rect 505904 386553 505964 386831
rect 505904 386519 505917 386553
rect 505951 386519 505964 386553
rect 505904 386153 505964 386519
rect 505904 386119 505917 386153
rect 505951 386119 505964 386153
rect 505904 385753 505964 386119
rect 505904 385719 505917 385753
rect 505951 385719 505964 385753
rect 505904 385356 505964 385719
rect 506238 386953 506298 387096
rect 506238 386919 506251 386953
rect 506285 386919 506298 386953
rect 506238 386553 506298 386919
rect 506238 386519 506251 386553
rect 506285 386519 506298 386553
rect 506238 386153 506298 386519
rect 506238 386119 506251 386153
rect 506285 386119 506298 386153
rect 506238 385753 506298 386119
rect 506238 385719 506251 385753
rect 506285 385719 506298 385753
rect 506238 385356 506298 385719
rect 508118 388567 508178 388750
rect 508118 388533 508131 388567
rect 508165 388533 508178 388567
rect 508118 388167 508178 388533
rect 508118 388133 508131 388167
rect 508165 388133 508178 388167
rect 508118 387767 508178 388133
rect 508118 387733 508131 387767
rect 508165 387733 508178 387767
rect 508118 387367 508178 387733
rect 508118 387333 508131 387367
rect 508165 387333 508178 387367
rect 508118 386967 508178 387333
rect 508118 386933 508131 386967
rect 508165 386933 508178 386967
rect 508118 386567 508178 386933
rect 508118 386533 508131 386567
rect 508165 386533 508178 386567
rect 508118 386167 508178 386533
rect 508118 386133 508131 386167
rect 508165 386133 508178 386167
rect 508118 385767 508178 386133
rect 508118 385733 508131 385767
rect 508165 385733 508178 385767
rect 508118 385367 508178 385733
rect 502478 384999 502491 385033
rect 502525 384999 502538 385033
rect 508118 385333 508131 385367
rect 508165 385333 508178 385367
rect 502478 384633 502538 384999
rect 502478 384599 502491 384633
rect 502525 384599 502538 384633
rect 502478 384233 502538 384599
rect 502478 384199 502491 384233
rect 502525 384199 502538 384233
rect 502478 383833 502538 384199
rect 502478 383799 502491 383833
rect 502525 383799 502538 383833
rect 502478 383433 502538 383799
rect 502478 383399 502491 383433
rect 502525 383399 502538 383433
rect 502478 383033 502538 383399
rect 502478 382999 502491 383033
rect 502525 382999 502538 383033
rect 502478 382633 502538 382999
rect 502478 382599 502491 382633
rect 502525 382599 502538 382633
rect 502478 382233 502538 382599
rect 502478 382199 502491 382233
rect 502525 382199 502538 382233
rect 502478 381833 502538 382199
rect 502478 381799 502491 381833
rect 502525 381799 502538 381833
rect 502478 381433 502538 381799
rect 502478 381399 502491 381433
rect 502525 381399 502538 381433
rect 502478 381033 502538 381399
rect 502478 380999 502491 381033
rect 502525 380999 502538 381033
rect 502478 380633 502538 380999
rect 502478 380599 502491 380633
rect 502525 380599 502538 380633
rect 502478 380233 502538 380599
rect 502478 380199 502491 380233
rect 502525 380199 502538 380233
rect 502478 379992 502538 380199
rect 504358 384843 504418 385026
rect 504358 384809 504371 384843
rect 504405 384809 504418 384843
rect 504358 384443 504418 384809
rect 504358 384409 504371 384443
rect 504405 384409 504418 384443
rect 504358 384043 504418 384409
rect 504358 384009 504371 384043
rect 504405 384009 504418 384043
rect 504358 383643 504418 384009
rect 504358 383609 504371 383643
rect 504405 383609 504418 383643
rect 504358 383243 504418 383609
rect 504358 383209 504371 383243
rect 504405 383209 504418 383243
rect 504358 382843 504418 383209
rect 504358 382809 504371 382843
rect 504405 382809 504418 382843
rect 504358 382443 504418 382809
rect 504358 382409 504371 382443
rect 504405 382409 504418 382443
rect 504358 382043 504418 382409
rect 504358 382009 504371 382043
rect 504405 382009 504418 382043
rect 504358 381643 504418 382009
rect 504358 381609 504371 381643
rect 504405 381609 504418 381643
rect 504358 381243 504418 381609
rect 504358 381209 504371 381243
rect 504405 381209 504418 381243
rect 504358 380843 504418 381209
rect 504358 380809 504371 380843
rect 504405 380809 504418 380843
rect 504358 380443 504418 380809
rect 504358 380409 504371 380443
rect 504405 380409 504418 380443
rect 504358 380043 504418 380409
rect 504358 380009 504371 380043
rect 504405 380009 504418 380043
rect 498718 379707 498731 379741
rect 498765 379707 498778 379741
rect 498718 379341 498778 379707
rect 498718 379307 498731 379341
rect 498765 379307 498778 379341
rect 498718 378941 498778 379307
rect 498718 378907 498731 378941
rect 498765 378907 498778 378941
rect 498718 378541 498778 378907
rect 498718 378507 498731 378541
rect 498765 378507 498778 378541
rect 498718 378141 498778 378507
rect 498718 378107 498731 378141
rect 498765 378107 498778 378141
rect 498718 377741 498778 378107
rect 504358 379643 504418 380009
rect 504358 379609 504371 379643
rect 504405 379609 504418 379643
rect 504358 379243 504418 379609
rect 504358 379209 504371 379243
rect 504405 379209 504418 379243
rect 504358 378843 504418 379209
rect 504358 378809 504371 378843
rect 504405 378809 504418 378843
rect 504358 378443 504418 378809
rect 504358 378409 504371 378443
rect 504405 378409 504418 378443
rect 504358 378043 504418 378409
rect 504358 378009 504371 378043
rect 504405 378009 504418 378043
rect 504358 377858 504418 378009
rect 506238 384843 506298 385026
rect 506238 384809 506251 384843
rect 506285 384809 506298 384843
rect 506238 384443 506298 384809
rect 506238 384409 506251 384443
rect 506285 384409 506298 384443
rect 506238 384043 506298 384409
rect 506238 384009 506251 384043
rect 506285 384009 506298 384043
rect 506238 383643 506298 384009
rect 506238 383609 506251 383643
rect 506285 383609 506298 383643
rect 506238 383243 506298 383609
rect 506238 383209 506251 383243
rect 506285 383209 506298 383243
rect 506238 382843 506298 383209
rect 506238 382809 506251 382843
rect 506285 382809 506298 382843
rect 506238 382443 506298 382809
rect 506238 382409 506251 382443
rect 506285 382409 506298 382443
rect 506238 382043 506298 382409
rect 506238 382009 506251 382043
rect 506285 382009 506298 382043
rect 506238 381643 506298 382009
rect 506238 381609 506251 381643
rect 506285 381609 506298 381643
rect 506238 381243 506298 381609
rect 508118 384967 508178 385333
rect 508118 384933 508131 384967
rect 508165 384933 508178 384967
rect 508118 384567 508178 384933
rect 508118 384533 508131 384567
rect 508165 384533 508178 384567
rect 508118 384167 508178 384533
rect 508118 384133 508131 384167
rect 508165 384133 508178 384167
rect 508118 383767 508178 384133
rect 508118 383733 508131 383767
rect 508165 383733 508178 383767
rect 508118 383367 508178 383733
rect 508118 383333 508131 383367
rect 508165 383333 508178 383367
rect 508118 382967 508178 383333
rect 508118 382933 508131 382967
rect 508165 382933 508178 382967
rect 508118 382567 508178 382933
rect 508118 382533 508131 382567
rect 508165 382533 508178 382567
rect 508118 382167 508178 382533
rect 508118 382133 508131 382167
rect 508165 382133 508178 382167
rect 508118 381767 508178 382133
rect 508118 381733 508131 381767
rect 508165 381733 508178 381767
rect 508118 381582 508178 381733
rect 509998 388567 510058 388750
rect 509998 388533 510011 388567
rect 510045 388533 510058 388567
rect 509998 388167 510058 388533
rect 509998 388133 510011 388167
rect 510045 388133 510058 388167
rect 509998 387767 510058 388133
rect 509998 387733 510011 387767
rect 510045 387733 510058 387767
rect 515638 388553 515698 388919
rect 515638 388519 515651 388553
rect 515685 388519 515698 388553
rect 515638 388153 515698 388519
rect 515638 388119 515651 388153
rect 515685 388119 515698 388153
rect 515638 387753 515698 388119
rect 509998 387367 510058 387733
rect 509998 387333 510011 387367
rect 510045 387333 510058 387367
rect 509998 386967 510058 387333
rect 509998 386933 510011 386967
rect 510045 386933 510058 386967
rect 509998 386567 510058 386933
rect 509998 386533 510011 386567
rect 510045 386533 510058 386567
rect 509998 386167 510058 386533
rect 509998 386133 510011 386167
rect 510045 386133 510058 386167
rect 509998 385767 510058 386133
rect 509998 385733 510011 385767
rect 510045 385733 510058 385767
rect 509998 385367 510058 385733
rect 509998 385333 510011 385367
rect 510045 385333 510058 385367
rect 509998 384967 510058 385333
rect 511878 387569 511938 387752
rect 511878 387535 511891 387569
rect 511925 387535 511938 387569
rect 511878 387369 511938 387535
rect 511878 387335 511891 387369
rect 511925 387335 511938 387369
rect 511878 387169 511938 387335
rect 513758 387569 513818 387752
rect 513758 387535 513771 387569
rect 513805 387535 513818 387569
rect 513758 387369 513818 387535
rect 513758 387335 513771 387369
rect 513805 387335 513818 387369
rect 511878 387135 511891 387169
rect 511925 387135 511938 387169
rect 511878 386969 511938 387135
rect 511878 386935 511891 386969
rect 511925 386935 511938 386969
rect 511878 386769 511938 386935
rect 513758 387169 513818 387335
rect 513758 387135 513771 387169
rect 513805 387135 513818 387169
rect 513758 386969 513818 387135
rect 513758 386935 513771 386969
rect 513805 386935 513818 386969
rect 513758 386840 513818 386935
rect 511878 386735 511891 386769
rect 511925 386735 511938 386769
rect 511878 386569 511938 386735
rect 511878 386535 511891 386569
rect 511925 386535 511938 386569
rect 511878 386369 511938 386535
rect 511878 386335 511891 386369
rect 511925 386335 511938 386369
rect 511878 386169 511938 386335
rect 512818 386769 513818 386840
rect 512818 386753 513771 386769
rect 512818 386311 512857 386753
rect 512959 386735 513771 386753
rect 513805 386735 513818 386769
rect 512959 386569 513818 386735
rect 512959 386535 513771 386569
rect 513805 386535 513818 386569
rect 512959 386369 513818 386535
rect 512959 386335 513771 386369
rect 513805 386335 513818 386369
rect 512959 386311 513818 386335
rect 512818 386224 513818 386311
rect 511878 386135 511891 386169
rect 511925 386135 511938 386169
rect 511878 385969 511938 386135
rect 511878 385935 511891 385969
rect 511925 385935 511938 385969
rect 511878 385769 511938 385935
rect 511878 385735 511891 385769
rect 511925 385735 511938 385769
rect 513758 386169 513818 386224
rect 513758 386135 513771 386169
rect 513805 386135 513818 386169
rect 513758 385969 513818 386135
rect 513758 385935 513771 385969
rect 513805 385935 513818 385969
rect 513758 385769 513818 385935
rect 511878 385569 511938 385735
rect 511878 385535 511891 385569
rect 511925 385535 511938 385569
rect 511878 385312 511938 385535
rect 512713 385312 513103 385744
rect 513758 385735 513771 385769
rect 513805 385735 513818 385769
rect 513758 385569 513818 385735
rect 513758 385535 513771 385569
rect 513805 385535 513818 385569
rect 513758 385312 513818 385535
rect 515638 387719 515651 387753
rect 515685 387719 515698 387753
rect 515638 387353 515698 387719
rect 515638 387319 515651 387353
rect 515685 387319 515698 387353
rect 515638 386953 515698 387319
rect 515638 386919 515651 386953
rect 515685 386919 515698 386953
rect 515638 386553 515698 386919
rect 515638 386519 515651 386553
rect 515685 386519 515698 386553
rect 515638 386153 515698 386519
rect 515638 386119 515651 386153
rect 515685 386119 515698 386153
rect 515638 385753 515698 386119
rect 515638 385719 515651 385753
rect 515685 385719 515698 385753
rect 515638 385356 515698 385719
rect 515798 389067 515858 389536
rect 517018 389525 517078 389536
rect 516894 389524 517078 389525
rect 516144 389490 516171 389524
rect 516225 389490 516243 389524
rect 516293 389490 516315 389524
rect 516361 389490 516387 389524
rect 516429 389490 516459 389524
rect 516497 389490 516531 389524
rect 516565 389490 516599 389524
rect 516637 389490 516667 389524
rect 516709 389490 516735 389524
rect 516781 389490 516803 389524
rect 516853 389490 516871 389524
rect 516925 389491 517078 389524
rect 516925 389490 516952 389491
rect 515798 389066 516162 389067
rect 515798 389033 516171 389066
rect 515798 388151 515858 389033
rect 516144 389032 516171 389033
rect 516225 389032 516243 389066
rect 516293 389032 516315 389066
rect 516361 389032 516387 389066
rect 516429 389032 516459 389066
rect 516497 389032 516531 389066
rect 516565 389032 516599 389066
rect 516637 389032 516667 389066
rect 516709 389032 516735 389066
rect 516781 389032 516803 389066
rect 516853 389032 516871 389066
rect 516925 389032 516952 389066
rect 517018 388609 517078 389491
rect 516894 388608 517078 388609
rect 516144 388574 516171 388608
rect 516225 388574 516243 388608
rect 516293 388574 516315 388608
rect 516361 388574 516387 388608
rect 516429 388574 516459 388608
rect 516497 388574 516531 388608
rect 516565 388574 516599 388608
rect 516637 388574 516667 388608
rect 516709 388574 516735 388608
rect 516781 388574 516803 388608
rect 516853 388574 516871 388608
rect 516925 388575 517078 388608
rect 516925 388574 516952 388575
rect 515798 388150 516162 388151
rect 515798 388117 516171 388150
rect 515798 387235 515858 388117
rect 516144 388116 516171 388117
rect 516225 388116 516243 388150
rect 516293 388116 516315 388150
rect 516361 388116 516387 388150
rect 516429 388116 516459 388150
rect 516497 388116 516531 388150
rect 516565 388116 516599 388150
rect 516637 388116 516667 388150
rect 516709 388116 516735 388150
rect 516781 388116 516803 388150
rect 516853 388116 516871 388150
rect 516925 388116 516952 388150
rect 517018 387693 517078 388575
rect 516894 387692 517078 387693
rect 516144 387658 516171 387692
rect 516225 387658 516243 387692
rect 516293 387658 516315 387692
rect 516361 387658 516387 387692
rect 516429 387658 516459 387692
rect 516497 387658 516531 387692
rect 516565 387658 516599 387692
rect 516637 387658 516667 387692
rect 516709 387658 516735 387692
rect 516781 387658 516803 387692
rect 516853 387658 516871 387692
rect 516925 387659 517078 387692
rect 516925 387658 516952 387659
rect 515798 387234 516162 387235
rect 515798 387201 516171 387234
rect 515798 386319 515858 387201
rect 516144 387200 516171 387201
rect 516225 387200 516243 387234
rect 516293 387200 516315 387234
rect 516361 387200 516387 387234
rect 516429 387200 516459 387234
rect 516497 387200 516531 387234
rect 516565 387200 516599 387234
rect 516637 387200 516667 387234
rect 516709 387200 516735 387234
rect 516781 387200 516803 387234
rect 516853 387200 516871 387234
rect 516925 387200 516952 387234
rect 517018 386777 517078 387659
rect 516894 386776 517078 386777
rect 516144 386742 516171 386776
rect 516225 386742 516243 386776
rect 516293 386742 516315 386776
rect 516361 386742 516387 386776
rect 516429 386742 516459 386776
rect 516497 386742 516531 386776
rect 516565 386742 516599 386776
rect 516637 386742 516667 386776
rect 516709 386742 516735 386776
rect 516781 386742 516803 386776
rect 516853 386742 516871 386776
rect 516925 386743 517078 386776
rect 516925 386742 516952 386743
rect 515798 386318 516162 386319
rect 515798 386285 516171 386318
rect 515798 385403 515858 386285
rect 516144 386284 516171 386285
rect 516225 386284 516243 386318
rect 516293 386284 516315 386318
rect 516361 386284 516387 386318
rect 516429 386284 516459 386318
rect 516497 386284 516531 386318
rect 516565 386284 516599 386318
rect 516637 386284 516667 386318
rect 516709 386284 516735 386318
rect 516781 386284 516803 386318
rect 516853 386284 516871 386318
rect 516925 386284 516952 386318
rect 517018 385861 517078 386743
rect 516894 385860 517078 385861
rect 516144 385826 516171 385860
rect 516225 385826 516243 385860
rect 516293 385826 516315 385860
rect 516361 385826 516387 385860
rect 516429 385826 516459 385860
rect 516497 385826 516531 385860
rect 516565 385826 516599 385860
rect 516637 385826 516667 385860
rect 516709 385826 516735 385860
rect 516781 385826 516803 385860
rect 516853 385826 516871 385860
rect 516925 385827 517078 385860
rect 516925 385826 516952 385827
rect 515798 385402 516162 385403
rect 515798 385369 516171 385402
rect 515798 385356 515858 385369
rect 516144 385368 516171 385369
rect 516225 385368 516243 385402
rect 516293 385368 516315 385402
rect 516361 385368 516387 385402
rect 516429 385368 516459 385402
rect 516497 385368 516531 385402
rect 516565 385368 516599 385402
rect 516637 385368 516667 385402
rect 516709 385368 516735 385402
rect 516781 385368 516803 385402
rect 516853 385368 516871 385402
rect 516925 385368 516952 385402
rect 517018 385356 517078 385827
rect 517184 389353 517244 389456
rect 517184 389319 517197 389353
rect 517231 389319 517244 389353
rect 517184 388953 517244 389319
rect 517184 388919 517197 388953
rect 517231 388919 517244 388953
rect 517184 388553 517244 388919
rect 517518 389353 517578 389546
rect 517518 389319 517531 389353
rect 517565 389319 517578 389353
rect 517518 388953 517578 389319
rect 517518 388919 517531 388953
rect 517565 388919 517578 388953
rect 517518 388556 517578 388919
rect 519398 389501 519458 389667
rect 520338 390101 521338 390172
rect 520338 390085 521291 390101
rect 520338 389643 520377 390085
rect 520479 390067 521291 390085
rect 521325 390067 521338 390101
rect 520479 389901 521338 390067
rect 520479 389867 521291 389901
rect 521325 389867 521338 389901
rect 520479 389701 521338 389867
rect 520479 389667 521291 389701
rect 521325 389667 521338 389701
rect 520479 389643 521338 389667
rect 520338 389556 521338 389643
rect 519398 389467 519411 389501
rect 519445 389467 519458 389501
rect 519398 389301 519458 389467
rect 519398 389267 519411 389301
rect 519445 389267 519458 389301
rect 519398 389101 519458 389267
rect 519398 389067 519411 389101
rect 519445 389067 519458 389101
rect 521278 389501 521338 389556
rect 521278 389467 521291 389501
rect 521325 389467 521338 389501
rect 521278 389301 521338 389467
rect 521278 389267 521291 389301
rect 521325 389267 521338 389301
rect 521278 389101 521338 389267
rect 519398 388901 519458 389067
rect 519398 388867 519411 388901
rect 519445 388867 519458 388901
rect 519398 388644 519458 388867
rect 520233 388644 520623 389076
rect 521278 389067 521291 389101
rect 521325 389067 521338 389101
rect 521278 388901 521338 389067
rect 521278 388867 521291 388901
rect 521325 388867 521338 388901
rect 521278 388644 521338 388867
rect 523158 390194 523218 390222
rect 523158 390181 523428 390194
rect 523158 390147 523311 390181
rect 523345 390147 523428 390181
rect 523158 390134 523428 390147
rect 523158 389941 523218 390134
rect 524798 390077 524858 390124
rect 523158 389907 523171 389941
rect 523205 389907 523218 389941
rect 523158 389541 523218 389907
rect 523158 389507 523171 389541
rect 523205 389507 523218 389541
rect 523158 389146 523218 389507
rect 523338 389619 523378 390064
rect 523419 390043 523439 390077
rect 523473 390043 523507 390077
rect 523545 390043 523575 390077
rect 523617 390043 523643 390077
rect 523689 390043 523711 390077
rect 523761 390043 523779 390077
rect 523833 390043 523847 390077
rect 523905 390043 523915 390077
rect 523977 390043 523983 390077
rect 524049 390043 524051 390077
rect 524085 390043 524087 390077
rect 524153 390043 524159 390077
rect 524221 390043 524231 390077
rect 524289 390043 524303 390077
rect 524357 390043 524375 390077
rect 524425 390043 524447 390077
rect 524493 390043 524519 390077
rect 524561 390043 524591 390077
rect 524629 390043 524663 390077
rect 524697 390043 524858 390077
rect 523338 389585 523439 389619
rect 523473 389585 523507 389619
rect 523545 389585 523575 389619
rect 523617 389585 523643 389619
rect 523689 389585 523711 389619
rect 523761 389585 523779 389619
rect 523833 389585 523847 389619
rect 523905 389585 523915 389619
rect 523977 389585 523983 389619
rect 524049 389585 524051 389619
rect 524085 389585 524087 389619
rect 524153 389585 524159 389619
rect 524221 389585 524231 389619
rect 524289 389585 524303 389619
rect 524357 389585 524375 389619
rect 524425 389585 524447 389619
rect 524493 389585 524519 389619
rect 524561 389585 524591 389619
rect 524629 389585 524663 389619
rect 524697 389585 524717 389619
rect 523158 389141 523298 389146
rect 523158 389107 523171 389141
rect 523205 389107 523298 389141
rect 523158 389081 523298 389107
rect 523158 389047 523261 389081
rect 523295 389047 523298 389081
rect 523158 388986 523298 389047
rect 523158 388741 523218 388986
rect 523158 388707 523171 388741
rect 523205 388707 523218 388741
rect 517184 388519 517197 388553
rect 517231 388519 517244 388553
rect 517184 388153 517244 388519
rect 517398 388553 517578 388556
rect 517398 388519 517531 388553
rect 517565 388519 517578 388553
rect 517398 388491 517578 388519
rect 517398 388457 517421 388491
rect 517455 388457 517578 388491
rect 517398 388396 517578 388457
rect 517184 388119 517197 388153
rect 517231 388119 517244 388153
rect 517184 387753 517244 388119
rect 517184 387719 517197 387753
rect 517231 387719 517244 387753
rect 517184 387417 517244 387719
rect 517184 387383 517189 387417
rect 517223 387383 517244 387417
rect 517184 387353 517244 387383
rect 517184 387319 517197 387353
rect 517231 387319 517244 387353
rect 517184 386953 517244 387319
rect 517518 388153 517578 388396
rect 517518 388119 517531 388153
rect 517565 388119 517578 388153
rect 517518 387753 517578 388119
rect 517518 387719 517531 387753
rect 517565 387719 517578 387753
rect 523158 388341 523218 388707
rect 523158 388307 523171 388341
rect 523205 388307 523218 388341
rect 523158 387941 523218 388307
rect 523158 387907 523171 387941
rect 523205 387907 523218 387941
rect 523158 387846 523218 387907
rect 523338 388703 523378 389585
rect 524798 389161 524858 390043
rect 523419 389127 523439 389161
rect 523473 389127 523507 389161
rect 523545 389127 523575 389161
rect 523617 389127 523643 389161
rect 523689 389127 523711 389161
rect 523761 389127 523779 389161
rect 523833 389127 523847 389161
rect 523905 389127 523915 389161
rect 523977 389127 523983 389161
rect 524049 389127 524051 389161
rect 524085 389127 524087 389161
rect 524153 389127 524159 389161
rect 524221 389127 524231 389161
rect 524289 389127 524303 389161
rect 524357 389127 524375 389161
rect 524425 389127 524447 389161
rect 524493 389127 524519 389161
rect 524561 389127 524591 389161
rect 524629 389127 524663 389161
rect 524697 389127 524858 389161
rect 523338 388669 523439 388703
rect 523473 388669 523507 388703
rect 523545 388669 523575 388703
rect 523617 388669 523643 388703
rect 523689 388669 523711 388703
rect 523761 388669 523779 388703
rect 523833 388669 523847 388703
rect 523905 388669 523915 388703
rect 523977 388669 523983 388703
rect 524049 388669 524051 388703
rect 524085 388669 524087 388703
rect 524153 388669 524159 388703
rect 524221 388669 524231 388703
rect 524289 388669 524303 388703
rect 524357 388669 524375 388703
rect 524425 388669 524447 388703
rect 524493 388669 524519 388703
rect 524561 388669 524591 388703
rect 524629 388669 524663 388703
rect 524697 388669 524717 388703
rect 523158 387781 523298 387846
rect 517518 387353 517578 387719
rect 517518 387319 517531 387353
rect 517565 387319 517578 387353
rect 517518 387256 517578 387319
rect 517398 387191 517578 387256
rect 517398 387157 517421 387191
rect 517455 387157 517578 387191
rect 517398 387096 517578 387157
rect 517184 386919 517197 386953
rect 517231 386919 517244 386953
rect 517184 386553 517244 386919
rect 517184 386519 517197 386553
rect 517231 386519 517244 386553
rect 517184 386153 517244 386519
rect 517184 386119 517197 386153
rect 517231 386119 517244 386153
rect 517184 385753 517244 386119
rect 517184 385719 517197 385753
rect 517231 385719 517244 385753
rect 517184 385356 517244 385719
rect 517518 386953 517578 387096
rect 517518 386919 517531 386953
rect 517565 386919 517578 386953
rect 517518 386553 517578 386919
rect 517518 386519 517531 386553
rect 517565 386519 517578 386553
rect 517518 386153 517578 386519
rect 517518 386119 517531 386153
rect 517565 386119 517578 386153
rect 517518 385753 517578 386119
rect 517518 385719 517531 385753
rect 517565 385719 517578 385753
rect 517518 385356 517578 385719
rect 519398 387569 519458 387752
rect 519398 387535 519411 387569
rect 519445 387535 519458 387569
rect 519398 387369 519458 387535
rect 519398 387335 519411 387369
rect 519445 387335 519458 387369
rect 519398 387169 519458 387335
rect 521278 387569 521338 387752
rect 521278 387535 521291 387569
rect 521325 387535 521338 387569
rect 521278 387369 521338 387535
rect 521278 387335 521291 387369
rect 521325 387335 521338 387369
rect 519398 387135 519411 387169
rect 519445 387135 519458 387169
rect 519398 386969 519458 387135
rect 519398 386935 519411 386969
rect 519445 386935 519458 386969
rect 519398 386769 519458 386935
rect 521278 387169 521338 387335
rect 521278 387135 521291 387169
rect 521325 387135 521338 387169
rect 521278 386969 521338 387135
rect 521278 386935 521291 386969
rect 521325 386935 521338 386969
rect 521278 386840 521338 386935
rect 519398 386735 519411 386769
rect 519445 386735 519458 386769
rect 519398 386569 519458 386735
rect 519398 386535 519411 386569
rect 519445 386535 519458 386569
rect 519398 386369 519458 386535
rect 519398 386335 519411 386369
rect 519445 386335 519458 386369
rect 519398 386169 519458 386335
rect 520338 386769 521338 386840
rect 520338 386753 521291 386769
rect 520338 386311 520377 386753
rect 520479 386735 521291 386753
rect 521325 386735 521338 386769
rect 520479 386569 521338 386735
rect 520479 386535 521291 386569
rect 521325 386535 521338 386569
rect 520479 386369 521338 386535
rect 520479 386335 521291 386369
rect 521325 386335 521338 386369
rect 520479 386311 521338 386335
rect 520338 386224 521338 386311
rect 519398 386135 519411 386169
rect 519445 386135 519458 386169
rect 519398 385969 519458 386135
rect 519398 385935 519411 385969
rect 519445 385935 519458 385969
rect 519398 385769 519458 385935
rect 519398 385735 519411 385769
rect 519445 385735 519458 385769
rect 521278 386169 521338 386224
rect 521278 386135 521291 386169
rect 521325 386135 521338 386169
rect 521278 385969 521338 386135
rect 521278 385935 521291 385969
rect 521325 385935 521338 385969
rect 521278 385769 521338 385935
rect 519398 385569 519458 385735
rect 519398 385535 519411 385569
rect 519445 385535 519458 385569
rect 519398 385312 519458 385535
rect 520233 385312 520623 385744
rect 521278 385735 521291 385769
rect 521325 385735 521338 385769
rect 521278 385569 521338 385735
rect 521278 385535 521291 385569
rect 521325 385535 521338 385569
rect 521278 385312 521338 385535
rect 523158 387747 523261 387781
rect 523295 387747 523298 387781
rect 523158 387686 523298 387747
rect 523338 387787 523378 388669
rect 524798 388245 524858 389127
rect 523419 388211 523439 388245
rect 523473 388211 523507 388245
rect 523545 388211 523575 388245
rect 523617 388211 523643 388245
rect 523689 388211 523711 388245
rect 523761 388211 523779 388245
rect 523833 388211 523847 388245
rect 523905 388211 523915 388245
rect 523977 388211 523983 388245
rect 524049 388211 524051 388245
rect 524085 388211 524087 388245
rect 524153 388211 524159 388245
rect 524221 388211 524231 388245
rect 524289 388211 524303 388245
rect 524357 388211 524375 388245
rect 524425 388211 524447 388245
rect 524493 388211 524519 388245
rect 524561 388211 524591 388245
rect 524629 388211 524663 388245
rect 524697 388211 524858 388245
rect 523338 387753 523439 387787
rect 523473 387753 523507 387787
rect 523545 387753 523575 387787
rect 523617 387753 523643 387787
rect 523689 387753 523711 387787
rect 523761 387753 523779 387787
rect 523833 387753 523847 387787
rect 523905 387753 523915 387787
rect 523977 387753 523983 387787
rect 524049 387753 524051 387787
rect 524085 387753 524087 387787
rect 524153 387753 524159 387787
rect 524221 387753 524231 387787
rect 524289 387753 524303 387787
rect 524357 387753 524375 387787
rect 524425 387753 524447 387787
rect 524493 387753 524519 387787
rect 524561 387753 524591 387787
rect 524629 387753 524663 387787
rect 524697 387753 524717 387787
rect 523158 387541 523218 387686
rect 523158 387507 523171 387541
rect 523205 387507 523218 387541
rect 523158 387141 523218 387507
rect 523158 387107 523171 387141
rect 523205 387107 523218 387141
rect 523158 386741 523218 387107
rect 523158 386707 523171 386741
rect 523205 386707 523218 386741
rect 523158 386546 523218 386707
rect 523338 386871 523378 387753
rect 524798 387329 524858 388211
rect 523419 387295 523439 387329
rect 523473 387295 523507 387329
rect 523545 387295 523575 387329
rect 523617 387295 523643 387329
rect 523689 387295 523711 387329
rect 523761 387295 523779 387329
rect 523833 387295 523847 387329
rect 523905 387295 523915 387329
rect 523977 387295 523983 387329
rect 524049 387295 524051 387329
rect 524085 387295 524087 387329
rect 524153 387295 524159 387329
rect 524221 387295 524231 387329
rect 524289 387295 524303 387329
rect 524357 387295 524375 387329
rect 524425 387295 524447 387329
rect 524493 387295 524519 387329
rect 524561 387295 524591 387329
rect 524629 387295 524663 387329
rect 524697 387295 524858 387329
rect 523338 386837 523439 386871
rect 523473 386837 523507 386871
rect 523545 386837 523575 386871
rect 523617 386837 523643 386871
rect 523689 386837 523711 386871
rect 523761 386837 523779 386871
rect 523833 386837 523847 386871
rect 523905 386837 523915 386871
rect 523977 386837 523983 386871
rect 524049 386837 524051 386871
rect 524085 386837 524087 386871
rect 524153 386837 524159 386871
rect 524221 386837 524231 386871
rect 524289 386837 524303 386871
rect 524357 386837 524375 386871
rect 524425 386837 524447 386871
rect 524493 386837 524519 386871
rect 524561 386837 524591 386871
rect 524629 386837 524663 386871
rect 524697 386837 524717 386871
rect 523158 386481 523298 386546
rect 523158 386447 523261 386481
rect 523295 386447 523298 386481
rect 523158 386386 523298 386447
rect 523158 386341 523218 386386
rect 523158 386307 523171 386341
rect 523205 386307 523218 386341
rect 523158 385941 523218 386307
rect 523158 385907 523171 385941
rect 523205 385907 523218 385941
rect 523158 385541 523218 385907
rect 523158 385507 523171 385541
rect 523205 385507 523218 385541
rect 523158 385246 523218 385507
rect 523338 385955 523378 386837
rect 524798 386413 524858 387295
rect 523419 386379 523439 386413
rect 523473 386379 523507 386413
rect 523545 386379 523575 386413
rect 523617 386379 523643 386413
rect 523689 386379 523711 386413
rect 523761 386379 523779 386413
rect 523833 386379 523847 386413
rect 523905 386379 523915 386413
rect 523977 386379 523983 386413
rect 524049 386379 524051 386413
rect 524085 386379 524087 386413
rect 524153 386379 524159 386413
rect 524221 386379 524231 386413
rect 524289 386379 524303 386413
rect 524357 386379 524375 386413
rect 524425 386379 524447 386413
rect 524493 386379 524519 386413
rect 524561 386379 524591 386413
rect 524629 386379 524663 386413
rect 524697 386379 524858 386413
rect 523338 385921 523439 385955
rect 523473 385921 523507 385955
rect 523545 385921 523575 385955
rect 523617 385921 523643 385955
rect 523689 385921 523711 385955
rect 523761 385921 523779 385955
rect 523833 385921 523847 385955
rect 523905 385921 523915 385955
rect 523977 385921 523983 385955
rect 524049 385921 524051 385955
rect 524085 385921 524087 385955
rect 524153 385921 524159 385955
rect 524221 385921 524231 385955
rect 524289 385921 524303 385955
rect 524357 385921 524375 385955
rect 524425 385921 524447 385955
rect 524493 385921 524519 385955
rect 524561 385921 524591 385955
rect 524629 385921 524663 385955
rect 524697 385921 524717 385955
rect 523158 385181 523298 385246
rect 523158 385147 523261 385181
rect 523295 385147 523298 385181
rect 523158 385141 523298 385147
rect 523158 385107 523171 385141
rect 523205 385107 523298 385141
rect 523158 385086 523298 385107
rect 509998 384933 510011 384967
rect 510045 384933 510058 384967
rect 509998 384567 510058 384933
rect 509998 384533 510011 384567
rect 510045 384533 510058 384567
rect 509998 384167 510058 384533
rect 509998 384133 510011 384167
rect 510045 384133 510058 384167
rect 509998 383767 510058 384133
rect 509998 383733 510011 383767
rect 510045 383733 510058 383767
rect 509998 383367 510058 383733
rect 509998 383333 510011 383367
rect 510045 383333 510058 383367
rect 509998 382967 510058 383333
rect 509998 382933 510011 382967
rect 510045 382933 510058 382967
rect 509998 382567 510058 382933
rect 509998 382533 510011 382567
rect 510045 382533 510058 382567
rect 509998 382167 510058 382533
rect 509998 382133 510011 382167
rect 510045 382133 510058 382167
rect 509998 381767 510058 382133
rect 509998 381733 510011 381767
rect 510045 381733 510058 381767
rect 509998 381582 510058 381733
rect 511878 384843 511938 385026
rect 511878 384809 511891 384843
rect 511925 384809 511938 384843
rect 511878 384443 511938 384809
rect 511878 384409 511891 384443
rect 511925 384409 511938 384443
rect 511878 384043 511938 384409
rect 511878 384009 511891 384043
rect 511925 384009 511938 384043
rect 511878 383643 511938 384009
rect 511878 383609 511891 383643
rect 511925 383609 511938 383643
rect 511878 383243 511938 383609
rect 511878 383209 511891 383243
rect 511925 383209 511938 383243
rect 511878 382843 511938 383209
rect 511878 382809 511891 382843
rect 511925 382809 511938 382843
rect 511878 382443 511938 382809
rect 511878 382409 511891 382443
rect 511925 382409 511938 382443
rect 511878 382043 511938 382409
rect 511878 382009 511891 382043
rect 511925 382009 511938 382043
rect 511878 381643 511938 382009
rect 511878 381609 511891 381643
rect 511925 381609 511938 381643
rect 506238 381209 506251 381243
rect 506285 381209 506298 381243
rect 506238 380843 506298 381209
rect 506238 380809 506251 380843
rect 506285 380809 506298 380843
rect 506238 380443 506298 380809
rect 506238 380409 506251 380443
rect 506285 380409 506298 380443
rect 506238 380043 506298 380409
rect 506238 380009 506251 380043
rect 506285 380009 506298 380043
rect 506238 379643 506298 380009
rect 506238 379609 506251 379643
rect 506285 379609 506298 379643
rect 506238 379243 506298 379609
rect 506238 379209 506251 379243
rect 506285 379209 506298 379243
rect 506238 378843 506298 379209
rect 506238 378809 506251 378843
rect 506285 378809 506298 378843
rect 506238 378443 506298 378809
rect 506238 378409 506251 378443
rect 506285 378409 506298 378443
rect 506238 378043 506298 378409
rect 506238 378009 506251 378043
rect 506285 378009 506298 378043
rect 506238 377858 506298 378009
rect 508118 381119 508178 381302
rect 508118 381085 508131 381119
rect 508165 381085 508178 381119
rect 508118 380719 508178 381085
rect 508118 380685 508131 380719
rect 508165 380685 508178 380719
rect 508118 380319 508178 380685
rect 508118 380285 508131 380319
rect 508165 380285 508178 380319
rect 508118 379919 508178 380285
rect 508118 379885 508131 379919
rect 508165 379885 508178 379919
rect 508118 379519 508178 379885
rect 508118 379485 508131 379519
rect 508165 379485 508178 379519
rect 508118 379119 508178 379485
rect 508118 379085 508131 379119
rect 508165 379085 508178 379119
rect 508118 378719 508178 379085
rect 508118 378685 508131 378719
rect 508165 378685 508178 378719
rect 508118 378319 508178 378685
rect 508118 378285 508131 378319
rect 508165 378285 508178 378319
rect 508118 377919 508178 378285
rect 508118 377885 508131 377919
rect 508165 377885 508178 377919
rect 498718 377707 498731 377741
rect 498765 377707 498778 377741
rect 498718 377341 498778 377707
rect 498718 377307 498731 377341
rect 498765 377307 498778 377341
rect 498718 376941 498778 377307
rect 498718 376907 498731 376941
rect 498765 376907 498778 376941
rect 498718 376541 498778 376907
rect 498718 376507 498731 376541
rect 498765 376507 498778 376541
rect 498718 376141 498778 376507
rect 498718 376107 498731 376141
rect 498765 376107 498778 376141
rect 498718 375741 498778 376107
rect 498718 375707 498731 375741
rect 498765 375707 498778 375741
rect 498718 375341 498778 375707
rect 498718 375307 498731 375341
rect 498765 375307 498778 375341
rect 498718 374941 498778 375307
rect 498718 374907 498731 374941
rect 498765 374907 498778 374941
rect 498718 374541 498778 374907
rect 498718 374507 498731 374541
rect 498765 374507 498778 374541
rect 498718 374141 498778 374507
rect 498718 374107 498731 374141
rect 498765 374107 498778 374141
rect 498718 373741 498778 374107
rect 498718 373707 498731 373741
rect 498765 373707 498778 373741
rect 498718 373341 498778 373707
rect 500598 377495 500658 377776
rect 502478 377748 502538 377776
rect 502268 377735 502538 377748
rect 502268 377701 502351 377735
rect 502385 377701 502538 377735
rect 502268 377688 502538 377701
rect 500598 377461 500611 377495
rect 500645 377461 500658 377495
rect 500598 377095 500658 377461
rect 500598 377061 500611 377095
rect 500645 377061 500658 377095
rect 500598 376695 500658 377061
rect 500598 376661 500611 376695
rect 500645 376661 500658 376695
rect 500598 376295 500658 376661
rect 500598 376261 500611 376295
rect 500645 376261 500658 376295
rect 500598 375895 500658 376261
rect 500598 375861 500611 375895
rect 500645 375861 500658 375895
rect 500598 375495 500658 375861
rect 500598 375461 500611 375495
rect 500645 375461 500658 375495
rect 500598 375095 500658 375461
rect 500598 375061 500611 375095
rect 500645 375061 500658 375095
rect 500598 374695 500658 375061
rect 500598 374661 500611 374695
rect 500645 374661 500658 374695
rect 500598 374295 500658 374661
rect 500598 374261 500611 374295
rect 500645 374261 500658 374295
rect 500598 373895 500658 374261
rect 500598 373861 500611 373895
rect 500645 373861 500658 373895
rect 500598 373498 500658 373861
rect 500758 377209 500818 377678
rect 501978 377667 502038 377678
rect 501854 377666 502038 377667
rect 501104 377632 501131 377666
rect 501185 377632 501203 377666
rect 501253 377632 501275 377666
rect 501321 377632 501347 377666
rect 501389 377632 501419 377666
rect 501457 377632 501491 377666
rect 501525 377632 501559 377666
rect 501597 377632 501627 377666
rect 501669 377632 501695 377666
rect 501741 377632 501763 377666
rect 501813 377632 501831 377666
rect 501885 377633 502038 377666
rect 501885 377632 501912 377633
rect 500758 377208 501122 377209
rect 500758 377175 501131 377208
rect 500758 376293 500818 377175
rect 501104 377174 501131 377175
rect 501185 377174 501203 377208
rect 501253 377174 501275 377208
rect 501321 377174 501347 377208
rect 501389 377174 501419 377208
rect 501457 377174 501491 377208
rect 501525 377174 501559 377208
rect 501597 377174 501627 377208
rect 501669 377174 501695 377208
rect 501741 377174 501763 377208
rect 501813 377174 501831 377208
rect 501885 377174 501912 377208
rect 501978 376751 502038 377633
rect 501854 376750 502038 376751
rect 501104 376716 501131 376750
rect 501185 376716 501203 376750
rect 501253 376716 501275 376750
rect 501321 376716 501347 376750
rect 501389 376716 501419 376750
rect 501457 376716 501491 376750
rect 501525 376716 501559 376750
rect 501597 376716 501627 376750
rect 501669 376716 501695 376750
rect 501741 376716 501763 376750
rect 501813 376716 501831 376750
rect 501885 376717 502038 376750
rect 501885 376716 501912 376717
rect 500758 376292 501122 376293
rect 500758 376259 501131 376292
rect 500758 375377 500818 376259
rect 501104 376258 501131 376259
rect 501185 376258 501203 376292
rect 501253 376258 501275 376292
rect 501321 376258 501347 376292
rect 501389 376258 501419 376292
rect 501457 376258 501491 376292
rect 501525 376258 501559 376292
rect 501597 376258 501627 376292
rect 501669 376258 501695 376292
rect 501741 376258 501763 376292
rect 501813 376258 501831 376292
rect 501885 376258 501912 376292
rect 501978 375835 502038 376717
rect 501854 375834 502038 375835
rect 501104 375800 501131 375834
rect 501185 375800 501203 375834
rect 501253 375800 501275 375834
rect 501321 375800 501347 375834
rect 501389 375800 501419 375834
rect 501457 375800 501491 375834
rect 501525 375800 501559 375834
rect 501597 375800 501627 375834
rect 501669 375800 501695 375834
rect 501741 375800 501763 375834
rect 501813 375800 501831 375834
rect 501885 375801 502038 375834
rect 501885 375800 501912 375801
rect 500758 375376 501122 375377
rect 500758 375343 501131 375376
rect 500758 374461 500818 375343
rect 501104 375342 501131 375343
rect 501185 375342 501203 375376
rect 501253 375342 501275 375376
rect 501321 375342 501347 375376
rect 501389 375342 501419 375376
rect 501457 375342 501491 375376
rect 501525 375342 501559 375376
rect 501597 375342 501627 375376
rect 501669 375342 501695 375376
rect 501741 375342 501763 375376
rect 501813 375342 501831 375376
rect 501885 375342 501912 375376
rect 501978 374919 502038 375801
rect 501854 374918 502038 374919
rect 501104 374884 501131 374918
rect 501185 374884 501203 374918
rect 501253 374884 501275 374918
rect 501321 374884 501347 374918
rect 501389 374884 501419 374918
rect 501457 374884 501491 374918
rect 501525 374884 501559 374918
rect 501597 374884 501627 374918
rect 501669 374884 501695 374918
rect 501741 374884 501763 374918
rect 501813 374884 501831 374918
rect 501885 374885 502038 374918
rect 501885 374884 501912 374885
rect 500758 374460 501122 374461
rect 500758 374427 501131 374460
rect 500758 373545 500818 374427
rect 501104 374426 501131 374427
rect 501185 374426 501203 374460
rect 501253 374426 501275 374460
rect 501321 374426 501347 374460
rect 501389 374426 501419 374460
rect 501457 374426 501491 374460
rect 501525 374426 501559 374460
rect 501597 374426 501627 374460
rect 501669 374426 501695 374460
rect 501741 374426 501763 374460
rect 501813 374426 501831 374460
rect 501885 374426 501912 374460
rect 501978 374003 502038 374885
rect 501854 374002 502038 374003
rect 501104 373968 501131 374002
rect 501185 373968 501203 374002
rect 501253 373968 501275 374002
rect 501321 373968 501347 374002
rect 501389 373968 501419 374002
rect 501457 373968 501491 374002
rect 501525 373968 501559 374002
rect 501597 373968 501627 374002
rect 501669 373968 501695 374002
rect 501741 373968 501763 374002
rect 501813 373968 501831 374002
rect 501885 373969 502038 374002
rect 501885 373968 501912 373969
rect 500758 373544 501122 373545
rect 500758 373511 501131 373544
rect 500758 373498 500818 373511
rect 501104 373510 501131 373511
rect 501185 373510 501203 373544
rect 501253 373510 501275 373544
rect 501321 373510 501347 373544
rect 501389 373510 501419 373544
rect 501457 373510 501491 373544
rect 501525 373510 501559 373544
rect 501597 373510 501627 373544
rect 501669 373510 501695 373544
rect 501741 373510 501763 373544
rect 501813 373510 501831 373544
rect 501885 373510 501912 373544
rect 501978 373498 502038 373969
rect 502144 377495 502204 377598
rect 502144 377461 502157 377495
rect 502191 377461 502204 377495
rect 502144 377095 502204 377461
rect 502144 377061 502157 377095
rect 502191 377061 502204 377095
rect 502144 376695 502204 377061
rect 502478 377495 502538 377688
rect 502478 377461 502491 377495
rect 502525 377461 502538 377495
rect 502478 377095 502538 377461
rect 502478 377061 502491 377095
rect 502525 377061 502538 377095
rect 502478 376698 502538 377061
rect 502144 376661 502157 376695
rect 502191 376661 502204 376695
rect 502144 376295 502204 376661
rect 502358 376695 502538 376698
rect 502358 376661 502491 376695
rect 502525 376661 502538 376695
rect 502358 376633 502538 376661
rect 502358 376599 502381 376633
rect 502415 376599 502538 376633
rect 502358 376538 502538 376599
rect 502144 376261 502157 376295
rect 502191 376261 502204 376295
rect 502144 375895 502204 376261
rect 502144 375861 502157 375895
rect 502191 375861 502204 375895
rect 502144 375495 502204 375861
rect 502144 375461 502157 375495
rect 502191 375461 502204 375495
rect 502144 375095 502204 375461
rect 502478 376295 502538 376538
rect 502478 376261 502491 376295
rect 502525 376261 502538 376295
rect 502478 375895 502538 376261
rect 502478 375861 502491 375895
rect 502525 375861 502538 375895
rect 502478 375495 502538 375861
rect 502478 375461 502491 375495
rect 502525 375461 502538 375495
rect 502478 375398 502538 375461
rect 502358 375333 502538 375398
rect 502358 375299 502381 375333
rect 502415 375299 502538 375333
rect 502358 375238 502538 375299
rect 502144 375061 502157 375095
rect 502191 375061 502204 375095
rect 502144 374695 502204 375061
rect 502144 374661 502157 374695
rect 502191 374661 502204 374695
rect 502144 374295 502204 374661
rect 502144 374261 502157 374295
rect 502191 374261 502204 374295
rect 502144 373895 502204 374261
rect 502144 373861 502157 373895
rect 502191 373861 502204 373895
rect 502144 373525 502204 373861
rect 502144 373498 502161 373525
rect 502195 373498 502204 373525
rect 502478 375095 502538 375238
rect 502478 375061 502491 375095
rect 502525 375061 502538 375095
rect 502478 374695 502538 375061
rect 502478 374661 502491 374695
rect 502525 374661 502538 374695
rect 502478 374295 502538 374661
rect 504358 377552 504418 377580
rect 504358 377539 504628 377552
rect 504358 377505 504511 377539
rect 504545 377505 504628 377539
rect 504358 377492 504628 377505
rect 504358 377299 504418 377492
rect 505998 377435 506058 377482
rect 504358 377265 504371 377299
rect 504405 377265 504418 377299
rect 504358 376899 504418 377265
rect 504358 376865 504371 376899
rect 504405 376865 504418 376899
rect 504358 376504 504418 376865
rect 504538 377389 504578 377422
rect 504619 377401 504639 377435
rect 504673 377401 504707 377435
rect 504745 377401 504775 377435
rect 504817 377401 504843 377435
rect 504889 377401 504911 377435
rect 504961 377401 504979 377435
rect 505033 377401 505047 377435
rect 505105 377401 505115 377435
rect 505177 377401 505183 377435
rect 505249 377401 505251 377435
rect 505285 377401 505287 377435
rect 505353 377401 505359 377435
rect 505421 377401 505431 377435
rect 505489 377401 505503 377435
rect 505557 377401 505575 377435
rect 505625 377401 505647 377435
rect 505693 377401 505719 377435
rect 505761 377401 505791 377435
rect 505829 377401 505863 377435
rect 505897 377401 506058 377435
rect 504538 377355 504541 377389
rect 504575 377355 504578 377389
rect 504538 376977 504578 377355
rect 505998 377389 506058 377401
rect 505998 377355 506003 377389
rect 506037 377355 506058 377389
rect 504538 376943 504639 376977
rect 504673 376943 504707 376977
rect 504745 376943 504775 376977
rect 504817 376943 504843 376977
rect 504889 376943 504911 376977
rect 504961 376943 504979 376977
rect 505033 376943 505047 376977
rect 505105 376943 505115 376977
rect 505177 376943 505183 376977
rect 505249 376943 505251 376977
rect 505285 376943 505287 376977
rect 505353 376943 505359 376977
rect 505421 376943 505431 376977
rect 505489 376943 505503 376977
rect 505557 376943 505575 376977
rect 505625 376943 505647 376977
rect 505693 376943 505719 376977
rect 505761 376943 505791 376977
rect 505829 376943 505863 376977
rect 505897 376943 505917 376977
rect 504358 376499 504498 376504
rect 504358 376465 504371 376499
rect 504405 376465 504498 376499
rect 504358 376439 504498 376465
rect 504358 376405 504461 376439
rect 504495 376405 504498 376439
rect 504358 376344 504498 376405
rect 504358 376099 504418 376344
rect 504358 376065 504371 376099
rect 504405 376065 504418 376099
rect 504358 375699 504418 376065
rect 504358 375665 504371 375699
rect 504405 375665 504418 375699
rect 504358 375299 504418 375665
rect 504358 375265 504371 375299
rect 504405 375265 504418 375299
rect 504358 374899 504418 375265
rect 504358 374865 504371 374899
rect 504405 374865 504418 374899
rect 504358 374606 504418 374865
rect 504538 376061 504578 376943
rect 505998 376519 506058 377355
rect 504619 376485 504639 376519
rect 504673 376485 504707 376519
rect 504745 376485 504775 376519
rect 504817 376485 504843 376519
rect 504889 376485 504911 376519
rect 504961 376485 504979 376519
rect 505033 376485 505047 376519
rect 505105 376485 505115 376519
rect 505177 376485 505183 376519
rect 505249 376485 505251 376519
rect 505285 376485 505287 376519
rect 505353 376485 505359 376519
rect 505421 376485 505431 376519
rect 505489 376485 505503 376519
rect 505557 376485 505575 376519
rect 505625 376485 505647 376519
rect 505693 376485 505719 376519
rect 505761 376485 505791 376519
rect 505829 376485 505863 376519
rect 505897 376485 506058 376519
rect 504538 376027 504639 376061
rect 504673 376027 504707 376061
rect 504745 376027 504775 376061
rect 504817 376027 504843 376061
rect 504889 376027 504911 376061
rect 504961 376027 504979 376061
rect 505033 376027 505047 376061
rect 505105 376027 505115 376061
rect 505177 376027 505183 376061
rect 505249 376027 505251 376061
rect 505285 376027 505287 376061
rect 505353 376027 505359 376061
rect 505421 376027 505431 376061
rect 505489 376027 505503 376061
rect 505557 376027 505575 376061
rect 505625 376027 505647 376061
rect 505693 376027 505719 376061
rect 505761 376027 505791 376061
rect 505829 376027 505863 376061
rect 505897 376027 505917 376061
rect 504538 375145 504578 376027
rect 505998 375603 506058 376485
rect 504619 375569 504639 375603
rect 504673 375569 504707 375603
rect 504745 375569 504775 375603
rect 504817 375569 504843 375603
rect 504889 375569 504911 375603
rect 504961 375569 504979 375603
rect 505033 375569 505047 375603
rect 505105 375569 505115 375603
rect 505177 375569 505183 375603
rect 505249 375569 505251 375603
rect 505285 375569 505287 375603
rect 505353 375569 505359 375603
rect 505421 375569 505431 375603
rect 505489 375569 505503 375603
rect 505557 375569 505575 375603
rect 505625 375569 505647 375603
rect 505693 375569 505719 375603
rect 505761 375569 505791 375603
rect 505829 375569 505863 375603
rect 505897 375569 506058 375603
rect 504538 375111 504639 375145
rect 504673 375111 504707 375145
rect 504745 375111 504775 375145
rect 504817 375111 504843 375145
rect 504889 375111 504911 375145
rect 504961 375111 504979 375145
rect 505033 375111 505047 375145
rect 505105 375111 505115 375145
rect 505177 375111 505183 375145
rect 505249 375111 505251 375145
rect 505285 375111 505287 375145
rect 505353 375111 505359 375145
rect 505421 375111 505431 375145
rect 505489 375111 505503 375145
rect 505557 375111 505575 375145
rect 505625 375111 505647 375145
rect 505693 375111 505719 375145
rect 505761 375111 505791 375145
rect 505829 375111 505863 375145
rect 505897 375111 505917 375145
rect 504538 374606 504578 375111
rect 505998 374687 506058 375569
rect 504619 374653 504639 374687
rect 504673 374653 504707 374687
rect 504745 374653 504775 374687
rect 504817 374653 504843 374687
rect 504889 374653 504911 374687
rect 504961 374653 504979 374687
rect 505033 374653 505047 374687
rect 505105 374653 505115 374687
rect 505177 374653 505183 374687
rect 505249 374653 505251 374687
rect 505285 374653 505287 374687
rect 505353 374653 505359 374687
rect 505421 374653 505431 374687
rect 505489 374653 505503 374687
rect 505557 374653 505575 374687
rect 505625 374653 505647 374687
rect 505693 374653 505719 374687
rect 505761 374653 505791 374687
rect 505829 374653 505863 374687
rect 505897 374653 506058 374687
rect 505998 374606 506058 374653
rect 506104 377299 506164 377482
rect 506104 377265 506117 377299
rect 506151 377265 506164 377299
rect 506104 376899 506164 377265
rect 506104 376865 506117 376899
rect 506151 376865 506164 376899
rect 506104 376499 506164 376865
rect 506104 376465 506117 376499
rect 506151 376465 506164 376499
rect 506104 376377 506164 376465
rect 506104 376343 506105 376377
rect 506139 376343 506164 376377
rect 506104 376099 506164 376343
rect 506104 376065 506117 376099
rect 506151 376065 506164 376099
rect 506104 375699 506164 376065
rect 506104 375665 506117 375699
rect 506151 375665 506164 375699
rect 506104 375299 506164 375665
rect 506104 375265 506117 375299
rect 506151 375265 506164 375299
rect 506104 374899 506164 375265
rect 506104 374865 506117 374899
rect 506151 374865 506164 374899
rect 506104 374606 506164 374865
rect 506238 377299 506298 377580
rect 506238 377265 506251 377299
rect 506285 377265 506298 377299
rect 506238 376899 506298 377265
rect 506238 376865 506251 376899
rect 506285 376865 506298 376899
rect 506238 376499 506298 376865
rect 506238 376465 506251 376499
rect 506285 376465 506298 376499
rect 506238 376099 506298 376465
rect 506238 376065 506251 376099
rect 506285 376065 506298 376099
rect 506238 375699 506298 376065
rect 506238 375665 506251 375699
rect 506285 375665 506298 375699
rect 506238 375299 506298 375665
rect 506238 375265 506251 375299
rect 506285 375265 506298 375299
rect 506238 374899 506298 375265
rect 506238 374865 506251 374899
rect 506285 374865 506298 374899
rect 506238 374606 506298 374865
rect 508118 377519 508178 377885
rect 508118 377485 508131 377519
rect 508165 377485 508178 377519
rect 508118 377119 508178 377485
rect 508118 377085 508131 377119
rect 508165 377085 508178 377119
rect 508118 376719 508178 377085
rect 508118 376685 508131 376719
rect 508165 376685 508178 376719
rect 508118 376319 508178 376685
rect 508118 376285 508131 376319
rect 508165 376285 508178 376319
rect 508118 375919 508178 376285
rect 508118 375885 508131 375919
rect 508165 375885 508178 375919
rect 508118 375519 508178 375885
rect 508118 375485 508131 375519
rect 508165 375485 508178 375519
rect 508118 375119 508178 375485
rect 508118 375085 508131 375119
rect 508165 375085 508178 375119
rect 508118 374719 508178 375085
rect 508118 374685 508131 374719
rect 508165 374685 508178 374719
rect 502478 374261 502491 374295
rect 502525 374261 502538 374295
rect 502478 373895 502538 374261
rect 508118 374319 508178 374685
rect 508118 374285 508131 374319
rect 508165 374285 508178 374319
rect 508118 374134 508178 374285
rect 509998 381119 510058 381302
rect 509998 381085 510011 381119
rect 510045 381085 510058 381119
rect 509998 380719 510058 381085
rect 509998 380685 510011 380719
rect 510045 380685 510058 380719
rect 509998 380319 510058 380685
rect 509998 380285 510011 380319
rect 510045 380285 510058 380319
rect 509998 379919 510058 380285
rect 509998 379885 510011 379919
rect 510045 379885 510058 379919
rect 509998 379519 510058 379885
rect 509998 379485 510011 379519
rect 510045 379485 510058 379519
rect 509998 379119 510058 379485
rect 509998 379085 510011 379119
rect 510045 379085 510058 379119
rect 509998 378719 510058 379085
rect 509998 378685 510011 378719
rect 510045 378685 510058 378719
rect 509998 378319 510058 378685
rect 509998 378285 510011 378319
rect 510045 378285 510058 378319
rect 509998 377919 510058 378285
rect 509998 377885 510011 377919
rect 510045 377885 510058 377919
rect 509998 377519 510058 377885
rect 511878 381243 511938 381609
rect 511878 381209 511891 381243
rect 511925 381209 511938 381243
rect 511878 380843 511938 381209
rect 511878 380809 511891 380843
rect 511925 380809 511938 380843
rect 511878 380443 511938 380809
rect 511878 380409 511891 380443
rect 511925 380409 511938 380443
rect 511878 380043 511938 380409
rect 511878 380009 511891 380043
rect 511925 380009 511938 380043
rect 511878 379643 511938 380009
rect 511878 379609 511891 379643
rect 511925 379609 511938 379643
rect 511878 379243 511938 379609
rect 511878 379209 511891 379243
rect 511925 379209 511938 379243
rect 511878 378843 511938 379209
rect 511878 378809 511891 378843
rect 511925 378809 511938 378843
rect 511878 378443 511938 378809
rect 511878 378409 511891 378443
rect 511925 378409 511938 378443
rect 511878 378043 511938 378409
rect 511878 378009 511891 378043
rect 511925 378009 511938 378043
rect 511878 377858 511938 378009
rect 513758 384843 513818 385026
rect 513758 384809 513771 384843
rect 513805 384809 513818 384843
rect 513758 384443 513818 384809
rect 513758 384409 513771 384443
rect 513805 384409 513818 384443
rect 513758 384043 513818 384409
rect 513758 384009 513771 384043
rect 513805 384009 513818 384043
rect 513758 383643 513818 384009
rect 513758 383609 513771 383643
rect 513805 383609 513818 383643
rect 513758 383243 513818 383609
rect 513758 383209 513771 383243
rect 513805 383209 513818 383243
rect 513758 382843 513818 383209
rect 513758 382809 513771 382843
rect 513805 382809 513818 382843
rect 513758 382443 513818 382809
rect 513758 382409 513771 382443
rect 513805 382409 513818 382443
rect 513758 382043 513818 382409
rect 513758 382009 513771 382043
rect 513805 382009 513818 382043
rect 513758 381643 513818 382009
rect 513758 381609 513771 381643
rect 513805 381609 513818 381643
rect 513758 381243 513818 381609
rect 513758 381209 513771 381243
rect 513805 381209 513818 381243
rect 513758 380843 513818 381209
rect 513758 380809 513771 380843
rect 513805 380809 513818 380843
rect 513758 380443 513818 380809
rect 513758 380409 513771 380443
rect 513805 380409 513818 380443
rect 513758 380043 513818 380409
rect 513758 380009 513771 380043
rect 513805 380009 513818 380043
rect 513758 379643 513818 380009
rect 513758 379609 513771 379643
rect 513805 379609 513818 379643
rect 513758 379243 513818 379609
rect 513758 379209 513771 379243
rect 513805 379209 513818 379243
rect 513758 378843 513818 379209
rect 513758 378809 513771 378843
rect 513805 378809 513818 378843
rect 513758 378443 513818 378809
rect 513758 378409 513771 378443
rect 513805 378409 513818 378443
rect 513758 378043 513818 378409
rect 513758 378009 513771 378043
rect 513805 378009 513818 378043
rect 513758 377858 513818 378009
rect 515638 384843 515698 385026
rect 515638 384809 515651 384843
rect 515685 384809 515698 384843
rect 515638 384443 515698 384809
rect 515638 384409 515651 384443
rect 515685 384409 515698 384443
rect 515638 384043 515698 384409
rect 515638 384009 515651 384043
rect 515685 384009 515698 384043
rect 515638 383643 515698 384009
rect 515638 383609 515651 383643
rect 515685 383609 515698 383643
rect 515638 383243 515698 383609
rect 515638 383209 515651 383243
rect 515685 383209 515698 383243
rect 515638 382843 515698 383209
rect 515638 382809 515651 382843
rect 515685 382809 515698 382843
rect 515638 382443 515698 382809
rect 515638 382409 515651 382443
rect 515685 382409 515698 382443
rect 515638 382043 515698 382409
rect 515638 382009 515651 382043
rect 515685 382009 515698 382043
rect 515638 381643 515698 382009
rect 515638 381609 515651 381643
rect 515685 381609 515698 381643
rect 515638 381243 515698 381609
rect 515638 381209 515651 381243
rect 515685 381209 515698 381243
rect 515638 380843 515698 381209
rect 515638 380809 515651 380843
rect 515685 380809 515698 380843
rect 515638 380443 515698 380809
rect 515638 380409 515651 380443
rect 515685 380409 515698 380443
rect 515638 380043 515698 380409
rect 515638 380009 515651 380043
rect 515685 380009 515698 380043
rect 515638 379643 515698 380009
rect 515638 379609 515651 379643
rect 515685 379609 515698 379643
rect 515638 379243 515698 379609
rect 515638 379209 515651 379243
rect 515685 379209 515698 379243
rect 515638 378843 515698 379209
rect 515638 378809 515651 378843
rect 515685 378809 515698 378843
rect 515638 378443 515698 378809
rect 515638 378409 515651 378443
rect 515685 378409 515698 378443
rect 515638 378043 515698 378409
rect 515638 378009 515651 378043
rect 515685 378009 515698 378043
rect 515638 377858 515698 378009
rect 517518 384843 517578 385026
rect 517518 384809 517531 384843
rect 517565 384809 517578 384843
rect 517518 384443 517578 384809
rect 517518 384409 517531 384443
rect 517565 384409 517578 384443
rect 517518 384043 517578 384409
rect 517518 384009 517531 384043
rect 517565 384009 517578 384043
rect 517518 383643 517578 384009
rect 517518 383609 517531 383643
rect 517565 383609 517578 383643
rect 517518 383243 517578 383609
rect 517518 383209 517531 383243
rect 517565 383209 517578 383243
rect 517518 382843 517578 383209
rect 517518 382809 517531 382843
rect 517565 382809 517578 382843
rect 517518 382443 517578 382809
rect 519398 384825 519458 385008
rect 519398 384791 519411 384825
rect 519445 384791 519458 384825
rect 519398 384625 519458 384791
rect 519398 384591 519411 384625
rect 519445 384591 519458 384625
rect 519398 384425 519458 384591
rect 521278 384825 521338 385008
rect 521278 384791 521291 384825
rect 521325 384791 521338 384825
rect 521278 384625 521338 384791
rect 521278 384591 521291 384625
rect 521325 384591 521338 384625
rect 519398 384391 519411 384425
rect 519445 384391 519458 384425
rect 519398 384225 519458 384391
rect 519398 384191 519411 384225
rect 519445 384191 519458 384225
rect 519398 384025 519458 384191
rect 521278 384425 521338 384591
rect 521278 384391 521291 384425
rect 521325 384391 521338 384425
rect 521278 384225 521338 384391
rect 521278 384191 521291 384225
rect 521325 384191 521338 384225
rect 521278 384096 521338 384191
rect 519398 383991 519411 384025
rect 519445 383991 519458 384025
rect 519398 383825 519458 383991
rect 519398 383791 519411 383825
rect 519445 383791 519458 383825
rect 519398 383625 519458 383791
rect 519398 383591 519411 383625
rect 519445 383591 519458 383625
rect 519398 383425 519458 383591
rect 520338 384025 521338 384096
rect 520338 384009 521291 384025
rect 520338 383567 520377 384009
rect 520479 383991 521291 384009
rect 521325 383991 521338 384025
rect 520479 383825 521338 383991
rect 520479 383791 521291 383825
rect 521325 383791 521338 383825
rect 520479 383625 521338 383791
rect 520479 383591 521291 383625
rect 521325 383591 521338 383625
rect 520479 383567 521338 383591
rect 520338 383480 521338 383567
rect 519398 383391 519411 383425
rect 519445 383391 519458 383425
rect 519398 383225 519458 383391
rect 519398 383191 519411 383225
rect 519445 383191 519458 383225
rect 519398 383025 519458 383191
rect 519398 382991 519411 383025
rect 519445 382991 519458 383025
rect 521278 383425 521338 383480
rect 521278 383391 521291 383425
rect 521325 383391 521338 383425
rect 521278 383225 521338 383391
rect 521278 383191 521291 383225
rect 521325 383191 521338 383225
rect 521278 383025 521338 383191
rect 519398 382825 519458 382991
rect 519398 382791 519411 382825
rect 519445 382791 519458 382825
rect 519398 382568 519458 382791
rect 520233 382568 520623 383000
rect 521278 382991 521291 383025
rect 521325 382991 521338 383025
rect 521278 382825 521338 382991
rect 521278 382791 521291 382825
rect 521325 382791 521338 382825
rect 521278 382568 521338 382791
rect 523158 384741 523218 385086
rect 523158 384707 523171 384741
rect 523205 384707 523218 384741
rect 523158 384341 523218 384707
rect 523158 384307 523171 384341
rect 523205 384307 523218 384341
rect 523158 383946 523218 384307
rect 523338 385039 523378 385921
rect 524798 385497 524858 386379
rect 523419 385463 523439 385497
rect 523473 385463 523507 385497
rect 523545 385463 523575 385497
rect 523617 385463 523643 385497
rect 523689 385463 523711 385497
rect 523761 385463 523779 385497
rect 523833 385463 523847 385497
rect 523905 385463 523915 385497
rect 523977 385463 523983 385497
rect 524049 385463 524051 385497
rect 524085 385463 524087 385497
rect 524153 385463 524159 385497
rect 524221 385463 524231 385497
rect 524289 385463 524303 385497
rect 524357 385463 524375 385497
rect 524425 385463 524447 385497
rect 524493 385463 524519 385497
rect 524561 385463 524591 385497
rect 524629 385463 524663 385497
rect 524697 385463 524858 385497
rect 523338 385005 523439 385039
rect 523473 385005 523507 385039
rect 523545 385005 523575 385039
rect 523617 385005 523643 385039
rect 523689 385005 523711 385039
rect 523761 385005 523779 385039
rect 523833 385005 523847 385039
rect 523905 385005 523915 385039
rect 523977 385005 523983 385039
rect 524049 385005 524051 385039
rect 524085 385005 524087 385039
rect 524153 385005 524159 385039
rect 524221 385005 524231 385039
rect 524289 385005 524303 385039
rect 524357 385005 524375 385039
rect 524425 385005 524447 385039
rect 524493 385005 524519 385039
rect 524561 385005 524591 385039
rect 524629 385005 524663 385039
rect 524697 385005 524717 385039
rect 523338 384123 523378 385005
rect 524798 384581 524858 385463
rect 523419 384547 523439 384581
rect 523473 384547 523507 384581
rect 523545 384547 523575 384581
rect 523617 384547 523643 384581
rect 523689 384547 523711 384581
rect 523761 384547 523779 384581
rect 523833 384547 523847 384581
rect 523905 384547 523915 384581
rect 523977 384547 523983 384581
rect 524049 384547 524051 384581
rect 524085 384547 524087 384581
rect 524153 384547 524159 384581
rect 524221 384547 524231 384581
rect 524289 384547 524303 384581
rect 524357 384547 524375 384581
rect 524425 384547 524447 384581
rect 524493 384547 524519 384581
rect 524561 384547 524591 384581
rect 524629 384547 524663 384581
rect 524697 384547 524858 384581
rect 523338 384089 523439 384123
rect 523473 384089 523507 384123
rect 523545 384089 523575 384123
rect 523617 384089 523643 384123
rect 523689 384089 523711 384123
rect 523761 384089 523779 384123
rect 523833 384089 523847 384123
rect 523905 384089 523915 384123
rect 523977 384089 523983 384123
rect 524049 384089 524051 384123
rect 524085 384089 524087 384123
rect 524153 384089 524159 384123
rect 524221 384089 524231 384123
rect 524289 384089 524303 384123
rect 524357 384089 524375 384123
rect 524425 384089 524447 384123
rect 524493 384089 524519 384123
rect 524561 384089 524591 384123
rect 524629 384089 524663 384123
rect 524697 384089 524717 384123
rect 523158 383941 523298 383946
rect 523158 383907 523171 383941
rect 523205 383907 523298 383941
rect 523158 383881 523298 383907
rect 523158 383847 523261 383881
rect 523295 383847 523298 383881
rect 523158 383786 523298 383847
rect 523158 383541 523218 383786
rect 523158 383507 523171 383541
rect 523205 383507 523218 383541
rect 523158 383141 523218 383507
rect 523158 383107 523171 383141
rect 523205 383107 523218 383141
rect 523158 382741 523218 383107
rect 523158 382707 523171 382741
rect 523205 382707 523218 382741
rect 523158 382646 523218 382707
rect 523338 383207 523378 384089
rect 524798 383665 524858 384547
rect 523419 383631 523439 383665
rect 523473 383631 523507 383665
rect 523545 383631 523575 383665
rect 523617 383631 523643 383665
rect 523689 383631 523711 383665
rect 523761 383631 523779 383665
rect 523833 383631 523847 383665
rect 523905 383631 523915 383665
rect 523977 383631 523983 383665
rect 524049 383631 524051 383665
rect 524085 383631 524087 383665
rect 524153 383631 524159 383665
rect 524221 383631 524231 383665
rect 524289 383631 524303 383665
rect 524357 383631 524375 383665
rect 524425 383631 524447 383665
rect 524493 383631 524519 383665
rect 524561 383631 524591 383665
rect 524629 383631 524663 383665
rect 524697 383631 524858 383665
rect 523338 383173 523439 383207
rect 523473 383173 523507 383207
rect 523545 383173 523575 383207
rect 523617 383173 523643 383207
rect 523689 383173 523711 383207
rect 523761 383173 523779 383207
rect 523833 383173 523847 383207
rect 523905 383173 523915 383207
rect 523977 383173 523983 383207
rect 524049 383173 524051 383207
rect 524085 383173 524087 383207
rect 524153 383173 524159 383207
rect 524221 383173 524231 383207
rect 524289 383173 524303 383207
rect 524357 383173 524375 383207
rect 524425 383173 524447 383207
rect 524493 383173 524519 383207
rect 524561 383173 524591 383207
rect 524629 383173 524663 383207
rect 524697 383173 524717 383207
rect 523158 382581 523298 382646
rect 517518 382409 517531 382443
rect 517565 382409 517578 382443
rect 517518 382043 517578 382409
rect 517518 382009 517531 382043
rect 517565 382009 517578 382043
rect 517518 381643 517578 382009
rect 523158 382547 523261 382581
rect 523295 382547 523298 382581
rect 523158 382486 523298 382547
rect 523158 382341 523218 382486
rect 523158 382307 523171 382341
rect 523205 382307 523218 382341
rect 523158 381941 523218 382307
rect 523158 381907 523171 381941
rect 523205 381907 523218 381941
rect 517518 381609 517531 381643
rect 517565 381609 517578 381643
rect 517518 381243 517578 381609
rect 517518 381209 517531 381243
rect 517565 381209 517578 381243
rect 517518 380843 517578 381209
rect 517518 380809 517531 380843
rect 517565 380809 517578 380843
rect 517518 380443 517578 380809
rect 517518 380409 517531 380443
rect 517565 380409 517578 380443
rect 517518 380043 517578 380409
rect 517518 380009 517531 380043
rect 517565 380009 517578 380043
rect 517518 379643 517578 380009
rect 517518 379609 517531 379643
rect 517565 379609 517578 379643
rect 517518 379243 517578 379609
rect 519398 381591 519458 381774
rect 519398 381557 519411 381591
rect 519445 381557 519458 381591
rect 519398 381391 519458 381557
rect 519398 381357 519411 381391
rect 519445 381357 519458 381391
rect 519398 381191 519458 381357
rect 521278 381591 521338 381774
rect 521278 381557 521291 381591
rect 521325 381557 521338 381591
rect 521278 381391 521338 381557
rect 521278 381357 521291 381391
rect 521325 381357 521338 381391
rect 519398 381157 519411 381191
rect 519445 381157 519458 381191
rect 519398 380991 519458 381157
rect 519398 380957 519411 380991
rect 519445 380957 519458 380991
rect 519398 380791 519458 380957
rect 521278 381191 521338 381357
rect 521278 381157 521291 381191
rect 521325 381157 521338 381191
rect 521278 380991 521338 381157
rect 521278 380957 521291 380991
rect 521325 380957 521338 380991
rect 521278 380862 521338 380957
rect 519398 380757 519411 380791
rect 519445 380757 519458 380791
rect 519398 380591 519458 380757
rect 519398 380557 519411 380591
rect 519445 380557 519458 380591
rect 519398 380391 519458 380557
rect 519398 380357 519411 380391
rect 519445 380357 519458 380391
rect 519398 380191 519458 380357
rect 520338 380791 521338 380862
rect 520338 380775 521291 380791
rect 520338 380333 520377 380775
rect 520479 380757 521291 380775
rect 521325 380757 521338 380791
rect 520479 380591 521338 380757
rect 520479 380557 521291 380591
rect 521325 380557 521338 380591
rect 520479 380391 521338 380557
rect 520479 380357 521291 380391
rect 521325 380357 521338 380391
rect 520479 380333 521338 380357
rect 520338 380246 521338 380333
rect 519398 380157 519411 380191
rect 519445 380157 519458 380191
rect 519398 379991 519458 380157
rect 519398 379957 519411 379991
rect 519445 379957 519458 379991
rect 519398 379791 519458 379957
rect 519398 379757 519411 379791
rect 519445 379757 519458 379791
rect 521278 380191 521338 380246
rect 521278 380157 521291 380191
rect 521325 380157 521338 380191
rect 521278 379991 521338 380157
rect 521278 379957 521291 379991
rect 521325 379957 521338 379991
rect 521278 379791 521338 379957
rect 519398 379591 519458 379757
rect 519398 379557 519411 379591
rect 519445 379557 519458 379591
rect 519398 379334 519458 379557
rect 520233 379334 520623 379766
rect 521278 379757 521291 379791
rect 521325 379757 521338 379791
rect 521278 379591 521338 379757
rect 521278 379557 521291 379591
rect 521325 379557 521338 379591
rect 521278 379334 521338 379557
rect 523158 381541 523218 381907
rect 523158 381507 523171 381541
rect 523205 381507 523218 381541
rect 523158 381346 523218 381507
rect 523338 382291 523378 383173
rect 524798 382749 524858 383631
rect 523419 382715 523439 382749
rect 523473 382715 523507 382749
rect 523545 382715 523575 382749
rect 523617 382715 523643 382749
rect 523689 382715 523711 382749
rect 523761 382715 523779 382749
rect 523833 382715 523847 382749
rect 523905 382715 523915 382749
rect 523977 382715 523983 382749
rect 524049 382715 524051 382749
rect 524085 382715 524087 382749
rect 524153 382715 524159 382749
rect 524221 382715 524231 382749
rect 524289 382715 524303 382749
rect 524357 382715 524375 382749
rect 524425 382715 524447 382749
rect 524493 382715 524519 382749
rect 524561 382715 524591 382749
rect 524629 382715 524663 382749
rect 524697 382715 524858 382749
rect 523338 382257 523439 382291
rect 523473 382257 523507 382291
rect 523545 382257 523575 382291
rect 523617 382257 523643 382291
rect 523689 382257 523711 382291
rect 523761 382257 523779 382291
rect 523833 382257 523847 382291
rect 523905 382257 523915 382291
rect 523977 382257 523983 382291
rect 524049 382257 524051 382291
rect 524085 382257 524087 382291
rect 524153 382257 524159 382291
rect 524221 382257 524231 382291
rect 524289 382257 524303 382291
rect 524357 382257 524375 382291
rect 524425 382257 524447 382291
rect 524493 382257 524519 382291
rect 524561 382257 524591 382291
rect 524629 382257 524663 382291
rect 524697 382257 524717 382291
rect 523338 381375 523378 382257
rect 524798 381833 524858 382715
rect 523419 381799 523439 381833
rect 523473 381799 523507 381833
rect 523545 381799 523575 381833
rect 523617 381799 523643 381833
rect 523689 381799 523711 381833
rect 523761 381799 523779 381833
rect 523833 381799 523847 381833
rect 523905 381799 523915 381833
rect 523977 381799 523983 381833
rect 524049 381799 524051 381833
rect 524085 381799 524087 381833
rect 524153 381799 524159 381833
rect 524221 381799 524231 381833
rect 524289 381799 524303 381833
rect 524357 381799 524375 381833
rect 524425 381799 524447 381833
rect 524493 381799 524519 381833
rect 524561 381799 524591 381833
rect 524629 381799 524663 381833
rect 524697 381799 524858 381833
rect 523158 381281 523298 381346
rect 523158 381247 523261 381281
rect 523295 381247 523298 381281
rect 523158 381186 523298 381247
rect 523338 381341 523439 381375
rect 523473 381341 523507 381375
rect 523545 381341 523575 381375
rect 523617 381341 523643 381375
rect 523689 381341 523711 381375
rect 523761 381341 523779 381375
rect 523833 381341 523847 381375
rect 523905 381341 523915 381375
rect 523977 381341 523983 381375
rect 524049 381341 524051 381375
rect 524085 381341 524087 381375
rect 524153 381341 524159 381375
rect 524221 381341 524231 381375
rect 524289 381341 524303 381375
rect 524357 381341 524375 381375
rect 524425 381341 524447 381375
rect 524493 381341 524519 381375
rect 524561 381341 524591 381375
rect 524629 381341 524663 381375
rect 524697 381341 524717 381375
rect 523158 381141 523218 381186
rect 523158 381107 523171 381141
rect 523205 381107 523218 381141
rect 523158 380741 523218 381107
rect 523158 380707 523171 380741
rect 523205 380707 523218 380741
rect 523158 380341 523218 380707
rect 523158 380307 523171 380341
rect 523205 380307 523218 380341
rect 523158 380046 523218 380307
rect 523338 380459 523378 381341
rect 524798 380917 524858 381799
rect 523419 380883 523439 380917
rect 523473 380883 523507 380917
rect 523545 380883 523575 380917
rect 523617 380883 523643 380917
rect 523689 380883 523711 380917
rect 523761 380883 523779 380917
rect 523833 380883 523847 380917
rect 523905 380883 523915 380917
rect 523977 380883 523983 380917
rect 524049 380883 524051 380917
rect 524085 380883 524087 380917
rect 524153 380883 524159 380917
rect 524221 380883 524231 380917
rect 524289 380883 524303 380917
rect 524357 380883 524375 380917
rect 524425 380883 524447 380917
rect 524493 380883 524519 380917
rect 524561 380883 524591 380917
rect 524629 380883 524663 380917
rect 524697 380883 524858 380917
rect 524798 380609 524858 380883
rect 524798 380575 524805 380609
rect 524839 380575 524858 380609
rect 523338 380425 523439 380459
rect 523473 380425 523507 380459
rect 523545 380425 523575 380459
rect 523617 380425 523643 380459
rect 523689 380425 523711 380459
rect 523761 380425 523779 380459
rect 523833 380425 523847 380459
rect 523905 380425 523915 380459
rect 523977 380425 523983 380459
rect 524049 380425 524051 380459
rect 524085 380425 524087 380459
rect 524153 380425 524159 380459
rect 524221 380425 524231 380459
rect 524289 380425 524303 380459
rect 524357 380425 524375 380459
rect 524425 380425 524447 380459
rect 524493 380425 524519 380459
rect 524561 380425 524591 380459
rect 524629 380425 524663 380459
rect 524697 380425 524717 380459
rect 523158 379981 523298 380046
rect 523158 379947 523261 379981
rect 523295 379947 523298 379981
rect 523158 379941 523298 379947
rect 523158 379907 523171 379941
rect 523205 379907 523298 379941
rect 523158 379886 523298 379907
rect 523158 379541 523218 379886
rect 523158 379507 523171 379541
rect 523205 379507 523218 379541
rect 517518 379209 517531 379243
rect 517565 379209 517578 379243
rect 517518 378843 517578 379209
rect 517518 378809 517531 378843
rect 517565 378809 517578 378843
rect 517518 378443 517578 378809
rect 517518 378409 517531 378443
rect 517565 378409 517578 378443
rect 517518 378043 517578 378409
rect 517518 378009 517531 378043
rect 517565 378009 517578 378043
rect 517518 377858 517578 378009
rect 523158 379141 523218 379507
rect 523158 379107 523171 379141
rect 523205 379107 523218 379141
rect 523158 378746 523218 379107
rect 523338 379543 523378 380425
rect 524798 380001 524858 380575
rect 523419 379967 523439 380001
rect 523473 379967 523507 380001
rect 523545 379967 523575 380001
rect 523617 379967 523643 380001
rect 523689 379967 523711 380001
rect 523761 379967 523779 380001
rect 523833 379967 523847 380001
rect 523905 379967 523915 380001
rect 523977 379967 523983 380001
rect 524049 379967 524051 380001
rect 524085 379967 524087 380001
rect 524153 379967 524159 380001
rect 524221 379967 524231 380001
rect 524289 379967 524303 380001
rect 524357 379967 524375 380001
rect 524425 379967 524447 380001
rect 524493 379967 524519 380001
rect 524561 379967 524591 380001
rect 524629 379967 524663 380001
rect 524697 379967 524858 380001
rect 523338 379509 523439 379543
rect 523473 379509 523507 379543
rect 523545 379509 523575 379543
rect 523617 379509 523643 379543
rect 523689 379509 523711 379543
rect 523761 379509 523779 379543
rect 523833 379509 523847 379543
rect 523905 379509 523915 379543
rect 523977 379509 523983 379543
rect 524049 379509 524051 379543
rect 524085 379509 524087 379543
rect 524153 379509 524159 379543
rect 524221 379509 524231 379543
rect 524289 379509 524303 379543
rect 524357 379509 524375 379543
rect 524425 379509 524447 379543
rect 524493 379509 524519 379543
rect 524561 379509 524591 379543
rect 524629 379509 524663 379543
rect 524697 379509 524717 379543
rect 523158 378741 523298 378746
rect 523158 378707 523171 378741
rect 523205 378707 523298 378741
rect 523158 378681 523298 378707
rect 523158 378647 523261 378681
rect 523295 378647 523298 378681
rect 523158 378586 523298 378647
rect 523338 378627 523378 379509
rect 524798 379085 524858 379967
rect 523419 379051 523439 379085
rect 523473 379051 523507 379085
rect 523545 379051 523575 379085
rect 523617 379051 523643 379085
rect 523689 379051 523711 379085
rect 523761 379051 523779 379085
rect 523833 379051 523847 379085
rect 523905 379051 523915 379085
rect 523977 379051 523983 379085
rect 524049 379051 524051 379085
rect 524085 379051 524087 379085
rect 524153 379051 524159 379085
rect 524221 379051 524231 379085
rect 524289 379051 524303 379085
rect 524357 379051 524375 379085
rect 524425 379051 524447 379085
rect 524493 379051 524519 379085
rect 524561 379051 524591 379085
rect 524629 379051 524663 379085
rect 524697 379051 524858 379085
rect 523338 378593 523439 378627
rect 523473 378593 523507 378627
rect 523545 378593 523575 378627
rect 523617 378593 523643 378627
rect 523689 378593 523711 378627
rect 523761 378593 523779 378627
rect 523833 378593 523847 378627
rect 523905 378593 523915 378627
rect 523977 378593 523983 378627
rect 524049 378593 524051 378627
rect 524085 378593 524087 378627
rect 524153 378593 524159 378627
rect 524221 378593 524231 378627
rect 524289 378593 524303 378627
rect 524357 378593 524375 378627
rect 524425 378593 524447 378627
rect 524493 378593 524519 378627
rect 524561 378593 524591 378627
rect 524629 378593 524663 378627
rect 524697 378593 524717 378627
rect 523158 378341 523218 378586
rect 523158 378307 523171 378341
rect 523205 378307 523218 378341
rect 523158 377941 523218 378307
rect 523158 377907 523171 377941
rect 523205 377907 523218 377941
rect 509998 377485 510011 377519
rect 510045 377485 510058 377519
rect 509998 377119 510058 377485
rect 509998 377085 510011 377119
rect 510045 377085 510058 377119
rect 509998 376719 510058 377085
rect 509998 376685 510011 376719
rect 510045 376685 510058 376719
rect 509998 376319 510058 376685
rect 509998 376285 510011 376319
rect 510045 376285 510058 376319
rect 509998 375919 510058 376285
rect 509998 375885 510011 375919
rect 510045 375885 510058 375919
rect 509998 375519 510058 375885
rect 509998 375485 510011 375519
rect 510045 375485 510058 375519
rect 509998 375119 510058 375485
rect 509998 375085 510011 375119
rect 510045 375085 510058 375119
rect 509998 374719 510058 375085
rect 509998 374685 510011 374719
rect 510045 374685 510058 374719
rect 509998 374319 510058 374685
rect 511878 377552 511938 377580
rect 511878 377539 512148 377552
rect 511878 377505 512031 377539
rect 512065 377505 512148 377539
rect 511878 377492 512148 377505
rect 511878 377299 511938 377492
rect 513518 377435 513578 377482
rect 511878 377265 511891 377299
rect 511925 377265 511938 377299
rect 511878 376899 511938 377265
rect 511878 376865 511891 376899
rect 511925 376865 511938 376899
rect 511878 376504 511938 376865
rect 512058 376977 512098 377422
rect 512139 377401 512159 377435
rect 512193 377401 512227 377435
rect 512265 377401 512295 377435
rect 512337 377401 512363 377435
rect 512409 377401 512431 377435
rect 512481 377401 512499 377435
rect 512553 377401 512567 377435
rect 512625 377401 512635 377435
rect 512697 377401 512703 377435
rect 512769 377401 512771 377435
rect 512805 377401 512807 377435
rect 512873 377401 512879 377435
rect 512941 377401 512951 377435
rect 513009 377401 513023 377435
rect 513077 377401 513095 377435
rect 513145 377401 513167 377435
rect 513213 377401 513239 377435
rect 513281 377401 513311 377435
rect 513349 377401 513383 377435
rect 513417 377401 513578 377435
rect 512058 376943 512159 376977
rect 512193 376943 512227 376977
rect 512265 376943 512295 376977
rect 512337 376943 512363 376977
rect 512409 376943 512431 376977
rect 512481 376943 512499 376977
rect 512553 376943 512567 376977
rect 512625 376943 512635 376977
rect 512697 376943 512703 376977
rect 512769 376943 512771 376977
rect 512805 376943 512807 376977
rect 512873 376943 512879 376977
rect 512941 376943 512951 376977
rect 513009 376943 513023 376977
rect 513077 376943 513095 376977
rect 513145 376943 513167 376977
rect 513213 376943 513239 376977
rect 513281 376943 513311 376977
rect 513349 376943 513383 376977
rect 513417 376943 513437 376977
rect 511878 376499 512018 376504
rect 511878 376465 511891 376499
rect 511925 376465 512018 376499
rect 511878 376439 512018 376465
rect 511878 376405 511981 376439
rect 512015 376405 512018 376439
rect 511878 376344 512018 376405
rect 511878 376099 511938 376344
rect 511878 376065 511891 376099
rect 511925 376065 511938 376099
rect 511878 375699 511938 376065
rect 511878 375665 511891 375699
rect 511925 375665 511938 375699
rect 511878 375299 511938 375665
rect 511878 375265 511891 375299
rect 511925 375265 511938 375299
rect 511878 374899 511938 375265
rect 511878 374865 511891 374899
rect 511925 374865 511938 374899
rect 511878 374606 511938 374865
rect 512058 376061 512098 376943
rect 513518 376519 513578 377401
rect 512139 376485 512159 376519
rect 512193 376485 512227 376519
rect 512265 376485 512295 376519
rect 512337 376485 512363 376519
rect 512409 376485 512431 376519
rect 512481 376485 512499 376519
rect 512553 376485 512567 376519
rect 512625 376485 512635 376519
rect 512697 376485 512703 376519
rect 512769 376485 512771 376519
rect 512805 376485 512807 376519
rect 512873 376485 512879 376519
rect 512941 376485 512951 376519
rect 513009 376485 513023 376519
rect 513077 376485 513095 376519
rect 513145 376485 513167 376519
rect 513213 376485 513239 376519
rect 513281 376485 513311 376519
rect 513349 376485 513383 376519
rect 513417 376485 513578 376519
rect 513518 376377 513578 376485
rect 513551 376343 513578 376377
rect 512058 376027 512159 376061
rect 512193 376027 512227 376061
rect 512265 376027 512295 376061
rect 512337 376027 512363 376061
rect 512409 376027 512431 376061
rect 512481 376027 512499 376061
rect 512553 376027 512567 376061
rect 512625 376027 512635 376061
rect 512697 376027 512703 376061
rect 512769 376027 512771 376061
rect 512805 376027 512807 376061
rect 512873 376027 512879 376061
rect 512941 376027 512951 376061
rect 513009 376027 513023 376061
rect 513077 376027 513095 376061
rect 513145 376027 513167 376061
rect 513213 376027 513239 376061
rect 513281 376027 513311 376061
rect 513349 376027 513383 376061
rect 513417 376027 513437 376061
rect 512058 375145 512098 376027
rect 513518 375603 513578 376343
rect 512139 375569 512159 375603
rect 512193 375569 512227 375603
rect 512265 375569 512295 375603
rect 512337 375569 512363 375603
rect 512409 375569 512431 375603
rect 512481 375569 512499 375603
rect 512553 375569 512567 375603
rect 512625 375569 512635 375603
rect 512697 375569 512703 375603
rect 512769 375569 512771 375603
rect 512805 375569 512807 375603
rect 512873 375569 512879 375603
rect 512941 375569 512951 375603
rect 513009 375569 513023 375603
rect 513077 375569 513095 375603
rect 513145 375569 513167 375603
rect 513213 375569 513239 375603
rect 513281 375569 513311 375603
rect 513349 375569 513383 375603
rect 513417 375569 513578 375603
rect 512058 375111 512159 375145
rect 512193 375111 512227 375145
rect 512265 375111 512295 375145
rect 512337 375111 512363 375145
rect 512409 375111 512431 375145
rect 512481 375111 512499 375145
rect 512553 375111 512567 375145
rect 512625 375111 512635 375145
rect 512697 375111 512703 375145
rect 512769 375111 512771 375145
rect 512805 375111 512807 375145
rect 512873 375111 512879 375145
rect 512941 375111 512951 375145
rect 513009 375111 513023 375145
rect 513077 375111 513095 375145
rect 513145 375111 513167 375145
rect 513213 375111 513239 375145
rect 513281 375111 513311 375145
rect 513349 375111 513383 375145
rect 513417 375111 513437 375145
rect 512058 374629 512098 375111
rect 513518 374687 513578 375569
rect 512139 374653 512159 374687
rect 512193 374653 512227 374687
rect 512265 374653 512295 374687
rect 512337 374653 512363 374687
rect 512409 374653 512431 374687
rect 512481 374653 512499 374687
rect 512553 374653 512567 374687
rect 512625 374653 512635 374687
rect 512697 374653 512703 374687
rect 512769 374653 512771 374687
rect 512805 374653 512807 374687
rect 512873 374653 512879 374687
rect 512941 374653 512951 374687
rect 513009 374653 513023 374687
rect 513077 374653 513095 374687
rect 513145 374653 513167 374687
rect 513213 374653 513239 374687
rect 513281 374653 513311 374687
rect 513349 374653 513383 374687
rect 513417 374653 513578 374687
rect 512058 374606 512061 374629
rect 512095 374606 512098 374629
rect 513518 374606 513578 374653
rect 513624 377299 513684 377482
rect 513624 377265 513637 377299
rect 513671 377265 513684 377299
rect 513624 376899 513684 377265
rect 513624 376865 513637 376899
rect 513671 376865 513684 376899
rect 513624 376499 513684 376865
rect 513624 376465 513637 376499
rect 513671 376465 513684 376499
rect 513624 376377 513684 376465
rect 513758 377299 513818 377580
rect 513758 377265 513771 377299
rect 513805 377265 513818 377299
rect 513758 376899 513818 377265
rect 513758 376865 513771 376899
rect 513805 376865 513818 376899
rect 513758 376499 513818 376865
rect 513758 376465 513771 376499
rect 513805 376465 513818 376499
rect 513624 376343 513653 376377
rect 513624 376099 513684 376343
rect 513624 376065 513637 376099
rect 513671 376065 513684 376099
rect 513624 375699 513684 376065
rect 513624 375665 513637 375699
rect 513671 375665 513684 375699
rect 513624 375299 513684 375665
rect 513624 375265 513637 375299
rect 513671 375265 513684 375299
rect 513624 374899 513684 375265
rect 513624 374865 513637 374899
rect 513671 374865 513684 374899
rect 513624 374606 513684 374865
rect 513758 376099 513818 376465
rect 513758 376065 513771 376099
rect 513805 376065 513818 376099
rect 513758 375699 513818 376065
rect 513758 375665 513771 375699
rect 513805 375665 513818 375699
rect 513758 375299 513818 375665
rect 513758 375265 513771 375299
rect 513805 375265 513818 375299
rect 513758 374899 513818 375265
rect 515638 377377 515698 377560
rect 515638 377343 515651 377377
rect 515685 377343 515698 377377
rect 515638 377177 515698 377343
rect 515638 377143 515651 377177
rect 515685 377143 515698 377177
rect 515638 376977 515698 377143
rect 517518 377377 517578 377560
rect 517518 377343 517531 377377
rect 517565 377343 517578 377377
rect 517518 377177 517578 377343
rect 517518 377143 517531 377177
rect 517565 377143 517578 377177
rect 515638 376943 515651 376977
rect 515685 376943 515698 376977
rect 515638 376777 515698 376943
rect 515638 376743 515651 376777
rect 515685 376743 515698 376777
rect 515638 376577 515698 376743
rect 517518 376977 517578 377143
rect 517518 376943 517531 376977
rect 517565 376943 517578 376977
rect 517518 376777 517578 376943
rect 517518 376743 517531 376777
rect 517565 376743 517578 376777
rect 517518 376648 517578 376743
rect 515638 376543 515651 376577
rect 515685 376543 515698 376577
rect 515638 376377 515698 376543
rect 515638 376343 515651 376377
rect 515685 376343 515698 376377
rect 515638 376177 515698 376343
rect 515638 376143 515651 376177
rect 515685 376143 515698 376177
rect 515638 375977 515698 376143
rect 516578 376577 517578 376648
rect 516578 376561 517531 376577
rect 516578 376119 516617 376561
rect 516719 376543 517531 376561
rect 517565 376543 517578 376577
rect 516719 376377 517578 376543
rect 516719 376343 517531 376377
rect 517565 376343 517578 376377
rect 516719 376177 517578 376343
rect 516719 376143 517531 376177
rect 517565 376143 517578 376177
rect 516719 376119 517578 376143
rect 516578 376032 517578 376119
rect 515638 375943 515651 375977
rect 515685 375943 515698 375977
rect 515638 375777 515698 375943
rect 515638 375743 515651 375777
rect 515685 375743 515698 375777
rect 515638 375577 515698 375743
rect 515638 375543 515651 375577
rect 515685 375543 515698 375577
rect 517518 375977 517578 376032
rect 517518 375943 517531 375977
rect 517565 375943 517578 375977
rect 517518 375777 517578 375943
rect 517518 375743 517531 375777
rect 517565 375743 517578 375777
rect 517518 375577 517578 375743
rect 515638 375377 515698 375543
rect 515638 375343 515651 375377
rect 515685 375343 515698 375377
rect 515638 375120 515698 375343
rect 516473 375120 516863 375552
rect 517518 375543 517531 375577
rect 517565 375543 517578 375577
rect 517518 375377 517578 375543
rect 517518 375343 517531 375377
rect 517565 375343 517578 375377
rect 517518 375120 517578 375343
rect 519398 377377 519458 377560
rect 519398 377343 519411 377377
rect 519445 377343 519458 377377
rect 519398 377177 519458 377343
rect 519398 377143 519411 377177
rect 519445 377143 519458 377177
rect 519398 376977 519458 377143
rect 521278 377377 521338 377560
rect 521278 377343 521291 377377
rect 521325 377343 521338 377377
rect 521278 377177 521338 377343
rect 521278 377143 521291 377177
rect 521325 377143 521338 377177
rect 519398 376943 519411 376977
rect 519445 376943 519458 376977
rect 519398 376777 519458 376943
rect 519398 376743 519411 376777
rect 519445 376743 519458 376777
rect 519398 376577 519458 376743
rect 521278 376977 521338 377143
rect 521278 376943 521291 376977
rect 521325 376943 521338 376977
rect 521278 376777 521338 376943
rect 521278 376743 521291 376777
rect 521325 376743 521338 376777
rect 521278 376648 521338 376743
rect 519398 376543 519411 376577
rect 519445 376543 519458 376577
rect 519398 376377 519458 376543
rect 519398 376343 519411 376377
rect 519445 376343 519458 376377
rect 519398 376177 519458 376343
rect 519398 376143 519411 376177
rect 519445 376143 519458 376177
rect 519398 375977 519458 376143
rect 520338 376577 521338 376648
rect 520338 376561 521291 376577
rect 520338 376119 520377 376561
rect 520479 376543 521291 376561
rect 521325 376543 521338 376577
rect 520479 376377 521338 376543
rect 520479 376343 521291 376377
rect 521325 376343 521338 376377
rect 520479 376177 521338 376343
rect 520479 376143 521291 376177
rect 521325 376143 521338 376177
rect 520479 376119 521338 376143
rect 520338 376032 521338 376119
rect 519398 375943 519411 375977
rect 519445 375943 519458 375977
rect 519398 375777 519458 375943
rect 519398 375743 519411 375777
rect 519445 375743 519458 375777
rect 519398 375577 519458 375743
rect 519398 375543 519411 375577
rect 519445 375543 519458 375577
rect 521278 375977 521338 376032
rect 521278 375943 521291 375977
rect 521325 375943 521338 375977
rect 521278 375777 521338 375943
rect 521278 375743 521291 375777
rect 521325 375743 521338 375777
rect 521278 375577 521338 375743
rect 519398 375377 519458 375543
rect 519398 375343 519411 375377
rect 519445 375343 519458 375377
rect 519398 375120 519458 375343
rect 520233 375120 520623 375552
rect 521278 375543 521291 375577
rect 521325 375543 521338 375577
rect 521278 375377 521338 375543
rect 521278 375343 521291 375377
rect 521325 375343 521338 375377
rect 521278 375120 521338 375343
rect 523158 377541 523218 377907
rect 523158 377507 523171 377541
rect 523205 377507 523218 377541
rect 523158 377446 523218 377507
rect 523338 377711 523378 378593
rect 524798 378169 524858 379051
rect 523419 378135 523439 378169
rect 523473 378135 523507 378169
rect 523545 378135 523575 378169
rect 523617 378135 523643 378169
rect 523689 378135 523711 378169
rect 523761 378135 523779 378169
rect 523833 378135 523847 378169
rect 523905 378135 523915 378169
rect 523977 378135 523983 378169
rect 524049 378135 524051 378169
rect 524085 378135 524087 378169
rect 524153 378135 524159 378169
rect 524221 378135 524231 378169
rect 524289 378135 524303 378169
rect 524357 378135 524375 378169
rect 524425 378135 524447 378169
rect 524493 378135 524519 378169
rect 524561 378135 524591 378169
rect 524629 378135 524663 378169
rect 524697 378135 524858 378169
rect 523338 377677 523439 377711
rect 523473 377677 523507 377711
rect 523545 377677 523575 377711
rect 523617 377677 523643 377711
rect 523689 377677 523711 377711
rect 523761 377677 523779 377711
rect 523833 377677 523847 377711
rect 523905 377677 523915 377711
rect 523977 377677 523983 377711
rect 524049 377677 524051 377711
rect 524085 377677 524087 377711
rect 524153 377677 524159 377711
rect 524221 377677 524231 377711
rect 524289 377677 524303 377711
rect 524357 377677 524375 377711
rect 524425 377677 524447 377711
rect 524493 377677 524519 377711
rect 524561 377677 524591 377711
rect 524629 377677 524663 377711
rect 524697 377677 524717 377711
rect 523158 377381 523298 377446
rect 523158 377347 523261 377381
rect 523295 377347 523298 377381
rect 523158 377286 523298 377347
rect 523158 377141 523218 377286
rect 523158 377107 523171 377141
rect 523205 377107 523218 377141
rect 523158 376741 523218 377107
rect 523158 376707 523171 376741
rect 523205 376707 523218 376741
rect 523158 376341 523218 376707
rect 523158 376307 523171 376341
rect 523205 376307 523218 376341
rect 523158 376146 523218 376307
rect 523338 376795 523378 377677
rect 524798 377253 524858 378135
rect 523419 377219 523439 377253
rect 523473 377219 523507 377253
rect 523545 377219 523575 377253
rect 523617 377219 523643 377253
rect 523689 377219 523711 377253
rect 523761 377219 523779 377253
rect 523833 377219 523847 377253
rect 523905 377219 523915 377253
rect 523977 377219 523983 377253
rect 524049 377219 524051 377253
rect 524085 377219 524087 377253
rect 524153 377219 524159 377253
rect 524221 377219 524231 377253
rect 524289 377219 524303 377253
rect 524357 377219 524375 377253
rect 524425 377219 524447 377253
rect 524493 377219 524519 377253
rect 524561 377219 524591 377253
rect 524629 377219 524663 377253
rect 524697 377219 524858 377253
rect 523338 376761 523439 376795
rect 523473 376761 523507 376795
rect 523545 376761 523575 376795
rect 523617 376761 523643 376795
rect 523689 376761 523711 376795
rect 523761 376761 523779 376795
rect 523833 376761 523847 376795
rect 523905 376761 523915 376795
rect 523977 376761 523983 376795
rect 524049 376761 524051 376795
rect 524085 376761 524087 376795
rect 524153 376761 524159 376795
rect 524221 376761 524231 376795
rect 524289 376761 524303 376795
rect 524357 376761 524375 376795
rect 524425 376761 524447 376795
rect 524493 376761 524519 376795
rect 524561 376761 524591 376795
rect 524629 376761 524663 376795
rect 524697 376761 524717 376795
rect 523158 376081 523298 376146
rect 523158 376047 523261 376081
rect 523295 376047 523298 376081
rect 523158 375986 523298 376047
rect 523158 375941 523218 375986
rect 523158 375907 523171 375941
rect 523205 375907 523218 375941
rect 523158 375541 523218 375907
rect 523158 375507 523171 375541
rect 523205 375507 523218 375541
rect 523158 375141 523218 375507
rect 513758 374865 513771 374899
rect 513805 374865 513818 374899
rect 513758 374606 513818 374865
rect 523158 375107 523171 375141
rect 523205 375107 523218 375141
rect 523158 374846 523218 375107
rect 523338 375879 523378 376761
rect 524798 376337 524858 377219
rect 523419 376303 523439 376337
rect 523473 376303 523507 376337
rect 523545 376303 523575 376337
rect 523617 376303 523643 376337
rect 523689 376303 523711 376337
rect 523761 376303 523779 376337
rect 523833 376303 523847 376337
rect 523905 376303 523915 376337
rect 523977 376303 523983 376337
rect 524049 376303 524051 376337
rect 524085 376303 524087 376337
rect 524153 376303 524159 376337
rect 524221 376303 524231 376337
rect 524289 376303 524303 376337
rect 524357 376303 524375 376337
rect 524425 376303 524447 376337
rect 524493 376303 524519 376337
rect 524561 376303 524591 376337
rect 524629 376303 524663 376337
rect 524697 376303 524858 376337
rect 523338 375845 523439 375879
rect 523473 375845 523507 375879
rect 523545 375845 523575 375879
rect 523617 375845 523643 375879
rect 523689 375845 523711 375879
rect 523761 375845 523779 375879
rect 523833 375845 523847 375879
rect 523905 375845 523915 375879
rect 523977 375845 523983 375879
rect 524049 375845 524051 375879
rect 524085 375845 524087 375879
rect 524153 375845 524159 375879
rect 524221 375845 524231 375879
rect 524289 375845 524303 375879
rect 524357 375845 524375 375879
rect 524425 375845 524447 375879
rect 524493 375845 524519 375879
rect 524561 375845 524591 375879
rect 524629 375845 524663 375879
rect 524697 375845 524717 375879
rect 523338 374963 523378 375845
rect 524798 375421 524858 376303
rect 523419 375387 523439 375421
rect 523473 375387 523507 375421
rect 523545 375387 523575 375421
rect 523617 375387 523643 375421
rect 523689 375387 523711 375421
rect 523761 375387 523779 375421
rect 523833 375387 523847 375421
rect 523905 375387 523915 375421
rect 523977 375387 523983 375421
rect 524049 375387 524051 375421
rect 524085 375387 524087 375421
rect 524153 375387 524159 375421
rect 524221 375387 524231 375421
rect 524289 375387 524303 375421
rect 524357 375387 524375 375421
rect 524425 375387 524447 375421
rect 524493 375387 524519 375421
rect 524561 375387 524591 375421
rect 524629 375387 524663 375421
rect 524697 375387 524858 375421
rect 523338 374929 523439 374963
rect 523473 374929 523507 374963
rect 523545 374929 523575 374963
rect 523617 374929 523643 374963
rect 523689 374929 523711 374963
rect 523761 374929 523779 374963
rect 523833 374929 523847 374963
rect 523905 374929 523915 374963
rect 523977 374929 523983 374963
rect 524049 374929 524051 374963
rect 524085 374929 524087 374963
rect 524153 374929 524159 374963
rect 524221 374929 524231 374963
rect 524289 374929 524303 374963
rect 524357 374929 524375 374963
rect 524425 374929 524447 374963
rect 524493 374929 524519 374963
rect 524561 374929 524591 374963
rect 524629 374929 524663 374963
rect 524697 374929 524717 374963
rect 515638 374633 515698 374816
rect 515638 374599 515651 374633
rect 515685 374599 515698 374633
rect 509998 374285 510011 374319
rect 510045 374285 510058 374319
rect 509998 374134 510058 374285
rect 515638 374433 515698 374599
rect 515638 374399 515651 374433
rect 515685 374399 515698 374433
rect 515638 374233 515698 374399
rect 517518 374633 517578 374816
rect 517518 374599 517531 374633
rect 517565 374599 517578 374633
rect 517518 374433 517578 374599
rect 517518 374399 517531 374433
rect 517565 374399 517578 374433
rect 515638 374199 515651 374233
rect 515685 374199 515698 374233
rect 502478 373861 502491 373895
rect 502525 373861 502538 373895
rect 502478 373498 502538 373861
rect 515638 374033 515698 374199
rect 515638 373999 515651 374033
rect 515685 373999 515698 374033
rect 515638 373833 515698 373999
rect 517518 374233 517578 374399
rect 517518 374199 517531 374233
rect 517565 374199 517578 374233
rect 517518 374033 517578 374199
rect 517518 373999 517531 374033
rect 517565 373999 517578 374033
rect 517518 373904 517578 373999
rect 515638 373799 515651 373833
rect 515685 373799 515698 373833
rect 515638 373633 515698 373799
rect 515638 373599 515651 373633
rect 515685 373599 515698 373633
rect 498718 373307 498731 373341
rect 498765 373307 498778 373341
rect 498718 372941 498778 373307
rect 515638 373433 515698 373599
rect 515638 373399 515651 373433
rect 515685 373399 515698 373433
rect 515638 373233 515698 373399
rect 516578 373833 517578 373904
rect 516578 373817 517531 373833
rect 516578 373375 516617 373817
rect 516719 373799 517531 373817
rect 517565 373799 517578 373833
rect 516719 373633 517578 373799
rect 516719 373599 517531 373633
rect 517565 373599 517578 373633
rect 516719 373433 517578 373599
rect 516719 373399 517531 373433
rect 517565 373399 517578 373433
rect 516719 373375 517578 373399
rect 516578 373288 517578 373375
rect 515638 373199 515651 373233
rect 515685 373199 515698 373233
rect 498718 372907 498731 372941
rect 498765 372907 498778 372941
rect 498718 372541 498778 372907
rect 498718 372507 498731 372541
rect 498765 372507 498778 372541
rect 498718 372316 498778 372507
rect 500598 372987 500658 373170
rect 500598 372953 500611 372987
rect 500645 372953 500658 372987
rect 500598 372787 500658 372953
rect 500598 372753 500611 372787
rect 500645 372753 500658 372787
rect 500598 372587 500658 372753
rect 500598 372553 500611 372587
rect 500645 372553 500658 372587
rect 500598 372387 500658 372553
rect 500598 372353 500611 372387
rect 500645 372353 500658 372387
rect 494958 371941 495018 372307
rect 500598 372187 500658 372353
rect 500598 372153 500611 372187
rect 500645 372153 500658 372187
rect 494958 371907 494971 371941
rect 495005 371907 495018 371941
rect 494958 371541 495018 371907
rect 494958 371507 494971 371541
rect 495005 371507 495018 371541
rect 494958 371141 495018 371507
rect 494958 371107 494971 371141
rect 495005 371107 495018 371141
rect 494958 370741 495018 371107
rect 494958 370707 494971 370741
rect 495005 370707 495018 370741
rect 494958 370341 495018 370707
rect 494958 370307 494971 370341
rect 495005 370307 495018 370341
rect 494958 369941 495018 370307
rect 494958 369907 494971 369941
rect 495005 369907 495018 369941
rect 494958 369541 495018 369907
rect 494958 369507 494971 369541
rect 495005 369507 495018 369541
rect 494958 369141 495018 369507
rect 494958 369107 494971 369141
rect 495005 369107 495018 369141
rect 494958 368741 495018 369107
rect 494958 368707 494971 368741
rect 495005 368707 495018 368741
rect 494958 368341 495018 368707
rect 494958 368307 494971 368341
rect 495005 368307 495018 368341
rect 494958 367941 495018 368307
rect 494958 367907 494971 367941
rect 495005 367907 495018 367941
rect 494958 367541 495018 367907
rect 494958 367507 494971 367541
rect 495005 367507 495018 367541
rect 494958 367141 495018 367507
rect 494958 367107 494971 367141
rect 495005 367107 495018 367141
rect 494958 366741 495018 367107
rect 494958 366707 494971 366741
rect 495005 366707 495018 366741
rect 494958 366341 495018 366707
rect 494958 366307 494971 366341
rect 495005 366307 495018 366341
rect 494958 365941 495018 366307
rect 494958 365907 494971 365941
rect 495005 365907 495018 365941
rect 494958 365541 495018 365907
rect 494958 365507 494971 365541
rect 495005 365507 495018 365541
rect 494958 365141 495018 365507
rect 494958 365107 494971 365141
rect 495005 365107 495018 365141
rect 494958 364741 495018 365107
rect 494958 364707 494971 364741
rect 495005 364707 495018 364741
rect 494958 364341 495018 364707
rect 494958 364307 494971 364341
rect 495005 364307 495018 364341
rect 494958 363941 495018 364307
rect 494958 363907 494971 363941
rect 495005 363907 495018 363941
rect 494958 363541 495018 363907
rect 494958 363507 494971 363541
rect 495005 363507 495018 363541
rect 494958 363141 495018 363507
rect 494958 363107 494971 363141
rect 495005 363107 495018 363141
rect 494958 362741 495018 363107
rect 494958 362707 494971 362741
rect 495005 362707 495018 362741
rect 494958 362516 495018 362707
rect 496838 371811 496898 371994
rect 496838 371777 496851 371811
rect 496885 371777 496898 371811
rect 496838 371611 496898 371777
rect 496838 371577 496851 371611
rect 496885 371577 496898 371611
rect 496838 371411 496898 371577
rect 496838 371377 496851 371411
rect 496885 371377 496898 371411
rect 496838 371211 496898 371377
rect 496838 371177 496851 371211
rect 496885 371177 496898 371211
rect 496838 371011 496898 371177
rect 496838 370977 496851 371011
rect 496885 370977 496898 371011
rect 496838 370811 496898 370977
rect 496838 370777 496851 370811
rect 496885 370777 496898 370811
rect 496838 370611 496898 370777
rect 496838 370577 496851 370611
rect 496885 370577 496898 370611
rect 496838 370411 496898 370577
rect 496838 370377 496851 370411
rect 496885 370377 496898 370411
rect 496838 370211 496898 370377
rect 496838 370177 496851 370211
rect 496885 370177 496898 370211
rect 496838 370011 496898 370177
rect 496838 369977 496851 370011
rect 496885 369977 496898 370011
rect 496838 369811 496898 369977
rect 496838 369777 496851 369811
rect 496885 369777 496898 369811
rect 496838 369611 496898 369777
rect 496838 369577 496851 369611
rect 496885 369577 496898 369611
rect 496838 369411 496898 369577
rect 496838 369377 496851 369411
rect 496885 369377 496898 369411
rect 496838 369211 496898 369377
rect 496838 369177 496851 369211
rect 496885 369177 496898 369211
rect 496838 369011 496898 369177
rect 496838 368977 496851 369011
rect 496885 368977 496898 369011
rect 496838 368811 496898 368977
rect 496838 368777 496851 368811
rect 496885 368777 496898 368811
rect 496838 368611 496898 368777
rect 496838 368577 496851 368611
rect 496885 368577 496898 368611
rect 496838 368411 496898 368577
rect 496838 368377 496851 368411
rect 496885 368377 496898 368411
rect 496838 368211 496898 368377
rect 496838 368177 496851 368211
rect 496885 368177 496898 368211
rect 496838 368011 496898 368177
rect 496838 367977 496851 368011
rect 496885 367977 496898 368011
rect 496838 367811 496898 367977
rect 496838 367777 496851 367811
rect 496885 367777 496898 367811
rect 496838 367611 496898 367777
rect 496838 367577 496851 367611
rect 496885 367577 496898 367611
rect 496838 367411 496898 367577
rect 496838 367377 496851 367411
rect 496885 367377 496898 367411
rect 496838 367211 496898 367377
rect 496838 367177 496851 367211
rect 496885 367177 496898 367211
rect 496838 367011 496898 367177
rect 496838 366977 496851 367011
rect 496885 366977 496898 367011
rect 496838 366811 496898 366977
rect 496838 366777 496851 366811
rect 496885 366777 496898 366811
rect 496838 366611 496898 366777
rect 496838 366577 496851 366611
rect 496885 366577 496898 366611
rect 496838 366411 496898 366577
rect 496838 366377 496851 366411
rect 496885 366377 496898 366411
rect 496838 366211 496898 366377
rect 496838 366177 496851 366211
rect 496885 366177 496898 366211
rect 496838 366011 496898 366177
rect 496838 365977 496851 366011
rect 496885 365977 496898 366011
rect 496838 365811 496898 365977
rect 496838 365777 496851 365811
rect 496885 365777 496898 365811
rect 496838 365611 496898 365777
rect 496838 365577 496851 365611
rect 496885 365577 496898 365611
rect 496838 365411 496898 365577
rect 496838 365377 496851 365411
rect 496885 365377 496898 365411
rect 496838 365211 496898 365377
rect 496838 365177 496851 365211
rect 496885 365177 496898 365211
rect 496838 365011 496898 365177
rect 496838 364977 496851 365011
rect 496885 364977 496898 365011
rect 496838 364811 496898 364977
rect 496838 364777 496851 364811
rect 496885 364777 496898 364811
rect 496838 364611 496898 364777
rect 496838 364577 496851 364611
rect 496885 364577 496898 364611
rect 496838 364411 496898 364577
rect 496838 364377 496851 364411
rect 496885 364377 496898 364411
rect 496838 364211 496898 364377
rect 496838 364177 496851 364211
rect 496885 364177 496898 364211
rect 496838 364011 496898 364177
rect 496838 363977 496851 364011
rect 496885 363977 496898 364011
rect 496838 363811 496898 363977
rect 496838 363777 496851 363811
rect 496885 363777 496898 363811
rect 496838 363611 496898 363777
rect 496838 363577 496851 363611
rect 496885 363577 496898 363611
rect 496838 363411 496898 363577
rect 496838 363377 496851 363411
rect 496885 363377 496898 363411
rect 496838 363211 496898 363377
rect 496838 363177 496851 363211
rect 496885 363177 496898 363211
rect 496838 363011 496898 363177
rect 496838 362977 496851 363011
rect 496885 362977 496898 363011
rect 496838 362811 496898 362977
rect 496838 362777 496851 362811
rect 496885 362777 496898 362811
rect 496838 362614 496898 362777
rect 497164 371948 498452 371968
rect 497164 371914 497184 371948
rect 497218 371934 498452 371948
rect 497218 371914 497222 371934
rect 497164 371900 497222 371914
rect 497256 371900 497312 371934
rect 497346 371900 497402 371934
rect 497436 371900 497492 371934
rect 497526 371900 497582 371934
rect 497616 371900 497672 371934
rect 497706 371900 497762 371934
rect 497796 371900 497852 371934
rect 497886 371900 497942 371934
rect 497976 371900 498032 371934
rect 498066 371900 498122 371934
rect 498156 371900 498212 371934
rect 498246 371900 498302 371934
rect 498336 371900 498452 371934
rect 497164 371869 498452 371900
rect 497164 371858 497263 371869
rect 497164 371824 497184 371858
rect 497218 371838 497263 371858
rect 497164 371804 497199 371824
rect 497233 371804 497263 371838
rect 498353 371838 498452 371869
rect 497164 371768 497263 371804
rect 497164 371734 497184 371768
rect 497218 371748 497263 371768
rect 497164 371714 497199 371734
rect 497233 371714 497263 371748
rect 497164 371678 497263 371714
rect 497164 371644 497184 371678
rect 497218 371658 497263 371678
rect 497164 371624 497199 371644
rect 497233 371624 497263 371658
rect 497164 371588 497263 371624
rect 497164 371554 497184 371588
rect 497218 371568 497263 371588
rect 497164 371534 497199 371554
rect 497233 371534 497263 371568
rect 497164 371498 497263 371534
rect 497164 371464 497184 371498
rect 497218 371478 497263 371498
rect 497164 371444 497199 371464
rect 497233 371444 497263 371478
rect 497164 371408 497263 371444
rect 497164 371374 497184 371408
rect 497218 371388 497263 371408
rect 497164 371354 497199 371374
rect 497233 371354 497263 371388
rect 497164 371318 497263 371354
rect 497164 371284 497184 371318
rect 497218 371298 497263 371318
rect 497164 371264 497199 371284
rect 497233 371264 497263 371298
rect 497164 371228 497263 371264
rect 497164 371194 497184 371228
rect 497218 371208 497263 371228
rect 497164 371174 497199 371194
rect 497233 371174 497263 371208
rect 497164 371138 497263 371174
rect 497164 371104 497184 371138
rect 497218 371118 497263 371138
rect 497164 371084 497199 371104
rect 497233 371084 497263 371118
rect 497164 371048 497263 371084
rect 497164 371014 497184 371048
rect 497218 371028 497263 371048
rect 497164 370994 497199 371014
rect 497233 370994 497263 371028
rect 497164 370958 497263 370994
rect 497164 370924 497184 370958
rect 497218 370938 497263 370958
rect 497164 370904 497199 370924
rect 497233 370904 497263 370938
rect 497164 370868 497263 370904
rect 497164 370834 497184 370868
rect 497218 370848 497263 370868
rect 497164 370814 497199 370834
rect 497233 370814 497263 370848
rect 497327 371786 498289 371805
rect 497327 371784 497403 371786
rect 497327 371750 497344 371784
rect 497378 371752 497403 371784
rect 497437 371752 497493 371786
rect 497527 371752 497583 371786
rect 497617 371752 497673 371786
rect 497707 371752 497763 371786
rect 497797 371752 497853 371786
rect 497887 371752 497943 371786
rect 497977 371752 498033 371786
rect 498067 371752 498123 371786
rect 498157 371752 498289 371786
rect 497378 371750 498289 371752
rect 497327 371733 498289 371750
rect 497327 371694 497399 371733
rect 497327 371660 497344 371694
rect 497378 371674 497399 371694
rect 497327 371640 497346 371660
rect 497380 371640 497399 371674
rect 498217 371708 498289 371733
rect 498217 371674 498236 371708
rect 498270 371674 498289 371708
rect 497327 371604 497399 371640
rect 497327 371570 497344 371604
rect 497378 371584 497399 371604
rect 497327 371550 497346 371570
rect 497380 371550 497399 371584
rect 497327 371514 497399 371550
rect 497327 371480 497344 371514
rect 497378 371494 497399 371514
rect 497327 371460 497346 371480
rect 497380 371460 497399 371494
rect 497327 371424 497399 371460
rect 497327 371390 497344 371424
rect 497378 371404 497399 371424
rect 497327 371370 497346 371390
rect 497380 371370 497399 371404
rect 497327 371334 497399 371370
rect 497327 371300 497344 371334
rect 497378 371314 497399 371334
rect 497327 371280 497346 371300
rect 497380 371280 497399 371314
rect 497327 371244 497399 371280
rect 497327 371210 497344 371244
rect 497378 371224 497399 371244
rect 497327 371190 497346 371210
rect 497380 371190 497399 371224
rect 497327 371154 497399 371190
rect 497327 371120 497344 371154
rect 497378 371134 497399 371154
rect 497327 371100 497346 371120
rect 497380 371100 497399 371134
rect 497327 371064 497399 371100
rect 497327 371030 497344 371064
rect 497378 371044 497399 371064
rect 497327 371010 497346 371030
rect 497380 371010 497399 371044
rect 497327 370974 497399 371010
rect 497461 371610 498155 371671
rect 497461 371576 497520 371610
rect 497554 371598 497610 371610
rect 497582 371576 497610 371598
rect 497644 371598 497700 371610
rect 497644 371576 497648 371598
rect 497461 371564 497548 371576
rect 497582 371564 497648 371576
rect 497682 371576 497700 371598
rect 497734 371598 497790 371610
rect 497734 371576 497748 371598
rect 497682 371564 497748 371576
rect 497782 371576 497790 371598
rect 497824 371598 497880 371610
rect 497914 371598 497970 371610
rect 498004 371598 498060 371610
rect 497824 371576 497848 371598
rect 497914 371576 497948 371598
rect 498004 371576 498048 371598
rect 498094 371576 498155 371610
rect 497782 371564 497848 371576
rect 497882 371564 497948 371576
rect 497982 371564 498048 371576
rect 498082 371564 498155 371576
rect 497461 371520 498155 371564
rect 497461 371486 497520 371520
rect 497554 371498 497610 371520
rect 497582 371486 497610 371498
rect 497644 371498 497700 371520
rect 497644 371486 497648 371498
rect 497461 371464 497548 371486
rect 497582 371464 497648 371486
rect 497682 371486 497700 371498
rect 497734 371498 497790 371520
rect 497734 371486 497748 371498
rect 497682 371464 497748 371486
rect 497782 371486 497790 371498
rect 497824 371498 497880 371520
rect 497914 371498 497970 371520
rect 498004 371498 498060 371520
rect 497824 371486 497848 371498
rect 497914 371486 497948 371498
rect 498004 371486 498048 371498
rect 498094 371486 498155 371520
rect 497782 371464 497848 371486
rect 497882 371464 497948 371486
rect 497982 371464 498048 371486
rect 498082 371464 498155 371486
rect 497461 371430 498155 371464
rect 497461 371396 497520 371430
rect 497554 371398 497610 371430
rect 497582 371396 497610 371398
rect 497644 371398 497700 371430
rect 497644 371396 497648 371398
rect 497461 371364 497548 371396
rect 497582 371364 497648 371396
rect 497682 371396 497700 371398
rect 497734 371398 497790 371430
rect 497734 371396 497748 371398
rect 497682 371364 497748 371396
rect 497782 371396 497790 371398
rect 497824 371398 497880 371430
rect 497914 371398 497970 371430
rect 498004 371398 498060 371430
rect 497824 371396 497848 371398
rect 497914 371396 497948 371398
rect 498004 371396 498048 371398
rect 498094 371396 498155 371430
rect 497782 371364 497848 371396
rect 497882 371364 497948 371396
rect 497982 371364 498048 371396
rect 498082 371364 498155 371396
rect 497461 371340 498155 371364
rect 497461 371306 497520 371340
rect 497554 371306 497610 371340
rect 497644 371306 497700 371340
rect 497734 371306 497790 371340
rect 497824 371306 497880 371340
rect 497914 371306 497970 371340
rect 498004 371306 498060 371340
rect 498094 371306 498155 371340
rect 497461 371298 498155 371306
rect 497461 371264 497548 371298
rect 497582 371264 497648 371298
rect 497682 371264 497748 371298
rect 497782 371264 497848 371298
rect 497882 371264 497948 371298
rect 497982 371264 498048 371298
rect 498082 371264 498155 371298
rect 497461 371250 498155 371264
rect 497461 371216 497520 371250
rect 497554 371216 497610 371250
rect 497644 371216 497700 371250
rect 497734 371216 497790 371250
rect 497824 371216 497880 371250
rect 497914 371216 497970 371250
rect 498004 371216 498060 371250
rect 498094 371216 498155 371250
rect 497461 371198 498155 371216
rect 497461 371164 497548 371198
rect 497582 371164 497648 371198
rect 497682 371164 497748 371198
rect 497782 371164 497848 371198
rect 497882 371164 497948 371198
rect 497982 371164 498048 371198
rect 498082 371164 498155 371198
rect 497461 371160 498155 371164
rect 497461 371126 497520 371160
rect 497554 371126 497610 371160
rect 497644 371126 497700 371160
rect 497734 371126 497790 371160
rect 497824 371126 497880 371160
rect 497914 371126 497970 371160
rect 498004 371126 498060 371160
rect 498094 371126 498155 371160
rect 497461 371098 498155 371126
rect 497461 371070 497548 371098
rect 497582 371070 497648 371098
rect 497461 371036 497520 371070
rect 497582 371064 497610 371070
rect 497554 371036 497610 371064
rect 497644 371064 497648 371070
rect 497682 371070 497748 371098
rect 497682 371064 497700 371070
rect 497644 371036 497700 371064
rect 497734 371064 497748 371070
rect 497782 371070 497848 371098
rect 497882 371070 497948 371098
rect 497982 371070 498048 371098
rect 498082 371070 498155 371098
rect 497782 371064 497790 371070
rect 497734 371036 497790 371064
rect 497824 371064 497848 371070
rect 497914 371064 497948 371070
rect 498004 371064 498048 371070
rect 497824 371036 497880 371064
rect 497914 371036 497970 371064
rect 498004 371036 498060 371064
rect 498094 371036 498155 371070
rect 497461 370977 498155 371036
rect 498217 371618 498289 371674
rect 498217 371584 498236 371618
rect 498270 371584 498289 371618
rect 498217 371528 498289 371584
rect 498217 371494 498236 371528
rect 498270 371494 498289 371528
rect 498217 371438 498289 371494
rect 498217 371404 498236 371438
rect 498270 371404 498289 371438
rect 498217 371348 498289 371404
rect 498217 371314 498236 371348
rect 498270 371314 498289 371348
rect 498217 371258 498289 371314
rect 498217 371224 498236 371258
rect 498270 371224 498289 371258
rect 498217 371168 498289 371224
rect 498217 371134 498236 371168
rect 498270 371134 498289 371168
rect 498217 371078 498289 371134
rect 498217 371044 498236 371078
rect 498270 371044 498289 371078
rect 498217 370988 498289 371044
rect 497327 370940 497344 370974
rect 497378 370954 497399 370974
rect 497327 370920 497346 370940
rect 497380 370920 497399 370954
rect 497327 370915 497399 370920
rect 498217 370954 498236 370988
rect 498270 370954 498289 370988
rect 498217 370915 498289 370954
rect 497327 370896 498289 370915
rect 497327 370884 497422 370896
rect 497327 370850 497344 370884
rect 497378 370862 497422 370884
rect 497456 370862 497512 370896
rect 497546 370862 497602 370896
rect 497636 370862 497692 370896
rect 497726 370862 497782 370896
rect 497816 370862 497872 370896
rect 497906 370862 497962 370896
rect 497996 370862 498052 370896
rect 498086 370862 498142 370896
rect 498176 370862 498289 370896
rect 497378 370850 498289 370862
rect 497327 370843 498289 370850
rect 498353 371804 498386 371838
rect 498420 371804 498452 371838
rect 498353 371748 498452 371804
rect 498353 371714 498386 371748
rect 498420 371714 498452 371748
rect 498353 371658 498452 371714
rect 498353 371624 498386 371658
rect 498420 371624 498452 371658
rect 498353 371568 498452 371624
rect 498353 371534 498386 371568
rect 498420 371534 498452 371568
rect 498353 371478 498452 371534
rect 498353 371444 498386 371478
rect 498420 371444 498452 371478
rect 498353 371388 498452 371444
rect 498353 371354 498386 371388
rect 498420 371354 498452 371388
rect 498353 371298 498452 371354
rect 498353 371264 498386 371298
rect 498420 371264 498452 371298
rect 498353 371208 498452 371264
rect 498353 371174 498386 371208
rect 498420 371174 498452 371208
rect 498353 371118 498452 371174
rect 498353 371084 498386 371118
rect 498420 371084 498452 371118
rect 498353 371028 498452 371084
rect 498353 370994 498386 371028
rect 498420 370994 498452 371028
rect 498353 370938 498452 370994
rect 498353 370904 498386 370938
rect 498420 370904 498452 370938
rect 498353 370848 498452 370904
rect 497164 370779 497263 370814
rect 498353 370814 498386 370848
rect 498420 370814 498452 370848
rect 498353 370779 498452 370814
rect 497164 370778 498452 370779
rect 497164 370744 497184 370778
rect 497218 370747 498452 370778
rect 497218 370744 497222 370747
rect 497164 370713 497222 370744
rect 497256 370713 497312 370747
rect 497346 370713 497402 370747
rect 497436 370713 497492 370747
rect 497526 370713 497582 370747
rect 497616 370713 497672 370747
rect 497706 370713 497762 370747
rect 497796 370713 497852 370747
rect 497886 370713 497942 370747
rect 497976 370713 498032 370747
rect 498066 370713 498122 370747
rect 498156 370713 498212 370747
rect 498246 370713 498302 370747
rect 498336 370713 498452 370747
rect 497164 370608 498452 370713
rect 497164 370574 497184 370608
rect 497218 370594 498452 370608
rect 497218 370574 497222 370594
rect 497164 370560 497222 370574
rect 497256 370560 497312 370594
rect 497346 370560 497402 370594
rect 497436 370560 497492 370594
rect 497526 370560 497582 370594
rect 497616 370560 497672 370594
rect 497706 370560 497762 370594
rect 497796 370560 497852 370594
rect 497886 370560 497942 370594
rect 497976 370560 498032 370594
rect 498066 370560 498122 370594
rect 498156 370560 498212 370594
rect 498246 370560 498302 370594
rect 498336 370560 498452 370594
rect 497164 370529 498452 370560
rect 497164 370518 497263 370529
rect 497164 370484 497184 370518
rect 497218 370498 497263 370518
rect 497164 370464 497199 370484
rect 497233 370464 497263 370498
rect 498353 370498 498452 370529
rect 497164 370428 497263 370464
rect 497164 370394 497184 370428
rect 497218 370408 497263 370428
rect 497164 370374 497199 370394
rect 497233 370374 497263 370408
rect 497164 370338 497263 370374
rect 497164 370304 497184 370338
rect 497218 370318 497263 370338
rect 497164 370284 497199 370304
rect 497233 370284 497263 370318
rect 497164 370248 497263 370284
rect 497164 370214 497184 370248
rect 497218 370228 497263 370248
rect 497164 370194 497199 370214
rect 497233 370194 497263 370228
rect 497164 370158 497263 370194
rect 497164 370124 497184 370158
rect 497218 370138 497263 370158
rect 497164 370104 497199 370124
rect 497233 370104 497263 370138
rect 497164 370068 497263 370104
rect 497164 370034 497184 370068
rect 497218 370048 497263 370068
rect 497164 370014 497199 370034
rect 497233 370014 497263 370048
rect 497164 369978 497263 370014
rect 497164 369944 497184 369978
rect 497218 369958 497263 369978
rect 497164 369924 497199 369944
rect 497233 369924 497263 369958
rect 497164 369888 497263 369924
rect 497164 369854 497184 369888
rect 497218 369868 497263 369888
rect 497164 369834 497199 369854
rect 497233 369834 497263 369868
rect 497164 369798 497263 369834
rect 497164 369764 497184 369798
rect 497218 369778 497263 369798
rect 497164 369744 497199 369764
rect 497233 369744 497263 369778
rect 497164 369708 497263 369744
rect 497164 369674 497184 369708
rect 497218 369688 497263 369708
rect 497164 369654 497199 369674
rect 497233 369654 497263 369688
rect 497164 369618 497263 369654
rect 497164 369584 497184 369618
rect 497218 369598 497263 369618
rect 497164 369564 497199 369584
rect 497233 369564 497263 369598
rect 497164 369528 497263 369564
rect 497164 369494 497184 369528
rect 497218 369508 497263 369528
rect 497164 369474 497199 369494
rect 497233 369474 497263 369508
rect 497327 370446 498289 370465
rect 497327 370444 497403 370446
rect 497327 370410 497344 370444
rect 497378 370412 497403 370444
rect 497437 370412 497493 370446
rect 497527 370412 497583 370446
rect 497617 370412 497673 370446
rect 497707 370412 497763 370446
rect 497797 370412 497853 370446
rect 497887 370412 497943 370446
rect 497977 370412 498033 370446
rect 498067 370412 498123 370446
rect 498157 370412 498289 370446
rect 497378 370410 498289 370412
rect 497327 370393 498289 370410
rect 497327 370354 497399 370393
rect 497327 370320 497344 370354
rect 497378 370334 497399 370354
rect 497327 370300 497346 370320
rect 497380 370300 497399 370334
rect 498217 370368 498289 370393
rect 498217 370334 498236 370368
rect 498270 370334 498289 370368
rect 497327 370264 497399 370300
rect 497327 370230 497344 370264
rect 497378 370244 497399 370264
rect 497327 370210 497346 370230
rect 497380 370210 497399 370244
rect 497327 370174 497399 370210
rect 497327 370140 497344 370174
rect 497378 370154 497399 370174
rect 497327 370120 497346 370140
rect 497380 370120 497399 370154
rect 497327 370084 497399 370120
rect 497327 370050 497344 370084
rect 497378 370064 497399 370084
rect 497327 370030 497346 370050
rect 497380 370030 497399 370064
rect 497327 369994 497399 370030
rect 497327 369960 497344 369994
rect 497378 369974 497399 369994
rect 497327 369940 497346 369960
rect 497380 369940 497399 369974
rect 497327 369904 497399 369940
rect 497327 369870 497344 369904
rect 497378 369884 497399 369904
rect 497327 369850 497346 369870
rect 497380 369850 497399 369884
rect 497327 369814 497399 369850
rect 497327 369780 497344 369814
rect 497378 369794 497399 369814
rect 497327 369760 497346 369780
rect 497380 369760 497399 369794
rect 497327 369724 497399 369760
rect 497327 369690 497344 369724
rect 497378 369704 497399 369724
rect 497327 369670 497346 369690
rect 497380 369670 497399 369704
rect 497327 369634 497399 369670
rect 497461 370270 498155 370331
rect 497461 370236 497520 370270
rect 497554 370258 497610 370270
rect 497582 370236 497610 370258
rect 497644 370258 497700 370270
rect 497644 370236 497648 370258
rect 497461 370224 497548 370236
rect 497582 370224 497648 370236
rect 497682 370236 497700 370258
rect 497734 370258 497790 370270
rect 497734 370236 497748 370258
rect 497682 370224 497748 370236
rect 497782 370236 497790 370258
rect 497824 370258 497880 370270
rect 497914 370258 497970 370270
rect 498004 370258 498060 370270
rect 497824 370236 497848 370258
rect 497914 370236 497948 370258
rect 498004 370236 498048 370258
rect 498094 370236 498155 370270
rect 497782 370224 497848 370236
rect 497882 370224 497948 370236
rect 497982 370224 498048 370236
rect 498082 370224 498155 370236
rect 497461 370180 498155 370224
rect 497461 370146 497520 370180
rect 497554 370158 497610 370180
rect 497582 370146 497610 370158
rect 497644 370158 497700 370180
rect 497644 370146 497648 370158
rect 497461 370124 497548 370146
rect 497582 370124 497648 370146
rect 497682 370146 497700 370158
rect 497734 370158 497790 370180
rect 497734 370146 497748 370158
rect 497682 370124 497748 370146
rect 497782 370146 497790 370158
rect 497824 370158 497880 370180
rect 497914 370158 497970 370180
rect 498004 370158 498060 370180
rect 497824 370146 497848 370158
rect 497914 370146 497948 370158
rect 498004 370146 498048 370158
rect 498094 370146 498155 370180
rect 497782 370124 497848 370146
rect 497882 370124 497948 370146
rect 497982 370124 498048 370146
rect 498082 370124 498155 370146
rect 497461 370090 498155 370124
rect 497461 370056 497520 370090
rect 497554 370058 497610 370090
rect 497582 370056 497610 370058
rect 497644 370058 497700 370090
rect 497644 370056 497648 370058
rect 497461 370024 497548 370056
rect 497582 370024 497648 370056
rect 497682 370056 497700 370058
rect 497734 370058 497790 370090
rect 497734 370056 497748 370058
rect 497682 370024 497748 370056
rect 497782 370056 497790 370058
rect 497824 370058 497880 370090
rect 497914 370058 497970 370090
rect 498004 370058 498060 370090
rect 497824 370056 497848 370058
rect 497914 370056 497948 370058
rect 498004 370056 498048 370058
rect 498094 370056 498155 370090
rect 497782 370024 497848 370056
rect 497882 370024 497948 370056
rect 497982 370024 498048 370056
rect 498082 370024 498155 370056
rect 497461 370000 498155 370024
rect 497461 369966 497520 370000
rect 497554 369966 497610 370000
rect 497644 369966 497700 370000
rect 497734 369966 497790 370000
rect 497824 369966 497880 370000
rect 497914 369966 497970 370000
rect 498004 369966 498060 370000
rect 498094 369966 498155 370000
rect 497461 369958 498155 369966
rect 497461 369924 497548 369958
rect 497582 369924 497648 369958
rect 497682 369924 497748 369958
rect 497782 369924 497848 369958
rect 497882 369924 497948 369958
rect 497982 369924 498048 369958
rect 498082 369924 498155 369958
rect 497461 369910 498155 369924
rect 497461 369876 497520 369910
rect 497554 369876 497610 369910
rect 497644 369876 497700 369910
rect 497734 369876 497790 369910
rect 497824 369876 497880 369910
rect 497914 369876 497970 369910
rect 498004 369876 498060 369910
rect 498094 369876 498155 369910
rect 497461 369858 498155 369876
rect 497461 369824 497548 369858
rect 497582 369824 497648 369858
rect 497682 369824 497748 369858
rect 497782 369824 497848 369858
rect 497882 369824 497948 369858
rect 497982 369824 498048 369858
rect 498082 369824 498155 369858
rect 497461 369820 498155 369824
rect 497461 369786 497520 369820
rect 497554 369786 497610 369820
rect 497644 369786 497700 369820
rect 497734 369786 497790 369820
rect 497824 369786 497880 369820
rect 497914 369786 497970 369820
rect 498004 369786 498060 369820
rect 498094 369786 498155 369820
rect 497461 369758 498155 369786
rect 497461 369730 497548 369758
rect 497582 369730 497648 369758
rect 497461 369696 497520 369730
rect 497582 369724 497610 369730
rect 497554 369696 497610 369724
rect 497644 369724 497648 369730
rect 497682 369730 497748 369758
rect 497682 369724 497700 369730
rect 497644 369696 497700 369724
rect 497734 369724 497748 369730
rect 497782 369730 497848 369758
rect 497882 369730 497948 369758
rect 497982 369730 498048 369758
rect 498082 369730 498155 369758
rect 497782 369724 497790 369730
rect 497734 369696 497790 369724
rect 497824 369724 497848 369730
rect 497914 369724 497948 369730
rect 498004 369724 498048 369730
rect 497824 369696 497880 369724
rect 497914 369696 497970 369724
rect 498004 369696 498060 369724
rect 498094 369696 498155 369730
rect 497461 369637 498155 369696
rect 498217 370278 498289 370334
rect 498217 370244 498236 370278
rect 498270 370244 498289 370278
rect 498217 370188 498289 370244
rect 498217 370154 498236 370188
rect 498270 370154 498289 370188
rect 498217 370098 498289 370154
rect 498217 370064 498236 370098
rect 498270 370064 498289 370098
rect 498217 370008 498289 370064
rect 498217 369974 498236 370008
rect 498270 369974 498289 370008
rect 498217 369918 498289 369974
rect 498217 369884 498236 369918
rect 498270 369884 498289 369918
rect 498217 369828 498289 369884
rect 498217 369794 498236 369828
rect 498270 369794 498289 369828
rect 498217 369738 498289 369794
rect 498217 369704 498236 369738
rect 498270 369704 498289 369738
rect 498217 369648 498289 369704
rect 497327 369600 497344 369634
rect 497378 369614 497399 369634
rect 497327 369580 497346 369600
rect 497380 369580 497399 369614
rect 497327 369575 497399 369580
rect 498217 369614 498236 369648
rect 498270 369614 498289 369648
rect 498217 369575 498289 369614
rect 497327 369556 498289 369575
rect 497327 369544 497422 369556
rect 497327 369510 497344 369544
rect 497378 369522 497422 369544
rect 497456 369522 497512 369556
rect 497546 369522 497602 369556
rect 497636 369522 497692 369556
rect 497726 369522 497782 369556
rect 497816 369522 497872 369556
rect 497906 369522 497962 369556
rect 497996 369522 498052 369556
rect 498086 369522 498142 369556
rect 498176 369522 498289 369556
rect 497378 369510 498289 369522
rect 497327 369503 498289 369510
rect 498353 370464 498386 370498
rect 498420 370464 498452 370498
rect 498353 370408 498452 370464
rect 498353 370374 498386 370408
rect 498420 370374 498452 370408
rect 498353 370318 498452 370374
rect 498353 370284 498386 370318
rect 498420 370284 498452 370318
rect 498353 370228 498452 370284
rect 498353 370194 498386 370228
rect 498420 370194 498452 370228
rect 498353 370138 498452 370194
rect 498353 370104 498386 370138
rect 498420 370104 498452 370138
rect 498353 370048 498452 370104
rect 498353 370014 498386 370048
rect 498420 370014 498452 370048
rect 498353 369958 498452 370014
rect 498353 369924 498386 369958
rect 498420 369924 498452 369958
rect 498353 369868 498452 369924
rect 498353 369834 498386 369868
rect 498420 369834 498452 369868
rect 498353 369778 498452 369834
rect 498353 369744 498386 369778
rect 498420 369744 498452 369778
rect 498353 369688 498452 369744
rect 498353 369654 498386 369688
rect 498420 369654 498452 369688
rect 498353 369598 498452 369654
rect 498353 369564 498386 369598
rect 498420 369564 498452 369598
rect 498353 369508 498452 369564
rect 497164 369439 497263 369474
rect 498353 369474 498386 369508
rect 498420 369474 498452 369508
rect 498353 369439 498452 369474
rect 497164 369438 498452 369439
rect 497164 369404 497184 369438
rect 497218 369407 498452 369438
rect 497218 369404 497222 369407
rect 497164 369373 497222 369404
rect 497256 369373 497312 369407
rect 497346 369373 497402 369407
rect 497436 369373 497492 369407
rect 497526 369373 497582 369407
rect 497616 369373 497672 369407
rect 497706 369373 497762 369407
rect 497796 369373 497852 369407
rect 497886 369373 497942 369407
rect 497976 369373 498032 369407
rect 498066 369373 498122 369407
rect 498156 369373 498212 369407
rect 498246 369373 498302 369407
rect 498336 369373 498452 369407
rect 497164 369268 498452 369373
rect 497164 369234 497184 369268
rect 497218 369254 498452 369268
rect 497218 369234 497222 369254
rect 497164 369220 497222 369234
rect 497256 369220 497312 369254
rect 497346 369220 497402 369254
rect 497436 369220 497492 369254
rect 497526 369220 497582 369254
rect 497616 369220 497672 369254
rect 497706 369220 497762 369254
rect 497796 369220 497852 369254
rect 497886 369220 497942 369254
rect 497976 369220 498032 369254
rect 498066 369220 498122 369254
rect 498156 369220 498212 369254
rect 498246 369220 498302 369254
rect 498336 369220 498452 369254
rect 497164 369189 498452 369220
rect 497164 369178 497263 369189
rect 497164 369144 497184 369178
rect 497218 369158 497263 369178
rect 497164 369124 497199 369144
rect 497233 369124 497263 369158
rect 498353 369158 498452 369189
rect 497164 369088 497263 369124
rect 497164 369054 497184 369088
rect 497218 369068 497263 369088
rect 497164 369034 497199 369054
rect 497233 369034 497263 369068
rect 497164 368998 497263 369034
rect 497164 368964 497184 368998
rect 497218 368978 497263 368998
rect 497164 368944 497199 368964
rect 497233 368944 497263 368978
rect 497164 368908 497263 368944
rect 497164 368874 497184 368908
rect 497218 368888 497263 368908
rect 497164 368854 497199 368874
rect 497233 368854 497263 368888
rect 497164 368818 497263 368854
rect 497164 368784 497184 368818
rect 497218 368798 497263 368818
rect 497164 368764 497199 368784
rect 497233 368764 497263 368798
rect 497164 368728 497263 368764
rect 497164 368694 497184 368728
rect 497218 368708 497263 368728
rect 497164 368674 497199 368694
rect 497233 368674 497263 368708
rect 497164 368638 497263 368674
rect 497164 368604 497184 368638
rect 497218 368618 497263 368638
rect 497164 368584 497199 368604
rect 497233 368584 497263 368618
rect 497164 368548 497263 368584
rect 497164 368514 497184 368548
rect 497218 368528 497263 368548
rect 497164 368494 497199 368514
rect 497233 368494 497263 368528
rect 497164 368458 497263 368494
rect 497164 368424 497184 368458
rect 497218 368438 497263 368458
rect 497164 368404 497199 368424
rect 497233 368404 497263 368438
rect 497164 368368 497263 368404
rect 497164 368334 497184 368368
rect 497218 368348 497263 368368
rect 497164 368314 497199 368334
rect 497233 368314 497263 368348
rect 497164 368278 497263 368314
rect 497164 368244 497184 368278
rect 497218 368258 497263 368278
rect 497164 368224 497199 368244
rect 497233 368224 497263 368258
rect 497164 368188 497263 368224
rect 497164 368154 497184 368188
rect 497218 368168 497263 368188
rect 497164 368134 497199 368154
rect 497233 368134 497263 368168
rect 497327 369106 498289 369125
rect 497327 369104 497403 369106
rect 497327 369070 497344 369104
rect 497378 369072 497403 369104
rect 497437 369072 497493 369106
rect 497527 369072 497583 369106
rect 497617 369072 497673 369106
rect 497707 369072 497763 369106
rect 497797 369072 497853 369106
rect 497887 369072 497943 369106
rect 497977 369072 498033 369106
rect 498067 369072 498123 369106
rect 498157 369072 498289 369106
rect 497378 369070 498289 369072
rect 497327 369053 498289 369070
rect 497327 369014 497399 369053
rect 497327 368980 497344 369014
rect 497378 368994 497399 369014
rect 497327 368960 497346 368980
rect 497380 368960 497399 368994
rect 498217 369028 498289 369053
rect 498217 368994 498236 369028
rect 498270 368994 498289 369028
rect 497327 368924 497399 368960
rect 497327 368890 497344 368924
rect 497378 368904 497399 368924
rect 497327 368870 497346 368890
rect 497380 368870 497399 368904
rect 497327 368834 497399 368870
rect 497327 368800 497344 368834
rect 497378 368814 497399 368834
rect 497327 368780 497346 368800
rect 497380 368780 497399 368814
rect 497327 368744 497399 368780
rect 497327 368710 497344 368744
rect 497378 368724 497399 368744
rect 497327 368690 497346 368710
rect 497380 368690 497399 368724
rect 497327 368654 497399 368690
rect 497327 368620 497344 368654
rect 497378 368634 497399 368654
rect 497327 368600 497346 368620
rect 497380 368600 497399 368634
rect 497327 368564 497399 368600
rect 497327 368530 497344 368564
rect 497378 368544 497399 368564
rect 497327 368510 497346 368530
rect 497380 368510 497399 368544
rect 497327 368474 497399 368510
rect 497327 368440 497344 368474
rect 497378 368454 497399 368474
rect 497327 368420 497346 368440
rect 497380 368420 497399 368454
rect 497327 368384 497399 368420
rect 497327 368350 497344 368384
rect 497378 368364 497399 368384
rect 497327 368330 497346 368350
rect 497380 368330 497399 368364
rect 497327 368294 497399 368330
rect 497461 368930 498155 368991
rect 497461 368896 497520 368930
rect 497554 368918 497610 368930
rect 497582 368896 497610 368918
rect 497644 368918 497700 368930
rect 497644 368896 497648 368918
rect 497461 368884 497548 368896
rect 497582 368884 497648 368896
rect 497682 368896 497700 368918
rect 497734 368918 497790 368930
rect 497734 368896 497748 368918
rect 497682 368884 497748 368896
rect 497782 368896 497790 368918
rect 497824 368918 497880 368930
rect 497914 368918 497970 368930
rect 498004 368918 498060 368930
rect 497824 368896 497848 368918
rect 497914 368896 497948 368918
rect 498004 368896 498048 368918
rect 498094 368896 498155 368930
rect 497782 368884 497848 368896
rect 497882 368884 497948 368896
rect 497982 368884 498048 368896
rect 498082 368884 498155 368896
rect 497461 368840 498155 368884
rect 497461 368806 497520 368840
rect 497554 368818 497610 368840
rect 497582 368806 497610 368818
rect 497644 368818 497700 368840
rect 497644 368806 497648 368818
rect 497461 368784 497548 368806
rect 497582 368784 497648 368806
rect 497682 368806 497700 368818
rect 497734 368818 497790 368840
rect 497734 368806 497748 368818
rect 497682 368784 497748 368806
rect 497782 368806 497790 368818
rect 497824 368818 497880 368840
rect 497914 368818 497970 368840
rect 498004 368818 498060 368840
rect 497824 368806 497848 368818
rect 497914 368806 497948 368818
rect 498004 368806 498048 368818
rect 498094 368806 498155 368840
rect 497782 368784 497848 368806
rect 497882 368784 497948 368806
rect 497982 368784 498048 368806
rect 498082 368784 498155 368806
rect 497461 368750 498155 368784
rect 497461 368716 497520 368750
rect 497554 368718 497610 368750
rect 497582 368716 497610 368718
rect 497644 368718 497700 368750
rect 497644 368716 497648 368718
rect 497461 368684 497548 368716
rect 497582 368684 497648 368716
rect 497682 368716 497700 368718
rect 497734 368718 497790 368750
rect 497734 368716 497748 368718
rect 497682 368684 497748 368716
rect 497782 368716 497790 368718
rect 497824 368718 497880 368750
rect 497914 368718 497970 368750
rect 498004 368718 498060 368750
rect 497824 368716 497848 368718
rect 497914 368716 497948 368718
rect 498004 368716 498048 368718
rect 498094 368716 498155 368750
rect 497782 368684 497848 368716
rect 497882 368684 497948 368716
rect 497982 368684 498048 368716
rect 498082 368684 498155 368716
rect 497461 368660 498155 368684
rect 497461 368626 497520 368660
rect 497554 368626 497610 368660
rect 497644 368626 497700 368660
rect 497734 368626 497790 368660
rect 497824 368626 497880 368660
rect 497914 368626 497970 368660
rect 498004 368626 498060 368660
rect 498094 368626 498155 368660
rect 497461 368618 498155 368626
rect 497461 368584 497548 368618
rect 497582 368584 497648 368618
rect 497682 368584 497748 368618
rect 497782 368584 497848 368618
rect 497882 368584 497948 368618
rect 497982 368584 498048 368618
rect 498082 368584 498155 368618
rect 497461 368570 498155 368584
rect 497461 368536 497520 368570
rect 497554 368536 497610 368570
rect 497644 368536 497700 368570
rect 497734 368536 497790 368570
rect 497824 368536 497880 368570
rect 497914 368536 497970 368570
rect 498004 368536 498060 368570
rect 498094 368536 498155 368570
rect 497461 368518 498155 368536
rect 497461 368484 497548 368518
rect 497582 368484 497648 368518
rect 497682 368484 497748 368518
rect 497782 368484 497848 368518
rect 497882 368484 497948 368518
rect 497982 368484 498048 368518
rect 498082 368484 498155 368518
rect 497461 368480 498155 368484
rect 497461 368446 497520 368480
rect 497554 368446 497610 368480
rect 497644 368446 497700 368480
rect 497734 368446 497790 368480
rect 497824 368446 497880 368480
rect 497914 368446 497970 368480
rect 498004 368446 498060 368480
rect 498094 368446 498155 368480
rect 497461 368418 498155 368446
rect 497461 368390 497548 368418
rect 497582 368390 497648 368418
rect 497461 368356 497520 368390
rect 497582 368384 497610 368390
rect 497554 368356 497610 368384
rect 497644 368384 497648 368390
rect 497682 368390 497748 368418
rect 497682 368384 497700 368390
rect 497644 368356 497700 368384
rect 497734 368384 497748 368390
rect 497782 368390 497848 368418
rect 497882 368390 497948 368418
rect 497982 368390 498048 368418
rect 498082 368390 498155 368418
rect 497782 368384 497790 368390
rect 497734 368356 497790 368384
rect 497824 368384 497848 368390
rect 497914 368384 497948 368390
rect 498004 368384 498048 368390
rect 497824 368356 497880 368384
rect 497914 368356 497970 368384
rect 498004 368356 498060 368384
rect 498094 368356 498155 368390
rect 497461 368297 498155 368356
rect 498217 368938 498289 368994
rect 498217 368904 498236 368938
rect 498270 368904 498289 368938
rect 498217 368848 498289 368904
rect 498217 368814 498236 368848
rect 498270 368814 498289 368848
rect 498217 368758 498289 368814
rect 498217 368724 498236 368758
rect 498270 368724 498289 368758
rect 498217 368668 498289 368724
rect 498217 368634 498236 368668
rect 498270 368634 498289 368668
rect 498217 368578 498289 368634
rect 498217 368544 498236 368578
rect 498270 368544 498289 368578
rect 498217 368488 498289 368544
rect 498217 368454 498236 368488
rect 498270 368454 498289 368488
rect 498217 368398 498289 368454
rect 498217 368364 498236 368398
rect 498270 368364 498289 368398
rect 498217 368308 498289 368364
rect 497327 368260 497344 368294
rect 497378 368274 497399 368294
rect 497327 368240 497346 368260
rect 497380 368240 497399 368274
rect 497327 368235 497399 368240
rect 498217 368274 498236 368308
rect 498270 368274 498289 368308
rect 498217 368235 498289 368274
rect 497327 368216 498289 368235
rect 497327 368204 497422 368216
rect 497327 368170 497344 368204
rect 497378 368182 497422 368204
rect 497456 368182 497512 368216
rect 497546 368182 497602 368216
rect 497636 368182 497692 368216
rect 497726 368182 497782 368216
rect 497816 368182 497872 368216
rect 497906 368182 497962 368216
rect 497996 368182 498052 368216
rect 498086 368182 498142 368216
rect 498176 368182 498289 368216
rect 497378 368170 498289 368182
rect 497327 368163 498289 368170
rect 498353 369124 498386 369158
rect 498420 369124 498452 369158
rect 498353 369068 498452 369124
rect 498353 369034 498386 369068
rect 498420 369034 498452 369068
rect 498353 368978 498452 369034
rect 498353 368944 498386 368978
rect 498420 368944 498452 368978
rect 498353 368888 498452 368944
rect 498353 368854 498386 368888
rect 498420 368854 498452 368888
rect 498353 368798 498452 368854
rect 498353 368764 498386 368798
rect 498420 368764 498452 368798
rect 498353 368708 498452 368764
rect 498353 368674 498386 368708
rect 498420 368674 498452 368708
rect 498353 368618 498452 368674
rect 498353 368584 498386 368618
rect 498420 368584 498452 368618
rect 498353 368528 498452 368584
rect 498353 368494 498386 368528
rect 498420 368494 498452 368528
rect 498353 368438 498452 368494
rect 498353 368404 498386 368438
rect 498420 368404 498452 368438
rect 498353 368348 498452 368404
rect 498353 368314 498386 368348
rect 498420 368314 498452 368348
rect 498353 368258 498452 368314
rect 498353 368224 498386 368258
rect 498420 368224 498452 368258
rect 498353 368168 498452 368224
rect 497164 368099 497263 368134
rect 498353 368134 498386 368168
rect 498420 368134 498452 368168
rect 498353 368099 498452 368134
rect 497164 368098 498452 368099
rect 497164 368064 497184 368098
rect 497218 368067 498452 368098
rect 497218 368064 497222 368067
rect 497164 368033 497222 368064
rect 497256 368033 497312 368067
rect 497346 368033 497402 368067
rect 497436 368033 497492 368067
rect 497526 368033 497582 368067
rect 497616 368033 497672 368067
rect 497706 368033 497762 368067
rect 497796 368033 497852 368067
rect 497886 368033 497942 368067
rect 497976 368033 498032 368067
rect 498066 368033 498122 368067
rect 498156 368033 498212 368067
rect 498246 368033 498302 368067
rect 498336 368033 498452 368067
rect 497164 367928 498452 368033
rect 497164 367894 497184 367928
rect 497218 367914 498452 367928
rect 497218 367894 497222 367914
rect 497164 367880 497222 367894
rect 497256 367880 497312 367914
rect 497346 367880 497402 367914
rect 497436 367880 497492 367914
rect 497526 367880 497582 367914
rect 497616 367880 497672 367914
rect 497706 367880 497762 367914
rect 497796 367880 497852 367914
rect 497886 367880 497942 367914
rect 497976 367880 498032 367914
rect 498066 367880 498122 367914
rect 498156 367880 498212 367914
rect 498246 367880 498302 367914
rect 498336 367880 498452 367914
rect 497164 367849 498452 367880
rect 497164 367838 497263 367849
rect 497164 367804 497184 367838
rect 497218 367818 497263 367838
rect 497164 367784 497199 367804
rect 497233 367784 497263 367818
rect 498353 367818 498452 367849
rect 497164 367748 497263 367784
rect 497164 367714 497184 367748
rect 497218 367728 497263 367748
rect 497164 367694 497199 367714
rect 497233 367694 497263 367728
rect 497164 367658 497263 367694
rect 497164 367624 497184 367658
rect 497218 367638 497263 367658
rect 497164 367604 497199 367624
rect 497233 367604 497263 367638
rect 497164 367568 497263 367604
rect 497164 367534 497184 367568
rect 497218 367548 497263 367568
rect 497164 367514 497199 367534
rect 497233 367514 497263 367548
rect 497164 367478 497263 367514
rect 497164 367444 497184 367478
rect 497218 367458 497263 367478
rect 497164 367424 497199 367444
rect 497233 367424 497263 367458
rect 497164 367388 497263 367424
rect 497164 367354 497184 367388
rect 497218 367368 497263 367388
rect 497164 367334 497199 367354
rect 497233 367334 497263 367368
rect 497164 367298 497263 367334
rect 497164 367264 497184 367298
rect 497218 367278 497263 367298
rect 497164 367244 497199 367264
rect 497233 367244 497263 367278
rect 497164 367208 497263 367244
rect 497164 367174 497184 367208
rect 497218 367188 497263 367208
rect 497164 367154 497199 367174
rect 497233 367154 497263 367188
rect 497164 367118 497263 367154
rect 497164 367084 497184 367118
rect 497218 367098 497263 367118
rect 497164 367064 497199 367084
rect 497233 367064 497263 367098
rect 497164 367028 497263 367064
rect 497164 366994 497184 367028
rect 497218 367008 497263 367028
rect 497164 366974 497199 366994
rect 497233 366974 497263 367008
rect 497164 366938 497263 366974
rect 497164 366904 497184 366938
rect 497218 366918 497263 366938
rect 497164 366884 497199 366904
rect 497233 366884 497263 366918
rect 497164 366848 497263 366884
rect 497164 366814 497184 366848
rect 497218 366828 497263 366848
rect 497164 366794 497199 366814
rect 497233 366794 497263 366828
rect 497327 367766 498289 367785
rect 497327 367764 497403 367766
rect 497327 367730 497344 367764
rect 497378 367732 497403 367764
rect 497437 367732 497493 367766
rect 497527 367732 497583 367766
rect 497617 367732 497673 367766
rect 497707 367732 497763 367766
rect 497797 367732 497853 367766
rect 497887 367732 497943 367766
rect 497977 367732 498033 367766
rect 498067 367732 498123 367766
rect 498157 367732 498289 367766
rect 497378 367730 498289 367732
rect 497327 367713 498289 367730
rect 497327 367674 497399 367713
rect 497327 367640 497344 367674
rect 497378 367654 497399 367674
rect 497327 367620 497346 367640
rect 497380 367620 497399 367654
rect 498217 367688 498289 367713
rect 498217 367654 498236 367688
rect 498270 367654 498289 367688
rect 497327 367584 497399 367620
rect 497327 367550 497344 367584
rect 497378 367564 497399 367584
rect 497327 367530 497346 367550
rect 497380 367530 497399 367564
rect 497327 367494 497399 367530
rect 497327 367460 497344 367494
rect 497378 367474 497399 367494
rect 497327 367440 497346 367460
rect 497380 367440 497399 367474
rect 497327 367404 497399 367440
rect 497327 367370 497344 367404
rect 497378 367384 497399 367404
rect 497327 367350 497346 367370
rect 497380 367350 497399 367384
rect 497327 367314 497399 367350
rect 497327 367280 497344 367314
rect 497378 367294 497399 367314
rect 497327 367260 497346 367280
rect 497380 367260 497399 367294
rect 497327 367224 497399 367260
rect 497327 367190 497344 367224
rect 497378 367204 497399 367224
rect 497327 367170 497346 367190
rect 497380 367170 497399 367204
rect 497327 367134 497399 367170
rect 497327 367100 497344 367134
rect 497378 367114 497399 367134
rect 497327 367080 497346 367100
rect 497380 367080 497399 367114
rect 497327 367044 497399 367080
rect 497327 367010 497344 367044
rect 497378 367024 497399 367044
rect 497327 366990 497346 367010
rect 497380 366990 497399 367024
rect 497327 366954 497399 366990
rect 497461 367590 498155 367651
rect 497461 367556 497520 367590
rect 497554 367578 497610 367590
rect 497582 367556 497610 367578
rect 497644 367578 497700 367590
rect 497644 367556 497648 367578
rect 497461 367544 497548 367556
rect 497582 367544 497648 367556
rect 497682 367556 497700 367578
rect 497734 367578 497790 367590
rect 497734 367556 497748 367578
rect 497682 367544 497748 367556
rect 497782 367556 497790 367578
rect 497824 367578 497880 367590
rect 497914 367578 497970 367590
rect 498004 367578 498060 367590
rect 497824 367556 497848 367578
rect 497914 367556 497948 367578
rect 498004 367556 498048 367578
rect 498094 367556 498155 367590
rect 497782 367544 497848 367556
rect 497882 367544 497948 367556
rect 497982 367544 498048 367556
rect 498082 367544 498155 367556
rect 497461 367500 498155 367544
rect 497461 367466 497520 367500
rect 497554 367478 497610 367500
rect 497582 367466 497610 367478
rect 497644 367478 497700 367500
rect 497644 367466 497648 367478
rect 497461 367444 497548 367466
rect 497582 367444 497648 367466
rect 497682 367466 497700 367478
rect 497734 367478 497790 367500
rect 497734 367466 497748 367478
rect 497682 367444 497748 367466
rect 497782 367466 497790 367478
rect 497824 367478 497880 367500
rect 497914 367478 497970 367500
rect 498004 367478 498060 367500
rect 497824 367466 497848 367478
rect 497914 367466 497948 367478
rect 498004 367466 498048 367478
rect 498094 367466 498155 367500
rect 497782 367444 497848 367466
rect 497882 367444 497948 367466
rect 497982 367444 498048 367466
rect 498082 367444 498155 367466
rect 497461 367410 498155 367444
rect 497461 367376 497520 367410
rect 497554 367378 497610 367410
rect 497582 367376 497610 367378
rect 497644 367378 497700 367410
rect 497644 367376 497648 367378
rect 497461 367344 497548 367376
rect 497582 367344 497648 367376
rect 497682 367376 497700 367378
rect 497734 367378 497790 367410
rect 497734 367376 497748 367378
rect 497682 367344 497748 367376
rect 497782 367376 497790 367378
rect 497824 367378 497880 367410
rect 497914 367378 497970 367410
rect 498004 367378 498060 367410
rect 497824 367376 497848 367378
rect 497914 367376 497948 367378
rect 498004 367376 498048 367378
rect 498094 367376 498155 367410
rect 497782 367344 497848 367376
rect 497882 367344 497948 367376
rect 497982 367344 498048 367376
rect 498082 367344 498155 367376
rect 497461 367320 498155 367344
rect 497461 367286 497520 367320
rect 497554 367286 497610 367320
rect 497644 367286 497700 367320
rect 497734 367286 497790 367320
rect 497824 367286 497880 367320
rect 497914 367286 497970 367320
rect 498004 367286 498060 367320
rect 498094 367286 498155 367320
rect 497461 367278 498155 367286
rect 497461 367244 497548 367278
rect 497582 367244 497648 367278
rect 497682 367244 497748 367278
rect 497782 367244 497848 367278
rect 497882 367244 497948 367278
rect 497982 367244 498048 367278
rect 498082 367244 498155 367278
rect 497461 367230 498155 367244
rect 497461 367196 497520 367230
rect 497554 367196 497610 367230
rect 497644 367196 497700 367230
rect 497734 367196 497790 367230
rect 497824 367196 497880 367230
rect 497914 367196 497970 367230
rect 498004 367196 498060 367230
rect 498094 367196 498155 367230
rect 497461 367178 498155 367196
rect 497461 367144 497548 367178
rect 497582 367144 497648 367178
rect 497682 367144 497748 367178
rect 497782 367144 497848 367178
rect 497882 367144 497948 367178
rect 497982 367144 498048 367178
rect 498082 367144 498155 367178
rect 497461 367140 498155 367144
rect 497461 367106 497520 367140
rect 497554 367106 497610 367140
rect 497644 367106 497700 367140
rect 497734 367106 497790 367140
rect 497824 367106 497880 367140
rect 497914 367106 497970 367140
rect 498004 367106 498060 367140
rect 498094 367106 498155 367140
rect 497461 367078 498155 367106
rect 497461 367050 497548 367078
rect 497582 367050 497648 367078
rect 497461 367016 497520 367050
rect 497582 367044 497610 367050
rect 497554 367016 497610 367044
rect 497644 367044 497648 367050
rect 497682 367050 497748 367078
rect 497682 367044 497700 367050
rect 497644 367016 497700 367044
rect 497734 367044 497748 367050
rect 497782 367050 497848 367078
rect 497882 367050 497948 367078
rect 497982 367050 498048 367078
rect 498082 367050 498155 367078
rect 497782 367044 497790 367050
rect 497734 367016 497790 367044
rect 497824 367044 497848 367050
rect 497914 367044 497948 367050
rect 498004 367044 498048 367050
rect 497824 367016 497880 367044
rect 497914 367016 497970 367044
rect 498004 367016 498060 367044
rect 498094 367016 498155 367050
rect 497461 366957 498155 367016
rect 498217 367598 498289 367654
rect 498217 367564 498236 367598
rect 498270 367564 498289 367598
rect 498217 367508 498289 367564
rect 498217 367474 498236 367508
rect 498270 367474 498289 367508
rect 498217 367418 498289 367474
rect 498217 367384 498236 367418
rect 498270 367384 498289 367418
rect 498217 367328 498289 367384
rect 498217 367294 498236 367328
rect 498270 367294 498289 367328
rect 498217 367238 498289 367294
rect 498217 367204 498236 367238
rect 498270 367204 498289 367238
rect 498217 367148 498289 367204
rect 498217 367114 498236 367148
rect 498270 367114 498289 367148
rect 498217 367058 498289 367114
rect 498217 367024 498236 367058
rect 498270 367024 498289 367058
rect 498217 366968 498289 367024
rect 497327 366920 497344 366954
rect 497378 366934 497399 366954
rect 497327 366900 497346 366920
rect 497380 366900 497399 366934
rect 497327 366895 497399 366900
rect 498217 366934 498236 366968
rect 498270 366934 498289 366968
rect 498217 366895 498289 366934
rect 497327 366876 498289 366895
rect 497327 366864 497422 366876
rect 497327 366830 497344 366864
rect 497378 366842 497422 366864
rect 497456 366842 497512 366876
rect 497546 366842 497602 366876
rect 497636 366842 497692 366876
rect 497726 366842 497782 366876
rect 497816 366842 497872 366876
rect 497906 366842 497962 366876
rect 497996 366842 498052 366876
rect 498086 366842 498142 366876
rect 498176 366842 498289 366876
rect 497378 366830 498289 366842
rect 497327 366823 498289 366830
rect 498353 367784 498386 367818
rect 498420 367784 498452 367818
rect 498353 367728 498452 367784
rect 498353 367694 498386 367728
rect 498420 367694 498452 367728
rect 498353 367638 498452 367694
rect 498353 367604 498386 367638
rect 498420 367604 498452 367638
rect 498353 367548 498452 367604
rect 498353 367514 498386 367548
rect 498420 367514 498452 367548
rect 498353 367458 498452 367514
rect 498353 367424 498386 367458
rect 498420 367424 498452 367458
rect 498353 367368 498452 367424
rect 498353 367334 498386 367368
rect 498420 367334 498452 367368
rect 498353 367278 498452 367334
rect 498353 367244 498386 367278
rect 498420 367244 498452 367278
rect 498353 367188 498452 367244
rect 498353 367154 498386 367188
rect 498420 367154 498452 367188
rect 498353 367098 498452 367154
rect 498353 367064 498386 367098
rect 498420 367064 498452 367098
rect 498353 367008 498452 367064
rect 498353 366974 498386 367008
rect 498420 366974 498452 367008
rect 498353 366918 498452 366974
rect 498353 366884 498386 366918
rect 498420 366884 498452 366918
rect 498353 366828 498452 366884
rect 497164 366759 497263 366794
rect 498353 366794 498386 366828
rect 498420 366794 498452 366828
rect 498353 366759 498452 366794
rect 497164 366758 498452 366759
rect 497164 366724 497184 366758
rect 497218 366727 498452 366758
rect 497218 366724 497222 366727
rect 497164 366693 497222 366724
rect 497256 366693 497312 366727
rect 497346 366693 497402 366727
rect 497436 366693 497492 366727
rect 497526 366693 497582 366727
rect 497616 366693 497672 366727
rect 497706 366693 497762 366727
rect 497796 366693 497852 366727
rect 497886 366693 497942 366727
rect 497976 366693 498032 366727
rect 498066 366693 498122 366727
rect 498156 366693 498212 366727
rect 498246 366693 498302 366727
rect 498336 366693 498452 366727
rect 497164 366588 498452 366693
rect 497164 366554 497184 366588
rect 497218 366574 498452 366588
rect 497218 366554 497222 366574
rect 497164 366540 497222 366554
rect 497256 366540 497312 366574
rect 497346 366540 497402 366574
rect 497436 366540 497492 366574
rect 497526 366540 497582 366574
rect 497616 366540 497672 366574
rect 497706 366540 497762 366574
rect 497796 366540 497852 366574
rect 497886 366540 497942 366574
rect 497976 366540 498032 366574
rect 498066 366540 498122 366574
rect 498156 366540 498212 366574
rect 498246 366540 498302 366574
rect 498336 366540 498452 366574
rect 497164 366509 498452 366540
rect 497164 366498 497263 366509
rect 497164 366464 497184 366498
rect 497218 366478 497263 366498
rect 497164 366444 497199 366464
rect 497233 366444 497263 366478
rect 498353 366478 498452 366509
rect 497164 366408 497263 366444
rect 497164 366374 497184 366408
rect 497218 366388 497263 366408
rect 497164 366354 497199 366374
rect 497233 366354 497263 366388
rect 497164 366318 497263 366354
rect 497164 366284 497184 366318
rect 497218 366298 497263 366318
rect 497164 366264 497199 366284
rect 497233 366264 497263 366298
rect 497164 366228 497263 366264
rect 497164 366194 497184 366228
rect 497218 366208 497263 366228
rect 497164 366174 497199 366194
rect 497233 366174 497263 366208
rect 497164 366138 497263 366174
rect 497164 366104 497184 366138
rect 497218 366118 497263 366138
rect 497164 366084 497199 366104
rect 497233 366084 497263 366118
rect 497164 366048 497263 366084
rect 497164 366014 497184 366048
rect 497218 366028 497263 366048
rect 497164 365994 497199 366014
rect 497233 365994 497263 366028
rect 497164 365958 497263 365994
rect 497164 365924 497184 365958
rect 497218 365938 497263 365958
rect 497164 365904 497199 365924
rect 497233 365904 497263 365938
rect 497164 365868 497263 365904
rect 497164 365834 497184 365868
rect 497218 365848 497263 365868
rect 497164 365814 497199 365834
rect 497233 365814 497263 365848
rect 497164 365778 497263 365814
rect 497164 365744 497184 365778
rect 497218 365758 497263 365778
rect 497164 365724 497199 365744
rect 497233 365724 497263 365758
rect 497164 365688 497263 365724
rect 497164 365654 497184 365688
rect 497218 365668 497263 365688
rect 497164 365634 497199 365654
rect 497233 365634 497263 365668
rect 497164 365598 497263 365634
rect 497164 365564 497184 365598
rect 497218 365578 497263 365598
rect 497164 365544 497199 365564
rect 497233 365544 497263 365578
rect 497164 365508 497263 365544
rect 497164 365474 497184 365508
rect 497218 365488 497263 365508
rect 497164 365454 497199 365474
rect 497233 365454 497263 365488
rect 497327 366426 498289 366445
rect 497327 366424 497403 366426
rect 497327 366390 497344 366424
rect 497378 366392 497403 366424
rect 497437 366392 497493 366426
rect 497527 366392 497583 366426
rect 497617 366392 497673 366426
rect 497707 366392 497763 366426
rect 497797 366392 497853 366426
rect 497887 366392 497943 366426
rect 497977 366392 498033 366426
rect 498067 366392 498123 366426
rect 498157 366392 498289 366426
rect 497378 366390 498289 366392
rect 497327 366373 498289 366390
rect 497327 366334 497399 366373
rect 497327 366300 497344 366334
rect 497378 366314 497399 366334
rect 497327 366280 497346 366300
rect 497380 366280 497399 366314
rect 498217 366348 498289 366373
rect 498217 366314 498236 366348
rect 498270 366314 498289 366348
rect 497327 366244 497399 366280
rect 497327 366210 497344 366244
rect 497378 366224 497399 366244
rect 497327 366190 497346 366210
rect 497380 366190 497399 366224
rect 497327 366154 497399 366190
rect 497327 366120 497344 366154
rect 497378 366134 497399 366154
rect 497327 366100 497346 366120
rect 497380 366100 497399 366134
rect 497327 366064 497399 366100
rect 497327 366030 497344 366064
rect 497378 366044 497399 366064
rect 497327 366010 497346 366030
rect 497380 366010 497399 366044
rect 497327 365974 497399 366010
rect 497327 365940 497344 365974
rect 497378 365954 497399 365974
rect 497327 365920 497346 365940
rect 497380 365920 497399 365954
rect 497327 365884 497399 365920
rect 497327 365850 497344 365884
rect 497378 365864 497399 365884
rect 497327 365830 497346 365850
rect 497380 365830 497399 365864
rect 497327 365794 497399 365830
rect 497327 365760 497344 365794
rect 497378 365774 497399 365794
rect 497327 365740 497346 365760
rect 497380 365740 497399 365774
rect 497327 365704 497399 365740
rect 497327 365670 497344 365704
rect 497378 365684 497399 365704
rect 497327 365650 497346 365670
rect 497380 365650 497399 365684
rect 497327 365614 497399 365650
rect 497461 366250 498155 366311
rect 497461 366216 497520 366250
rect 497554 366238 497610 366250
rect 497582 366216 497610 366238
rect 497644 366238 497700 366250
rect 497644 366216 497648 366238
rect 497461 366204 497548 366216
rect 497582 366204 497648 366216
rect 497682 366216 497700 366238
rect 497734 366238 497790 366250
rect 497734 366216 497748 366238
rect 497682 366204 497748 366216
rect 497782 366216 497790 366238
rect 497824 366238 497880 366250
rect 497914 366238 497970 366250
rect 498004 366238 498060 366250
rect 497824 366216 497848 366238
rect 497914 366216 497948 366238
rect 498004 366216 498048 366238
rect 498094 366216 498155 366250
rect 497782 366204 497848 366216
rect 497882 366204 497948 366216
rect 497982 366204 498048 366216
rect 498082 366204 498155 366216
rect 497461 366160 498155 366204
rect 497461 366126 497520 366160
rect 497554 366138 497610 366160
rect 497582 366126 497610 366138
rect 497644 366138 497700 366160
rect 497644 366126 497648 366138
rect 497461 366104 497548 366126
rect 497582 366104 497648 366126
rect 497682 366126 497700 366138
rect 497734 366138 497790 366160
rect 497734 366126 497748 366138
rect 497682 366104 497748 366126
rect 497782 366126 497790 366138
rect 497824 366138 497880 366160
rect 497914 366138 497970 366160
rect 498004 366138 498060 366160
rect 497824 366126 497848 366138
rect 497914 366126 497948 366138
rect 498004 366126 498048 366138
rect 498094 366126 498155 366160
rect 497782 366104 497848 366126
rect 497882 366104 497948 366126
rect 497982 366104 498048 366126
rect 498082 366104 498155 366126
rect 497461 366070 498155 366104
rect 497461 366036 497520 366070
rect 497554 366038 497610 366070
rect 497582 366036 497610 366038
rect 497644 366038 497700 366070
rect 497644 366036 497648 366038
rect 497461 366004 497548 366036
rect 497582 366004 497648 366036
rect 497682 366036 497700 366038
rect 497734 366038 497790 366070
rect 497734 366036 497748 366038
rect 497682 366004 497748 366036
rect 497782 366036 497790 366038
rect 497824 366038 497880 366070
rect 497914 366038 497970 366070
rect 498004 366038 498060 366070
rect 497824 366036 497848 366038
rect 497914 366036 497948 366038
rect 498004 366036 498048 366038
rect 498094 366036 498155 366070
rect 497782 366004 497848 366036
rect 497882 366004 497948 366036
rect 497982 366004 498048 366036
rect 498082 366004 498155 366036
rect 497461 365980 498155 366004
rect 497461 365946 497520 365980
rect 497554 365946 497610 365980
rect 497644 365946 497700 365980
rect 497734 365946 497790 365980
rect 497824 365946 497880 365980
rect 497914 365946 497970 365980
rect 498004 365946 498060 365980
rect 498094 365946 498155 365980
rect 497461 365938 498155 365946
rect 497461 365904 497548 365938
rect 497582 365904 497648 365938
rect 497682 365904 497748 365938
rect 497782 365904 497848 365938
rect 497882 365904 497948 365938
rect 497982 365904 498048 365938
rect 498082 365904 498155 365938
rect 497461 365890 498155 365904
rect 497461 365856 497520 365890
rect 497554 365856 497610 365890
rect 497644 365856 497700 365890
rect 497734 365856 497790 365890
rect 497824 365856 497880 365890
rect 497914 365856 497970 365890
rect 498004 365856 498060 365890
rect 498094 365856 498155 365890
rect 497461 365838 498155 365856
rect 497461 365804 497548 365838
rect 497582 365804 497648 365838
rect 497682 365804 497748 365838
rect 497782 365804 497848 365838
rect 497882 365804 497948 365838
rect 497982 365804 498048 365838
rect 498082 365804 498155 365838
rect 497461 365800 498155 365804
rect 497461 365766 497520 365800
rect 497554 365766 497610 365800
rect 497644 365766 497700 365800
rect 497734 365766 497790 365800
rect 497824 365766 497880 365800
rect 497914 365766 497970 365800
rect 498004 365766 498060 365800
rect 498094 365766 498155 365800
rect 497461 365738 498155 365766
rect 497461 365710 497548 365738
rect 497582 365710 497648 365738
rect 497461 365676 497520 365710
rect 497582 365704 497610 365710
rect 497554 365676 497610 365704
rect 497644 365704 497648 365710
rect 497682 365710 497748 365738
rect 497682 365704 497700 365710
rect 497644 365676 497700 365704
rect 497734 365704 497748 365710
rect 497782 365710 497848 365738
rect 497882 365710 497948 365738
rect 497982 365710 498048 365738
rect 498082 365710 498155 365738
rect 497782 365704 497790 365710
rect 497734 365676 497790 365704
rect 497824 365704 497848 365710
rect 497914 365704 497948 365710
rect 498004 365704 498048 365710
rect 497824 365676 497880 365704
rect 497914 365676 497970 365704
rect 498004 365676 498060 365704
rect 498094 365676 498155 365710
rect 497461 365617 498155 365676
rect 498217 366258 498289 366314
rect 498217 366224 498236 366258
rect 498270 366224 498289 366258
rect 498217 366168 498289 366224
rect 498217 366134 498236 366168
rect 498270 366134 498289 366168
rect 498217 366078 498289 366134
rect 498217 366044 498236 366078
rect 498270 366044 498289 366078
rect 498217 365988 498289 366044
rect 498217 365954 498236 365988
rect 498270 365954 498289 365988
rect 498217 365898 498289 365954
rect 498217 365864 498236 365898
rect 498270 365864 498289 365898
rect 498217 365808 498289 365864
rect 498217 365774 498236 365808
rect 498270 365774 498289 365808
rect 498217 365718 498289 365774
rect 498217 365684 498236 365718
rect 498270 365684 498289 365718
rect 498217 365628 498289 365684
rect 497327 365580 497344 365614
rect 497378 365594 497399 365614
rect 497327 365560 497346 365580
rect 497380 365560 497399 365594
rect 497327 365555 497399 365560
rect 498217 365594 498236 365628
rect 498270 365594 498289 365628
rect 498217 365555 498289 365594
rect 497327 365536 498289 365555
rect 497327 365524 497422 365536
rect 497327 365490 497344 365524
rect 497378 365502 497422 365524
rect 497456 365502 497512 365536
rect 497546 365502 497602 365536
rect 497636 365502 497692 365536
rect 497726 365502 497782 365536
rect 497816 365502 497872 365536
rect 497906 365502 497962 365536
rect 497996 365502 498052 365536
rect 498086 365502 498142 365536
rect 498176 365502 498289 365536
rect 497378 365490 498289 365502
rect 497327 365483 498289 365490
rect 498353 366444 498386 366478
rect 498420 366444 498452 366478
rect 498353 366388 498452 366444
rect 498353 366354 498386 366388
rect 498420 366354 498452 366388
rect 498353 366298 498452 366354
rect 498353 366264 498386 366298
rect 498420 366264 498452 366298
rect 498353 366208 498452 366264
rect 498353 366174 498386 366208
rect 498420 366174 498452 366208
rect 498353 366118 498452 366174
rect 498353 366084 498386 366118
rect 498420 366084 498452 366118
rect 498353 366028 498452 366084
rect 498353 365994 498386 366028
rect 498420 365994 498452 366028
rect 498353 365938 498452 365994
rect 498353 365904 498386 365938
rect 498420 365904 498452 365938
rect 498353 365848 498452 365904
rect 498353 365814 498386 365848
rect 498420 365814 498452 365848
rect 498353 365758 498452 365814
rect 498353 365724 498386 365758
rect 498420 365724 498452 365758
rect 498353 365668 498452 365724
rect 498353 365634 498386 365668
rect 498420 365634 498452 365668
rect 498353 365578 498452 365634
rect 498353 365544 498386 365578
rect 498420 365544 498452 365578
rect 498353 365488 498452 365544
rect 497164 365419 497263 365454
rect 498353 365454 498386 365488
rect 498420 365454 498452 365488
rect 498353 365419 498452 365454
rect 497164 365418 498452 365419
rect 497164 365384 497184 365418
rect 497218 365387 498452 365418
rect 497218 365384 497222 365387
rect 497164 365353 497222 365384
rect 497256 365353 497312 365387
rect 497346 365353 497402 365387
rect 497436 365353 497492 365387
rect 497526 365353 497582 365387
rect 497616 365353 497672 365387
rect 497706 365353 497762 365387
rect 497796 365353 497852 365387
rect 497886 365353 497942 365387
rect 497976 365353 498032 365387
rect 498066 365353 498122 365387
rect 498156 365353 498212 365387
rect 498246 365353 498302 365387
rect 498336 365353 498452 365387
rect 497164 365248 498452 365353
rect 497164 365214 497184 365248
rect 497218 365234 498452 365248
rect 497218 365214 497222 365234
rect 497164 365200 497222 365214
rect 497256 365200 497312 365234
rect 497346 365200 497402 365234
rect 497436 365200 497492 365234
rect 497526 365200 497582 365234
rect 497616 365200 497672 365234
rect 497706 365200 497762 365234
rect 497796 365200 497852 365234
rect 497886 365200 497942 365234
rect 497976 365200 498032 365234
rect 498066 365200 498122 365234
rect 498156 365200 498212 365234
rect 498246 365200 498302 365234
rect 498336 365200 498452 365234
rect 497164 365169 498452 365200
rect 497164 365158 497263 365169
rect 497164 365124 497184 365158
rect 497218 365138 497263 365158
rect 497164 365104 497199 365124
rect 497233 365104 497263 365138
rect 498353 365138 498452 365169
rect 497164 365068 497263 365104
rect 497164 365034 497184 365068
rect 497218 365048 497263 365068
rect 497164 365014 497199 365034
rect 497233 365014 497263 365048
rect 497164 364978 497263 365014
rect 497164 364944 497184 364978
rect 497218 364958 497263 364978
rect 497164 364924 497199 364944
rect 497233 364924 497263 364958
rect 497164 364888 497263 364924
rect 497164 364854 497184 364888
rect 497218 364868 497263 364888
rect 497164 364834 497199 364854
rect 497233 364834 497263 364868
rect 497164 364798 497263 364834
rect 497164 364764 497184 364798
rect 497218 364778 497263 364798
rect 497164 364744 497199 364764
rect 497233 364744 497263 364778
rect 497164 364708 497263 364744
rect 497164 364674 497184 364708
rect 497218 364688 497263 364708
rect 497164 364654 497199 364674
rect 497233 364654 497263 364688
rect 497164 364618 497263 364654
rect 497164 364584 497184 364618
rect 497218 364598 497263 364618
rect 497164 364564 497199 364584
rect 497233 364564 497263 364598
rect 497164 364528 497263 364564
rect 497164 364494 497184 364528
rect 497218 364508 497263 364528
rect 497164 364474 497199 364494
rect 497233 364474 497263 364508
rect 497164 364438 497263 364474
rect 497164 364404 497184 364438
rect 497218 364418 497263 364438
rect 497164 364384 497199 364404
rect 497233 364384 497263 364418
rect 497164 364348 497263 364384
rect 497164 364314 497184 364348
rect 497218 364328 497263 364348
rect 497164 364294 497199 364314
rect 497233 364294 497263 364328
rect 497164 364258 497263 364294
rect 497164 364224 497184 364258
rect 497218 364238 497263 364258
rect 497164 364204 497199 364224
rect 497233 364204 497263 364238
rect 497164 364168 497263 364204
rect 497164 364134 497184 364168
rect 497218 364148 497263 364168
rect 497164 364114 497199 364134
rect 497233 364114 497263 364148
rect 497327 365086 498289 365105
rect 497327 365084 497403 365086
rect 497327 365050 497344 365084
rect 497378 365052 497403 365084
rect 497437 365052 497493 365086
rect 497527 365052 497583 365086
rect 497617 365052 497673 365086
rect 497707 365052 497763 365086
rect 497797 365052 497853 365086
rect 497887 365052 497943 365086
rect 497977 365052 498033 365086
rect 498067 365052 498123 365086
rect 498157 365052 498289 365086
rect 497378 365050 498289 365052
rect 497327 365033 498289 365050
rect 497327 364994 497399 365033
rect 497327 364960 497344 364994
rect 497378 364974 497399 364994
rect 497327 364940 497346 364960
rect 497380 364940 497399 364974
rect 498217 365008 498289 365033
rect 498217 364974 498236 365008
rect 498270 364974 498289 365008
rect 497327 364904 497399 364940
rect 497327 364870 497344 364904
rect 497378 364884 497399 364904
rect 497327 364850 497346 364870
rect 497380 364850 497399 364884
rect 497327 364814 497399 364850
rect 497327 364780 497344 364814
rect 497378 364794 497399 364814
rect 497327 364760 497346 364780
rect 497380 364760 497399 364794
rect 497327 364724 497399 364760
rect 497327 364690 497344 364724
rect 497378 364704 497399 364724
rect 497327 364670 497346 364690
rect 497380 364670 497399 364704
rect 497327 364634 497399 364670
rect 497327 364600 497344 364634
rect 497378 364614 497399 364634
rect 497327 364580 497346 364600
rect 497380 364580 497399 364614
rect 497327 364544 497399 364580
rect 497327 364510 497344 364544
rect 497378 364524 497399 364544
rect 497327 364490 497346 364510
rect 497380 364490 497399 364524
rect 497327 364454 497399 364490
rect 497327 364420 497344 364454
rect 497378 364434 497399 364454
rect 497327 364400 497346 364420
rect 497380 364400 497399 364434
rect 497327 364364 497399 364400
rect 497327 364330 497344 364364
rect 497378 364344 497399 364364
rect 497327 364310 497346 364330
rect 497380 364310 497399 364344
rect 497327 364274 497399 364310
rect 497461 364910 498155 364971
rect 497461 364876 497520 364910
rect 497554 364898 497610 364910
rect 497582 364876 497610 364898
rect 497644 364898 497700 364910
rect 497644 364876 497648 364898
rect 497461 364864 497548 364876
rect 497582 364864 497648 364876
rect 497682 364876 497700 364898
rect 497734 364898 497790 364910
rect 497734 364876 497748 364898
rect 497682 364864 497748 364876
rect 497782 364876 497790 364898
rect 497824 364898 497880 364910
rect 497914 364898 497970 364910
rect 498004 364898 498060 364910
rect 497824 364876 497848 364898
rect 497914 364876 497948 364898
rect 498004 364876 498048 364898
rect 498094 364876 498155 364910
rect 497782 364864 497848 364876
rect 497882 364864 497948 364876
rect 497982 364864 498048 364876
rect 498082 364864 498155 364876
rect 497461 364820 498155 364864
rect 497461 364786 497520 364820
rect 497554 364798 497610 364820
rect 497582 364786 497610 364798
rect 497644 364798 497700 364820
rect 497644 364786 497648 364798
rect 497461 364764 497548 364786
rect 497582 364764 497648 364786
rect 497682 364786 497700 364798
rect 497734 364798 497790 364820
rect 497734 364786 497748 364798
rect 497682 364764 497748 364786
rect 497782 364786 497790 364798
rect 497824 364798 497880 364820
rect 497914 364798 497970 364820
rect 498004 364798 498060 364820
rect 497824 364786 497848 364798
rect 497914 364786 497948 364798
rect 498004 364786 498048 364798
rect 498094 364786 498155 364820
rect 497782 364764 497848 364786
rect 497882 364764 497948 364786
rect 497982 364764 498048 364786
rect 498082 364764 498155 364786
rect 497461 364730 498155 364764
rect 497461 364696 497520 364730
rect 497554 364698 497610 364730
rect 497582 364696 497610 364698
rect 497644 364698 497700 364730
rect 497644 364696 497648 364698
rect 497461 364664 497548 364696
rect 497582 364664 497648 364696
rect 497682 364696 497700 364698
rect 497734 364698 497790 364730
rect 497734 364696 497748 364698
rect 497682 364664 497748 364696
rect 497782 364696 497790 364698
rect 497824 364698 497880 364730
rect 497914 364698 497970 364730
rect 498004 364698 498060 364730
rect 497824 364696 497848 364698
rect 497914 364696 497948 364698
rect 498004 364696 498048 364698
rect 498094 364696 498155 364730
rect 497782 364664 497848 364696
rect 497882 364664 497948 364696
rect 497982 364664 498048 364696
rect 498082 364664 498155 364696
rect 497461 364640 498155 364664
rect 497461 364606 497520 364640
rect 497554 364606 497610 364640
rect 497644 364606 497700 364640
rect 497734 364606 497790 364640
rect 497824 364606 497880 364640
rect 497914 364606 497970 364640
rect 498004 364606 498060 364640
rect 498094 364606 498155 364640
rect 497461 364598 498155 364606
rect 497461 364564 497548 364598
rect 497582 364564 497648 364598
rect 497682 364564 497748 364598
rect 497782 364564 497848 364598
rect 497882 364564 497948 364598
rect 497982 364564 498048 364598
rect 498082 364564 498155 364598
rect 497461 364550 498155 364564
rect 497461 364516 497520 364550
rect 497554 364516 497610 364550
rect 497644 364516 497700 364550
rect 497734 364516 497790 364550
rect 497824 364516 497880 364550
rect 497914 364516 497970 364550
rect 498004 364516 498060 364550
rect 498094 364516 498155 364550
rect 497461 364498 498155 364516
rect 497461 364464 497548 364498
rect 497582 364464 497648 364498
rect 497682 364464 497748 364498
rect 497782 364464 497848 364498
rect 497882 364464 497948 364498
rect 497982 364464 498048 364498
rect 498082 364464 498155 364498
rect 497461 364460 498155 364464
rect 497461 364426 497520 364460
rect 497554 364426 497610 364460
rect 497644 364426 497700 364460
rect 497734 364426 497790 364460
rect 497824 364426 497880 364460
rect 497914 364426 497970 364460
rect 498004 364426 498060 364460
rect 498094 364426 498155 364460
rect 497461 364398 498155 364426
rect 497461 364370 497548 364398
rect 497582 364370 497648 364398
rect 497461 364336 497520 364370
rect 497582 364364 497610 364370
rect 497554 364336 497610 364364
rect 497644 364364 497648 364370
rect 497682 364370 497748 364398
rect 497682 364364 497700 364370
rect 497644 364336 497700 364364
rect 497734 364364 497748 364370
rect 497782 364370 497848 364398
rect 497882 364370 497948 364398
rect 497982 364370 498048 364398
rect 498082 364370 498155 364398
rect 497782 364364 497790 364370
rect 497734 364336 497790 364364
rect 497824 364364 497848 364370
rect 497914 364364 497948 364370
rect 498004 364364 498048 364370
rect 497824 364336 497880 364364
rect 497914 364336 497970 364364
rect 498004 364336 498060 364364
rect 498094 364336 498155 364370
rect 497461 364277 498155 364336
rect 498217 364918 498289 364974
rect 498217 364884 498236 364918
rect 498270 364884 498289 364918
rect 498217 364828 498289 364884
rect 498217 364794 498236 364828
rect 498270 364794 498289 364828
rect 498217 364738 498289 364794
rect 498217 364704 498236 364738
rect 498270 364704 498289 364738
rect 498217 364648 498289 364704
rect 498217 364614 498236 364648
rect 498270 364614 498289 364648
rect 498217 364558 498289 364614
rect 498217 364524 498236 364558
rect 498270 364524 498289 364558
rect 498217 364468 498289 364524
rect 498217 364434 498236 364468
rect 498270 364434 498289 364468
rect 498217 364378 498289 364434
rect 498217 364344 498236 364378
rect 498270 364344 498289 364378
rect 498217 364288 498289 364344
rect 497327 364240 497344 364274
rect 497378 364254 497399 364274
rect 497327 364220 497346 364240
rect 497380 364220 497399 364254
rect 497327 364215 497399 364220
rect 498217 364254 498236 364288
rect 498270 364254 498289 364288
rect 498217 364215 498289 364254
rect 497327 364196 498289 364215
rect 497327 364184 497422 364196
rect 497327 364150 497344 364184
rect 497378 364162 497422 364184
rect 497456 364162 497512 364196
rect 497546 364162 497602 364196
rect 497636 364162 497692 364196
rect 497726 364162 497782 364196
rect 497816 364162 497872 364196
rect 497906 364162 497962 364196
rect 497996 364162 498052 364196
rect 498086 364162 498142 364196
rect 498176 364162 498289 364196
rect 497378 364150 498289 364162
rect 497327 364143 498289 364150
rect 498353 365104 498386 365138
rect 498420 365104 498452 365138
rect 498353 365048 498452 365104
rect 498353 365014 498386 365048
rect 498420 365014 498452 365048
rect 498353 364958 498452 365014
rect 498353 364924 498386 364958
rect 498420 364924 498452 364958
rect 498353 364868 498452 364924
rect 498353 364834 498386 364868
rect 498420 364834 498452 364868
rect 498353 364778 498452 364834
rect 498353 364744 498386 364778
rect 498420 364744 498452 364778
rect 498353 364688 498452 364744
rect 498353 364654 498386 364688
rect 498420 364654 498452 364688
rect 498353 364598 498452 364654
rect 498353 364564 498386 364598
rect 498420 364564 498452 364598
rect 498353 364508 498452 364564
rect 498353 364474 498386 364508
rect 498420 364474 498452 364508
rect 498353 364418 498452 364474
rect 498353 364384 498386 364418
rect 498420 364384 498452 364418
rect 498353 364328 498452 364384
rect 498353 364294 498386 364328
rect 498420 364294 498452 364328
rect 498353 364238 498452 364294
rect 498353 364204 498386 364238
rect 498420 364204 498452 364238
rect 498353 364148 498452 364204
rect 497164 364079 497263 364114
rect 498353 364114 498386 364148
rect 498420 364114 498452 364148
rect 498353 364079 498452 364114
rect 497164 364078 498452 364079
rect 497164 364044 497184 364078
rect 497218 364047 498452 364078
rect 497218 364044 497222 364047
rect 497164 364013 497222 364044
rect 497256 364013 497312 364047
rect 497346 364013 497402 364047
rect 497436 364013 497492 364047
rect 497526 364013 497582 364047
rect 497616 364013 497672 364047
rect 497706 364013 497762 364047
rect 497796 364013 497852 364047
rect 497886 364013 497942 364047
rect 497976 364013 498032 364047
rect 498066 364013 498122 364047
rect 498156 364013 498212 364047
rect 498246 364013 498302 364047
rect 498336 364013 498452 364047
rect 497164 363908 498452 364013
rect 497164 363874 497184 363908
rect 497218 363894 498452 363908
rect 497218 363874 497222 363894
rect 497164 363860 497222 363874
rect 497256 363860 497312 363894
rect 497346 363860 497402 363894
rect 497436 363860 497492 363894
rect 497526 363860 497582 363894
rect 497616 363860 497672 363894
rect 497706 363860 497762 363894
rect 497796 363860 497852 363894
rect 497886 363860 497942 363894
rect 497976 363860 498032 363894
rect 498066 363860 498122 363894
rect 498156 363860 498212 363894
rect 498246 363860 498302 363894
rect 498336 363860 498452 363894
rect 497164 363829 498452 363860
rect 497164 363818 497263 363829
rect 497164 363784 497184 363818
rect 497218 363798 497263 363818
rect 497164 363764 497199 363784
rect 497233 363764 497263 363798
rect 498353 363798 498452 363829
rect 497164 363728 497263 363764
rect 497164 363694 497184 363728
rect 497218 363708 497263 363728
rect 497164 363674 497199 363694
rect 497233 363674 497263 363708
rect 497164 363638 497263 363674
rect 497164 363604 497184 363638
rect 497218 363618 497263 363638
rect 497164 363584 497199 363604
rect 497233 363584 497263 363618
rect 497164 363548 497263 363584
rect 497164 363514 497184 363548
rect 497218 363528 497263 363548
rect 497164 363494 497199 363514
rect 497233 363494 497263 363528
rect 497164 363458 497263 363494
rect 497164 363424 497184 363458
rect 497218 363438 497263 363458
rect 497164 363404 497199 363424
rect 497233 363404 497263 363438
rect 497164 363368 497263 363404
rect 497164 363334 497184 363368
rect 497218 363348 497263 363368
rect 497164 363314 497199 363334
rect 497233 363314 497263 363348
rect 497164 363278 497263 363314
rect 497164 363244 497184 363278
rect 497218 363258 497263 363278
rect 497164 363224 497199 363244
rect 497233 363224 497263 363258
rect 497164 363188 497263 363224
rect 497164 363154 497184 363188
rect 497218 363168 497263 363188
rect 497164 363134 497199 363154
rect 497233 363134 497263 363168
rect 497164 363098 497263 363134
rect 497164 363064 497184 363098
rect 497218 363078 497263 363098
rect 497164 363044 497199 363064
rect 497233 363044 497263 363078
rect 497164 363008 497263 363044
rect 497164 362974 497184 363008
rect 497218 362988 497263 363008
rect 497164 362954 497199 362974
rect 497233 362954 497263 362988
rect 497164 362918 497263 362954
rect 497164 362884 497184 362918
rect 497218 362898 497263 362918
rect 497164 362864 497199 362884
rect 497233 362864 497263 362898
rect 497164 362828 497263 362864
rect 497164 362794 497184 362828
rect 497218 362808 497263 362828
rect 497164 362774 497199 362794
rect 497233 362774 497263 362808
rect 497327 363746 498289 363765
rect 497327 363744 497403 363746
rect 497327 363710 497344 363744
rect 497378 363712 497403 363744
rect 497437 363712 497493 363746
rect 497527 363712 497583 363746
rect 497617 363712 497673 363746
rect 497707 363712 497763 363746
rect 497797 363712 497853 363746
rect 497887 363712 497943 363746
rect 497977 363712 498033 363746
rect 498067 363712 498123 363746
rect 498157 363712 498289 363746
rect 497378 363710 498289 363712
rect 497327 363693 498289 363710
rect 497327 363654 497399 363693
rect 497327 363620 497344 363654
rect 497378 363634 497399 363654
rect 497327 363600 497346 363620
rect 497380 363600 497399 363634
rect 498217 363668 498289 363693
rect 498217 363634 498236 363668
rect 498270 363634 498289 363668
rect 497327 363564 497399 363600
rect 497327 363530 497344 363564
rect 497378 363544 497399 363564
rect 497327 363510 497346 363530
rect 497380 363510 497399 363544
rect 497327 363474 497399 363510
rect 497327 363440 497344 363474
rect 497378 363454 497399 363474
rect 497327 363420 497346 363440
rect 497380 363420 497399 363454
rect 497327 363384 497399 363420
rect 497327 363350 497344 363384
rect 497378 363364 497399 363384
rect 497327 363330 497346 363350
rect 497380 363330 497399 363364
rect 497327 363294 497399 363330
rect 497327 363260 497344 363294
rect 497378 363274 497399 363294
rect 497327 363240 497346 363260
rect 497380 363240 497399 363274
rect 497327 363204 497399 363240
rect 497327 363170 497344 363204
rect 497378 363184 497399 363204
rect 497327 363150 497346 363170
rect 497380 363150 497399 363184
rect 497327 363114 497399 363150
rect 497327 363080 497344 363114
rect 497378 363094 497399 363114
rect 497327 363060 497346 363080
rect 497380 363060 497399 363094
rect 497327 363024 497399 363060
rect 497327 362990 497344 363024
rect 497378 363004 497399 363024
rect 497327 362970 497346 362990
rect 497380 362970 497399 363004
rect 497327 362934 497399 362970
rect 497461 363570 498155 363631
rect 497461 363536 497520 363570
rect 497554 363558 497610 363570
rect 497582 363536 497610 363558
rect 497644 363558 497700 363570
rect 497644 363536 497648 363558
rect 497461 363524 497548 363536
rect 497582 363524 497648 363536
rect 497682 363536 497700 363558
rect 497734 363558 497790 363570
rect 497734 363536 497748 363558
rect 497682 363524 497748 363536
rect 497782 363536 497790 363558
rect 497824 363558 497880 363570
rect 497914 363558 497970 363570
rect 498004 363558 498060 363570
rect 497824 363536 497848 363558
rect 497914 363536 497948 363558
rect 498004 363536 498048 363558
rect 498094 363536 498155 363570
rect 497782 363524 497848 363536
rect 497882 363524 497948 363536
rect 497982 363524 498048 363536
rect 498082 363524 498155 363536
rect 497461 363480 498155 363524
rect 497461 363446 497520 363480
rect 497554 363458 497610 363480
rect 497582 363446 497610 363458
rect 497644 363458 497700 363480
rect 497644 363446 497648 363458
rect 497461 363424 497548 363446
rect 497582 363424 497648 363446
rect 497682 363446 497700 363458
rect 497734 363458 497790 363480
rect 497734 363446 497748 363458
rect 497682 363424 497748 363446
rect 497782 363446 497790 363458
rect 497824 363458 497880 363480
rect 497914 363458 497970 363480
rect 498004 363458 498060 363480
rect 497824 363446 497848 363458
rect 497914 363446 497948 363458
rect 498004 363446 498048 363458
rect 498094 363446 498155 363480
rect 497782 363424 497848 363446
rect 497882 363424 497948 363446
rect 497982 363424 498048 363446
rect 498082 363424 498155 363446
rect 497461 363390 498155 363424
rect 497461 363356 497520 363390
rect 497554 363358 497610 363390
rect 497582 363356 497610 363358
rect 497644 363358 497700 363390
rect 497644 363356 497648 363358
rect 497461 363324 497548 363356
rect 497582 363324 497648 363356
rect 497682 363356 497700 363358
rect 497734 363358 497790 363390
rect 497734 363356 497748 363358
rect 497682 363324 497748 363356
rect 497782 363356 497790 363358
rect 497824 363358 497880 363390
rect 497914 363358 497970 363390
rect 498004 363358 498060 363390
rect 497824 363356 497848 363358
rect 497914 363356 497948 363358
rect 498004 363356 498048 363358
rect 498094 363356 498155 363390
rect 497782 363324 497848 363356
rect 497882 363324 497948 363356
rect 497982 363324 498048 363356
rect 498082 363324 498155 363356
rect 497461 363300 498155 363324
rect 497461 363266 497520 363300
rect 497554 363266 497610 363300
rect 497644 363266 497700 363300
rect 497734 363266 497790 363300
rect 497824 363266 497880 363300
rect 497914 363266 497970 363300
rect 498004 363266 498060 363300
rect 498094 363266 498155 363300
rect 497461 363258 498155 363266
rect 497461 363224 497548 363258
rect 497582 363224 497648 363258
rect 497682 363224 497748 363258
rect 497782 363224 497848 363258
rect 497882 363224 497948 363258
rect 497982 363224 498048 363258
rect 498082 363224 498155 363258
rect 497461 363210 498155 363224
rect 497461 363176 497520 363210
rect 497554 363176 497610 363210
rect 497644 363176 497700 363210
rect 497734 363176 497790 363210
rect 497824 363176 497880 363210
rect 497914 363176 497970 363210
rect 498004 363176 498060 363210
rect 498094 363176 498155 363210
rect 497461 363158 498155 363176
rect 497461 363124 497548 363158
rect 497582 363124 497648 363158
rect 497682 363124 497748 363158
rect 497782 363124 497848 363158
rect 497882 363124 497948 363158
rect 497982 363124 498048 363158
rect 498082 363124 498155 363158
rect 497461 363120 498155 363124
rect 497461 363086 497520 363120
rect 497554 363086 497610 363120
rect 497644 363086 497700 363120
rect 497734 363086 497790 363120
rect 497824 363086 497880 363120
rect 497914 363086 497970 363120
rect 498004 363086 498060 363120
rect 498094 363086 498155 363120
rect 497461 363058 498155 363086
rect 497461 363030 497548 363058
rect 497582 363030 497648 363058
rect 497461 362996 497520 363030
rect 497582 363024 497610 363030
rect 497554 362996 497610 363024
rect 497644 363024 497648 363030
rect 497682 363030 497748 363058
rect 497682 363024 497700 363030
rect 497644 362996 497700 363024
rect 497734 363024 497748 363030
rect 497782 363030 497848 363058
rect 497882 363030 497948 363058
rect 497982 363030 498048 363058
rect 498082 363030 498155 363058
rect 497782 363024 497790 363030
rect 497734 362996 497790 363024
rect 497824 363024 497848 363030
rect 497914 363024 497948 363030
rect 498004 363024 498048 363030
rect 497824 362996 497880 363024
rect 497914 362996 497970 363024
rect 498004 362996 498060 363024
rect 498094 362996 498155 363030
rect 497461 362937 498155 362996
rect 498217 363578 498289 363634
rect 498217 363544 498236 363578
rect 498270 363544 498289 363578
rect 498217 363488 498289 363544
rect 498217 363454 498236 363488
rect 498270 363454 498289 363488
rect 498217 363398 498289 363454
rect 498217 363364 498236 363398
rect 498270 363364 498289 363398
rect 498217 363308 498289 363364
rect 498217 363274 498236 363308
rect 498270 363274 498289 363308
rect 498217 363218 498289 363274
rect 498217 363184 498236 363218
rect 498270 363184 498289 363218
rect 498217 363128 498289 363184
rect 498217 363094 498236 363128
rect 498270 363094 498289 363128
rect 498217 363038 498289 363094
rect 498217 363004 498236 363038
rect 498270 363004 498289 363038
rect 498217 362948 498289 363004
rect 497327 362900 497344 362934
rect 497378 362914 497399 362934
rect 497327 362880 497346 362900
rect 497380 362880 497399 362914
rect 497327 362875 497399 362880
rect 498217 362914 498236 362948
rect 498270 362914 498289 362948
rect 498217 362875 498289 362914
rect 497327 362856 498289 362875
rect 497327 362844 497422 362856
rect 497327 362810 497344 362844
rect 497378 362822 497422 362844
rect 497456 362822 497512 362856
rect 497546 362822 497602 362856
rect 497636 362822 497692 362856
rect 497726 362822 497782 362856
rect 497816 362822 497872 362856
rect 497906 362822 497962 362856
rect 497996 362822 498052 362856
rect 498086 362822 498142 362856
rect 498176 362822 498289 362856
rect 497378 362810 498289 362822
rect 497327 362803 498289 362810
rect 498353 363764 498386 363798
rect 498420 363764 498452 363798
rect 498353 363708 498452 363764
rect 498353 363674 498386 363708
rect 498420 363674 498452 363708
rect 498353 363618 498452 363674
rect 498353 363584 498386 363618
rect 498420 363584 498452 363618
rect 498353 363528 498452 363584
rect 498353 363494 498386 363528
rect 498420 363494 498452 363528
rect 498353 363438 498452 363494
rect 498353 363404 498386 363438
rect 498420 363404 498452 363438
rect 498353 363348 498452 363404
rect 498353 363314 498386 363348
rect 498420 363314 498452 363348
rect 498353 363258 498452 363314
rect 498353 363224 498386 363258
rect 498420 363224 498452 363258
rect 498353 363168 498452 363224
rect 498353 363134 498386 363168
rect 498420 363134 498452 363168
rect 498353 363078 498452 363134
rect 498353 363044 498386 363078
rect 498420 363044 498452 363078
rect 498353 362988 498452 363044
rect 498353 362954 498386 362988
rect 498420 362954 498452 362988
rect 498353 362898 498452 362954
rect 498353 362864 498386 362898
rect 498420 362864 498452 362898
rect 498353 362808 498452 362864
rect 497164 362739 497263 362774
rect 498353 362774 498386 362808
rect 498420 362774 498452 362808
rect 498353 362739 498452 362774
rect 497164 362738 498452 362739
rect 497164 362704 497184 362738
rect 497218 362707 498452 362738
rect 497218 362704 497222 362707
rect 497164 362673 497222 362704
rect 497256 362673 497312 362707
rect 497346 362673 497402 362707
rect 497436 362673 497492 362707
rect 497526 362673 497582 362707
rect 497616 362673 497672 362707
rect 497706 362673 497762 362707
rect 497796 362673 497852 362707
rect 497886 362673 497942 362707
rect 497976 362673 498032 362707
rect 498066 362673 498122 362707
rect 498156 362673 498212 362707
rect 498246 362673 498302 362707
rect 498336 362673 498452 362707
rect 497164 362640 498452 362673
rect 498718 371811 498778 371994
rect 498718 371777 498731 371811
rect 498765 371777 498778 371811
rect 498718 371611 498778 371777
rect 498718 371577 498731 371611
rect 498765 371577 498778 371611
rect 498718 371411 498778 371577
rect 498718 371377 498731 371411
rect 498765 371377 498778 371411
rect 498718 371211 498778 371377
rect 498718 371177 498731 371211
rect 498765 371177 498778 371211
rect 498718 371011 498778 371177
rect 498718 370977 498731 371011
rect 498765 370977 498778 371011
rect 498718 370811 498778 370977
rect 498718 370777 498731 370811
rect 498765 370777 498778 370811
rect 498718 370611 498778 370777
rect 498718 370577 498731 370611
rect 498765 370577 498778 370611
rect 498718 370411 498778 370577
rect 498718 370377 498731 370411
rect 498765 370377 498778 370411
rect 498718 370211 498778 370377
rect 498718 370177 498731 370211
rect 498765 370177 498778 370211
rect 498718 370011 498778 370177
rect 498718 369977 498731 370011
rect 498765 369977 498778 370011
rect 498718 369811 498778 369977
rect 498718 369777 498731 369811
rect 498765 369777 498778 369811
rect 498718 369611 498778 369777
rect 498718 369577 498731 369611
rect 498765 369577 498778 369611
rect 498718 369411 498778 369577
rect 498718 369377 498731 369411
rect 498765 369377 498778 369411
rect 498718 369211 498778 369377
rect 498718 369177 498731 369211
rect 498765 369177 498778 369211
rect 498718 369011 498778 369177
rect 498718 368977 498731 369011
rect 498765 368977 498778 369011
rect 498718 368811 498778 368977
rect 498718 368777 498731 368811
rect 498765 368777 498778 368811
rect 498718 368611 498778 368777
rect 498718 368577 498731 368611
rect 498765 368577 498778 368611
rect 498718 368411 498778 368577
rect 498718 368377 498731 368411
rect 498765 368377 498778 368411
rect 498718 368211 498778 368377
rect 498718 368177 498731 368211
rect 498765 368177 498778 368211
rect 498718 368011 498778 368177
rect 498718 367977 498731 368011
rect 498765 367977 498778 368011
rect 498718 367811 498778 367977
rect 498718 367777 498731 367811
rect 498765 367777 498778 367811
rect 498718 367611 498778 367777
rect 498718 367577 498731 367611
rect 498765 367577 498778 367611
rect 498718 367411 498778 367577
rect 498718 367377 498731 367411
rect 498765 367377 498778 367411
rect 498718 367211 498778 367377
rect 498718 367177 498731 367211
rect 498765 367177 498778 367211
rect 498718 367011 498778 367177
rect 498718 366977 498731 367011
rect 498765 366977 498778 367011
rect 498718 366811 498778 366977
rect 498718 366777 498731 366811
rect 498765 366777 498778 366811
rect 498718 366611 498778 366777
rect 498718 366577 498731 366611
rect 498765 366577 498778 366611
rect 498718 366411 498778 366577
rect 498718 366377 498731 366411
rect 498765 366377 498778 366411
rect 498718 366211 498778 366377
rect 498718 366177 498731 366211
rect 498765 366177 498778 366211
rect 498718 366011 498778 366177
rect 498718 365977 498731 366011
rect 498765 365977 498778 366011
rect 498718 365811 498778 365977
rect 498718 365777 498731 365811
rect 498765 365777 498778 365811
rect 498718 365611 498778 365777
rect 498718 365577 498731 365611
rect 498765 365577 498778 365611
rect 498718 365411 498778 365577
rect 498718 365377 498731 365411
rect 498765 365377 498778 365411
rect 498718 365211 498778 365377
rect 498718 365177 498731 365211
rect 498765 365177 498778 365211
rect 498718 365011 498778 365177
rect 498718 364977 498731 365011
rect 498765 364977 498778 365011
rect 498718 364811 498778 364977
rect 498718 364777 498731 364811
rect 498765 364777 498778 364811
rect 498718 364611 498778 364777
rect 498718 364577 498731 364611
rect 498765 364577 498778 364611
rect 498718 364411 498778 364577
rect 498718 364377 498731 364411
rect 498765 364377 498778 364411
rect 498718 364211 498778 364377
rect 498718 364177 498731 364211
rect 498765 364177 498778 364211
rect 498718 364011 498778 364177
rect 498718 363977 498731 364011
rect 498765 363977 498778 364011
rect 498718 363811 498778 363977
rect 498718 363777 498731 363811
rect 498765 363777 498778 363811
rect 498718 363611 498778 363777
rect 498718 363577 498731 363611
rect 498765 363577 498778 363611
rect 498718 363411 498778 363577
rect 498718 363377 498731 363411
rect 498765 363377 498778 363411
rect 498718 363211 498778 363377
rect 498718 363177 498731 363211
rect 498765 363177 498778 363211
rect 498718 363011 498778 363177
rect 498718 362977 498731 363011
rect 498765 362977 498778 363011
rect 498718 362811 498778 362977
rect 498718 362777 498731 362811
rect 498765 362777 498778 362811
rect 498718 362614 498778 362777
rect 500598 371987 500658 372153
rect 500598 371953 500611 371987
rect 500645 371953 500658 371987
rect 500598 371787 500658 371953
rect 500598 371753 500611 371787
rect 500645 371753 500658 371787
rect 500598 371587 500658 371753
rect 500598 371553 500611 371587
rect 500645 371553 500658 371587
rect 500598 371387 500658 371553
rect 500598 371353 500611 371387
rect 500645 371353 500658 371387
rect 500598 371187 500658 371353
rect 500598 371153 500611 371187
rect 500645 371153 500658 371187
rect 500598 370987 500658 371153
rect 500598 370953 500611 370987
rect 500645 370953 500658 370987
rect 500598 370787 500658 370953
rect 500598 370753 500611 370787
rect 500645 370753 500658 370787
rect 500598 370587 500658 370753
rect 500598 370553 500611 370587
rect 500645 370553 500658 370587
rect 500598 370387 500658 370553
rect 500598 370353 500611 370387
rect 500645 370353 500658 370387
rect 500598 370187 500658 370353
rect 500598 370153 500611 370187
rect 500645 370153 500658 370187
rect 500598 369987 500658 370153
rect 500598 369953 500611 369987
rect 500645 369953 500658 369987
rect 500598 369787 500658 369953
rect 500598 369753 500611 369787
rect 500645 369753 500658 369787
rect 500598 369587 500658 369753
rect 500598 369553 500611 369587
rect 500645 369553 500658 369587
rect 500598 369387 500658 369553
rect 500598 369353 500611 369387
rect 500645 369353 500658 369387
rect 500598 369187 500658 369353
rect 500598 369153 500611 369187
rect 500645 369153 500658 369187
rect 500598 368987 500658 369153
rect 500598 368953 500611 368987
rect 500645 368953 500658 368987
rect 500598 368787 500658 368953
rect 500598 368753 500611 368787
rect 500645 368753 500658 368787
rect 500598 368587 500658 368753
rect 500598 368553 500611 368587
rect 500645 368553 500658 368587
rect 500598 368387 500658 368553
rect 500598 368353 500611 368387
rect 500645 368353 500658 368387
rect 500598 368187 500658 368353
rect 500598 368153 500611 368187
rect 500645 368153 500658 368187
rect 500598 367987 500658 368153
rect 500598 367953 500611 367987
rect 500645 367953 500658 367987
rect 500598 367787 500658 367953
rect 500598 367753 500611 367787
rect 500645 367753 500658 367787
rect 500598 367587 500658 367753
rect 500598 367553 500611 367587
rect 500645 367553 500658 367587
rect 500598 367387 500658 367553
rect 500598 367353 500611 367387
rect 500645 367353 500658 367387
rect 500598 367187 500658 367353
rect 500598 367153 500611 367187
rect 500645 367153 500658 367187
rect 500598 366987 500658 367153
rect 500598 366953 500611 366987
rect 500645 366953 500658 366987
rect 500598 366787 500658 366953
rect 500598 366753 500611 366787
rect 500645 366753 500658 366787
rect 500598 366587 500658 366753
rect 500598 366553 500611 366587
rect 500645 366553 500658 366587
rect 500598 366387 500658 366553
rect 500598 366353 500611 366387
rect 500645 366353 500658 366387
rect 500598 366187 500658 366353
rect 500598 366153 500611 366187
rect 500645 366153 500658 366187
rect 500598 365987 500658 366153
rect 500598 365953 500611 365987
rect 500645 365953 500658 365987
rect 500598 365787 500658 365953
rect 500598 365753 500611 365787
rect 500645 365753 500658 365787
rect 500598 365587 500658 365753
rect 500598 365553 500611 365587
rect 500645 365553 500658 365587
rect 500598 365387 500658 365553
rect 500598 365353 500611 365387
rect 500645 365353 500658 365387
rect 500598 365187 500658 365353
rect 500598 365153 500611 365187
rect 500645 365153 500658 365187
rect 500598 364987 500658 365153
rect 500598 364953 500611 364987
rect 500645 364953 500658 364987
rect 500598 364787 500658 364953
rect 500598 364753 500611 364787
rect 500645 364753 500658 364787
rect 500598 364587 500658 364753
rect 500598 364553 500611 364587
rect 500645 364553 500658 364587
rect 500598 364387 500658 364553
rect 500598 364353 500611 364387
rect 500645 364353 500658 364387
rect 500598 364187 500658 364353
rect 500598 364153 500611 364187
rect 500645 364153 500658 364187
rect 500598 363987 500658 364153
rect 500598 363953 500611 363987
rect 500645 363953 500658 363987
rect 500598 363787 500658 363953
rect 500598 363753 500611 363787
rect 500645 363753 500658 363787
rect 500598 363587 500658 363753
rect 500598 363553 500611 363587
rect 500645 363553 500658 363587
rect 500598 363387 500658 363553
rect 500598 363353 500611 363387
rect 500645 363353 500658 363387
rect 500598 363187 500658 363353
rect 500598 363153 500611 363187
rect 500645 363153 500658 363187
rect 500598 362987 500658 363153
rect 500598 362953 500611 362987
rect 500645 362953 500658 362987
rect 500598 362787 500658 362953
rect 500598 362753 500611 362787
rect 500645 362753 500658 362787
rect 500598 362587 500658 362753
rect 500598 362553 500611 362587
rect 500645 362553 500658 362587
rect 500598 362450 500658 362553
rect 500924 373124 502212 373144
rect 500924 373090 500944 373124
rect 500978 373110 502212 373124
rect 500978 373090 500982 373110
rect 500924 373076 500982 373090
rect 501016 373076 501072 373110
rect 501106 373076 501162 373110
rect 501196 373076 501252 373110
rect 501286 373076 501342 373110
rect 501376 373076 501432 373110
rect 501466 373076 501522 373110
rect 501556 373076 501612 373110
rect 501646 373076 501702 373110
rect 501736 373076 501792 373110
rect 501826 373076 501882 373110
rect 501916 373076 501972 373110
rect 502006 373076 502062 373110
rect 502096 373076 502212 373110
rect 500924 373045 502212 373076
rect 500924 373034 501023 373045
rect 500924 373000 500944 373034
rect 500978 373014 501023 373034
rect 500924 372980 500959 373000
rect 500993 372980 501023 373014
rect 502113 373014 502212 373045
rect 500924 372944 501023 372980
rect 500924 372910 500944 372944
rect 500978 372924 501023 372944
rect 500924 372890 500959 372910
rect 500993 372890 501023 372924
rect 500924 372854 501023 372890
rect 500924 372820 500944 372854
rect 500978 372834 501023 372854
rect 500924 372800 500959 372820
rect 500993 372800 501023 372834
rect 500924 372764 501023 372800
rect 500924 372730 500944 372764
rect 500978 372744 501023 372764
rect 500924 372710 500959 372730
rect 500993 372710 501023 372744
rect 500924 372674 501023 372710
rect 500924 372640 500944 372674
rect 500978 372654 501023 372674
rect 500924 372620 500959 372640
rect 500993 372620 501023 372654
rect 500924 372584 501023 372620
rect 500924 372550 500944 372584
rect 500978 372564 501023 372584
rect 500924 372530 500959 372550
rect 500993 372530 501023 372564
rect 500924 372494 501023 372530
rect 500924 372460 500944 372494
rect 500978 372474 501023 372494
rect 500924 372440 500959 372460
rect 500993 372440 501023 372474
rect 500924 372404 501023 372440
rect 500924 372370 500944 372404
rect 500978 372384 501023 372404
rect 500924 372350 500959 372370
rect 500993 372350 501023 372384
rect 500924 372314 501023 372350
rect 500924 372280 500944 372314
rect 500978 372294 501023 372314
rect 500924 372260 500959 372280
rect 500993 372260 501023 372294
rect 500924 372224 501023 372260
rect 500924 372190 500944 372224
rect 500978 372204 501023 372224
rect 500924 372170 500959 372190
rect 500993 372170 501023 372204
rect 500924 372134 501023 372170
rect 500924 372100 500944 372134
rect 500978 372114 501023 372134
rect 500924 372080 500959 372100
rect 500993 372080 501023 372114
rect 500924 372044 501023 372080
rect 500924 372010 500944 372044
rect 500978 372024 501023 372044
rect 500924 371990 500959 372010
rect 500993 371990 501023 372024
rect 501087 372962 502049 372981
rect 501087 372960 501163 372962
rect 501087 372926 501104 372960
rect 501138 372928 501163 372960
rect 501197 372928 501253 372962
rect 501287 372928 501343 372962
rect 501377 372928 501433 372962
rect 501467 372928 501523 372962
rect 501557 372928 501613 372962
rect 501647 372928 501703 372962
rect 501737 372928 501793 372962
rect 501827 372928 501883 372962
rect 501917 372928 502049 372962
rect 501138 372926 502049 372928
rect 501087 372909 502049 372926
rect 501087 372870 501159 372909
rect 501087 372836 501104 372870
rect 501138 372850 501159 372870
rect 501087 372816 501106 372836
rect 501140 372816 501159 372850
rect 501977 372884 502049 372909
rect 501977 372850 501996 372884
rect 502030 372850 502049 372884
rect 501087 372780 501159 372816
rect 501087 372746 501104 372780
rect 501138 372760 501159 372780
rect 501087 372726 501106 372746
rect 501140 372726 501159 372760
rect 501087 372690 501159 372726
rect 501087 372656 501104 372690
rect 501138 372670 501159 372690
rect 501087 372636 501106 372656
rect 501140 372636 501159 372670
rect 501087 372600 501159 372636
rect 501087 372566 501104 372600
rect 501138 372580 501159 372600
rect 501087 372546 501106 372566
rect 501140 372546 501159 372580
rect 501087 372510 501159 372546
rect 501087 372476 501104 372510
rect 501138 372490 501159 372510
rect 501087 372456 501106 372476
rect 501140 372456 501159 372490
rect 501087 372420 501159 372456
rect 501087 372386 501104 372420
rect 501138 372400 501159 372420
rect 501087 372366 501106 372386
rect 501140 372366 501159 372400
rect 501087 372330 501159 372366
rect 501087 372296 501104 372330
rect 501138 372310 501159 372330
rect 501087 372276 501106 372296
rect 501140 372276 501159 372310
rect 501087 372240 501159 372276
rect 501087 372206 501104 372240
rect 501138 372220 501159 372240
rect 501087 372186 501106 372206
rect 501140 372186 501159 372220
rect 501087 372150 501159 372186
rect 501221 372786 501915 372847
rect 501221 372752 501280 372786
rect 501314 372774 501370 372786
rect 501342 372752 501370 372774
rect 501404 372774 501460 372786
rect 501404 372752 501408 372774
rect 501221 372740 501308 372752
rect 501342 372740 501408 372752
rect 501442 372752 501460 372774
rect 501494 372774 501550 372786
rect 501494 372752 501508 372774
rect 501442 372740 501508 372752
rect 501542 372752 501550 372774
rect 501584 372774 501640 372786
rect 501674 372774 501730 372786
rect 501764 372774 501820 372786
rect 501584 372752 501608 372774
rect 501674 372752 501708 372774
rect 501764 372752 501808 372774
rect 501854 372752 501915 372786
rect 501542 372740 501608 372752
rect 501642 372740 501708 372752
rect 501742 372740 501808 372752
rect 501842 372740 501915 372752
rect 501221 372696 501915 372740
rect 501221 372662 501280 372696
rect 501314 372674 501370 372696
rect 501342 372662 501370 372674
rect 501404 372674 501460 372696
rect 501404 372662 501408 372674
rect 501221 372640 501308 372662
rect 501342 372640 501408 372662
rect 501442 372662 501460 372674
rect 501494 372674 501550 372696
rect 501494 372662 501508 372674
rect 501442 372640 501508 372662
rect 501542 372662 501550 372674
rect 501584 372674 501640 372696
rect 501674 372674 501730 372696
rect 501764 372674 501820 372696
rect 501584 372662 501608 372674
rect 501674 372662 501708 372674
rect 501764 372662 501808 372674
rect 501854 372662 501915 372696
rect 501542 372640 501608 372662
rect 501642 372640 501708 372662
rect 501742 372640 501808 372662
rect 501842 372640 501915 372662
rect 501221 372606 501915 372640
rect 501221 372572 501280 372606
rect 501314 372574 501370 372606
rect 501342 372572 501370 372574
rect 501404 372574 501460 372606
rect 501404 372572 501408 372574
rect 501221 372540 501308 372572
rect 501342 372540 501408 372572
rect 501442 372572 501460 372574
rect 501494 372574 501550 372606
rect 501494 372572 501508 372574
rect 501442 372540 501508 372572
rect 501542 372572 501550 372574
rect 501584 372574 501640 372606
rect 501674 372574 501730 372606
rect 501764 372574 501820 372606
rect 501584 372572 501608 372574
rect 501674 372572 501708 372574
rect 501764 372572 501808 372574
rect 501854 372572 501915 372606
rect 501542 372540 501608 372572
rect 501642 372540 501708 372572
rect 501742 372540 501808 372572
rect 501842 372540 501915 372572
rect 501221 372516 501915 372540
rect 501221 372482 501280 372516
rect 501314 372482 501370 372516
rect 501404 372482 501460 372516
rect 501494 372482 501550 372516
rect 501584 372482 501640 372516
rect 501674 372482 501730 372516
rect 501764 372482 501820 372516
rect 501854 372482 501915 372516
rect 501221 372474 501915 372482
rect 501221 372440 501308 372474
rect 501342 372440 501408 372474
rect 501442 372440 501508 372474
rect 501542 372440 501608 372474
rect 501642 372440 501708 372474
rect 501742 372440 501808 372474
rect 501842 372440 501915 372474
rect 501221 372426 501915 372440
rect 501221 372392 501280 372426
rect 501314 372392 501370 372426
rect 501404 372392 501460 372426
rect 501494 372392 501550 372426
rect 501584 372392 501640 372426
rect 501674 372392 501730 372426
rect 501764 372392 501820 372426
rect 501854 372392 501915 372426
rect 501221 372374 501915 372392
rect 501221 372340 501308 372374
rect 501342 372340 501408 372374
rect 501442 372340 501508 372374
rect 501542 372340 501608 372374
rect 501642 372340 501708 372374
rect 501742 372340 501808 372374
rect 501842 372340 501915 372374
rect 501221 372336 501915 372340
rect 501221 372302 501280 372336
rect 501314 372302 501370 372336
rect 501404 372302 501460 372336
rect 501494 372302 501550 372336
rect 501584 372302 501640 372336
rect 501674 372302 501730 372336
rect 501764 372302 501820 372336
rect 501854 372302 501915 372336
rect 501221 372274 501915 372302
rect 501221 372246 501308 372274
rect 501342 372246 501408 372274
rect 501221 372212 501280 372246
rect 501342 372240 501370 372246
rect 501314 372212 501370 372240
rect 501404 372240 501408 372246
rect 501442 372246 501508 372274
rect 501442 372240 501460 372246
rect 501404 372212 501460 372240
rect 501494 372240 501508 372246
rect 501542 372246 501608 372274
rect 501642 372246 501708 372274
rect 501742 372246 501808 372274
rect 501842 372246 501915 372274
rect 501542 372240 501550 372246
rect 501494 372212 501550 372240
rect 501584 372240 501608 372246
rect 501674 372240 501708 372246
rect 501764 372240 501808 372246
rect 501584 372212 501640 372240
rect 501674 372212 501730 372240
rect 501764 372212 501820 372240
rect 501854 372212 501915 372246
rect 501221 372153 501915 372212
rect 501977 372794 502049 372850
rect 501977 372760 501996 372794
rect 502030 372760 502049 372794
rect 501977 372704 502049 372760
rect 501977 372670 501996 372704
rect 502030 372670 502049 372704
rect 501977 372614 502049 372670
rect 501977 372580 501996 372614
rect 502030 372580 502049 372614
rect 501977 372524 502049 372580
rect 501977 372490 501996 372524
rect 502030 372490 502049 372524
rect 501977 372434 502049 372490
rect 501977 372400 501996 372434
rect 502030 372400 502049 372434
rect 501977 372344 502049 372400
rect 501977 372310 501996 372344
rect 502030 372310 502049 372344
rect 501977 372254 502049 372310
rect 501977 372220 501996 372254
rect 502030 372220 502049 372254
rect 501977 372164 502049 372220
rect 501087 372116 501104 372150
rect 501138 372130 501159 372150
rect 501087 372096 501106 372116
rect 501140 372096 501159 372130
rect 501087 372091 501159 372096
rect 501977 372130 501996 372164
rect 502030 372130 502049 372164
rect 501977 372091 502049 372130
rect 501087 372072 502049 372091
rect 501087 372060 501182 372072
rect 501087 372026 501104 372060
rect 501138 372038 501182 372060
rect 501216 372038 501272 372072
rect 501306 372038 501362 372072
rect 501396 372038 501452 372072
rect 501486 372038 501542 372072
rect 501576 372038 501632 372072
rect 501666 372038 501722 372072
rect 501756 372038 501812 372072
rect 501846 372038 501902 372072
rect 501936 372038 502049 372072
rect 501138 372026 502049 372038
rect 501087 372019 502049 372026
rect 502113 372980 502146 373014
rect 502180 372980 502212 373014
rect 502113 372924 502212 372980
rect 502113 372890 502146 372924
rect 502180 372890 502212 372924
rect 502113 372834 502212 372890
rect 502113 372800 502146 372834
rect 502180 372800 502212 372834
rect 502113 372744 502212 372800
rect 502113 372710 502146 372744
rect 502180 372710 502212 372744
rect 502113 372654 502212 372710
rect 502113 372620 502146 372654
rect 502180 372620 502212 372654
rect 502113 372564 502212 372620
rect 502113 372530 502146 372564
rect 502180 372530 502212 372564
rect 502113 372474 502212 372530
rect 502113 372440 502146 372474
rect 502180 372440 502212 372474
rect 502113 372384 502212 372440
rect 502113 372350 502146 372384
rect 502180 372350 502212 372384
rect 502113 372294 502212 372350
rect 502113 372260 502146 372294
rect 502180 372260 502212 372294
rect 502113 372204 502212 372260
rect 502113 372170 502146 372204
rect 502180 372170 502212 372204
rect 502113 372114 502212 372170
rect 502113 372080 502146 372114
rect 502180 372080 502212 372114
rect 502113 372024 502212 372080
rect 500924 371955 501023 371990
rect 502113 371990 502146 372024
rect 502180 371990 502212 372024
rect 502113 371955 502212 371990
rect 500924 371954 502212 371955
rect 500924 371920 500944 371954
rect 500978 371923 502212 371954
rect 500978 371920 500982 371923
rect 500924 371889 500982 371920
rect 501016 371889 501072 371923
rect 501106 371889 501162 371923
rect 501196 371889 501252 371923
rect 501286 371889 501342 371923
rect 501376 371889 501432 371923
rect 501466 371889 501522 371923
rect 501556 371889 501612 371923
rect 501646 371889 501702 371923
rect 501736 371889 501792 371923
rect 501826 371889 501882 371923
rect 501916 371889 501972 371923
rect 502006 371889 502062 371923
rect 502096 371889 502212 371923
rect 500924 371784 502212 371889
rect 500924 371750 500944 371784
rect 500978 371770 502212 371784
rect 500978 371750 500982 371770
rect 500924 371736 500982 371750
rect 501016 371736 501072 371770
rect 501106 371736 501162 371770
rect 501196 371736 501252 371770
rect 501286 371736 501342 371770
rect 501376 371736 501432 371770
rect 501466 371736 501522 371770
rect 501556 371736 501612 371770
rect 501646 371736 501702 371770
rect 501736 371736 501792 371770
rect 501826 371736 501882 371770
rect 501916 371736 501972 371770
rect 502006 371736 502062 371770
rect 502096 371736 502212 371770
rect 500924 371705 502212 371736
rect 500924 371694 501023 371705
rect 500924 371660 500944 371694
rect 500978 371674 501023 371694
rect 500924 371640 500959 371660
rect 500993 371640 501023 371674
rect 502113 371674 502212 371705
rect 500924 371604 501023 371640
rect 500924 371570 500944 371604
rect 500978 371584 501023 371604
rect 500924 371550 500959 371570
rect 500993 371550 501023 371584
rect 500924 371514 501023 371550
rect 500924 371480 500944 371514
rect 500978 371494 501023 371514
rect 500924 371460 500959 371480
rect 500993 371460 501023 371494
rect 500924 371424 501023 371460
rect 500924 371390 500944 371424
rect 500978 371404 501023 371424
rect 500924 371370 500959 371390
rect 500993 371370 501023 371404
rect 500924 371334 501023 371370
rect 500924 371300 500944 371334
rect 500978 371314 501023 371334
rect 500924 371280 500959 371300
rect 500993 371280 501023 371314
rect 500924 371244 501023 371280
rect 500924 371210 500944 371244
rect 500978 371224 501023 371244
rect 500924 371190 500959 371210
rect 500993 371190 501023 371224
rect 500924 371154 501023 371190
rect 500924 371120 500944 371154
rect 500978 371134 501023 371154
rect 500924 371100 500959 371120
rect 500993 371100 501023 371134
rect 500924 371064 501023 371100
rect 500924 371030 500944 371064
rect 500978 371044 501023 371064
rect 500924 371010 500959 371030
rect 500993 371010 501023 371044
rect 500924 370974 501023 371010
rect 500924 370940 500944 370974
rect 500978 370954 501023 370974
rect 500924 370920 500959 370940
rect 500993 370920 501023 370954
rect 500924 370884 501023 370920
rect 500924 370850 500944 370884
rect 500978 370864 501023 370884
rect 500924 370830 500959 370850
rect 500993 370830 501023 370864
rect 500924 370794 501023 370830
rect 500924 370760 500944 370794
rect 500978 370774 501023 370794
rect 500924 370740 500959 370760
rect 500993 370740 501023 370774
rect 500924 370704 501023 370740
rect 500924 370670 500944 370704
rect 500978 370684 501023 370704
rect 500924 370650 500959 370670
rect 500993 370650 501023 370684
rect 501087 371622 502049 371641
rect 501087 371620 501163 371622
rect 501087 371586 501104 371620
rect 501138 371588 501163 371620
rect 501197 371588 501253 371622
rect 501287 371588 501343 371622
rect 501377 371588 501433 371622
rect 501467 371588 501523 371622
rect 501557 371588 501613 371622
rect 501647 371588 501703 371622
rect 501737 371588 501793 371622
rect 501827 371588 501883 371622
rect 501917 371588 502049 371622
rect 501138 371586 502049 371588
rect 501087 371569 502049 371586
rect 501087 371530 501159 371569
rect 501087 371496 501104 371530
rect 501138 371510 501159 371530
rect 501087 371476 501106 371496
rect 501140 371476 501159 371510
rect 501977 371544 502049 371569
rect 501977 371510 501996 371544
rect 502030 371510 502049 371544
rect 501087 371440 501159 371476
rect 501087 371406 501104 371440
rect 501138 371420 501159 371440
rect 501087 371386 501106 371406
rect 501140 371386 501159 371420
rect 501087 371350 501159 371386
rect 501087 371316 501104 371350
rect 501138 371330 501159 371350
rect 501087 371296 501106 371316
rect 501140 371296 501159 371330
rect 501087 371260 501159 371296
rect 501087 371226 501104 371260
rect 501138 371240 501159 371260
rect 501087 371206 501106 371226
rect 501140 371206 501159 371240
rect 501087 371170 501159 371206
rect 501087 371136 501104 371170
rect 501138 371150 501159 371170
rect 501087 371116 501106 371136
rect 501140 371116 501159 371150
rect 501087 371080 501159 371116
rect 501087 371046 501104 371080
rect 501138 371060 501159 371080
rect 501087 371026 501106 371046
rect 501140 371026 501159 371060
rect 501087 370990 501159 371026
rect 501087 370956 501104 370990
rect 501138 370970 501159 370990
rect 501087 370936 501106 370956
rect 501140 370936 501159 370970
rect 501087 370900 501159 370936
rect 501087 370866 501104 370900
rect 501138 370880 501159 370900
rect 501087 370846 501106 370866
rect 501140 370846 501159 370880
rect 501087 370810 501159 370846
rect 501221 371446 501915 371507
rect 501221 371412 501280 371446
rect 501314 371434 501370 371446
rect 501342 371412 501370 371434
rect 501404 371434 501460 371446
rect 501404 371412 501408 371434
rect 501221 371400 501308 371412
rect 501342 371400 501408 371412
rect 501442 371412 501460 371434
rect 501494 371434 501550 371446
rect 501494 371412 501508 371434
rect 501442 371400 501508 371412
rect 501542 371412 501550 371434
rect 501584 371434 501640 371446
rect 501674 371434 501730 371446
rect 501764 371434 501820 371446
rect 501584 371412 501608 371434
rect 501674 371412 501708 371434
rect 501764 371412 501808 371434
rect 501854 371412 501915 371446
rect 501542 371400 501608 371412
rect 501642 371400 501708 371412
rect 501742 371400 501808 371412
rect 501842 371400 501915 371412
rect 501221 371356 501915 371400
rect 501221 371322 501280 371356
rect 501314 371334 501370 371356
rect 501342 371322 501370 371334
rect 501404 371334 501460 371356
rect 501404 371322 501408 371334
rect 501221 371300 501308 371322
rect 501342 371300 501408 371322
rect 501442 371322 501460 371334
rect 501494 371334 501550 371356
rect 501494 371322 501508 371334
rect 501442 371300 501508 371322
rect 501542 371322 501550 371334
rect 501584 371334 501640 371356
rect 501674 371334 501730 371356
rect 501764 371334 501820 371356
rect 501584 371322 501608 371334
rect 501674 371322 501708 371334
rect 501764 371322 501808 371334
rect 501854 371322 501915 371356
rect 501542 371300 501608 371322
rect 501642 371300 501708 371322
rect 501742 371300 501808 371322
rect 501842 371300 501915 371322
rect 501221 371266 501915 371300
rect 501221 371232 501280 371266
rect 501314 371234 501370 371266
rect 501342 371232 501370 371234
rect 501404 371234 501460 371266
rect 501404 371232 501408 371234
rect 501221 371200 501308 371232
rect 501342 371200 501408 371232
rect 501442 371232 501460 371234
rect 501494 371234 501550 371266
rect 501494 371232 501508 371234
rect 501442 371200 501508 371232
rect 501542 371232 501550 371234
rect 501584 371234 501640 371266
rect 501674 371234 501730 371266
rect 501764 371234 501820 371266
rect 501584 371232 501608 371234
rect 501674 371232 501708 371234
rect 501764 371232 501808 371234
rect 501854 371232 501915 371266
rect 501542 371200 501608 371232
rect 501642 371200 501708 371232
rect 501742 371200 501808 371232
rect 501842 371200 501915 371232
rect 501221 371176 501915 371200
rect 501221 371142 501280 371176
rect 501314 371142 501370 371176
rect 501404 371142 501460 371176
rect 501494 371142 501550 371176
rect 501584 371142 501640 371176
rect 501674 371142 501730 371176
rect 501764 371142 501820 371176
rect 501854 371142 501915 371176
rect 501221 371134 501915 371142
rect 501221 371100 501308 371134
rect 501342 371100 501408 371134
rect 501442 371100 501508 371134
rect 501542 371100 501608 371134
rect 501642 371100 501708 371134
rect 501742 371100 501808 371134
rect 501842 371100 501915 371134
rect 501221 371086 501915 371100
rect 501221 371052 501280 371086
rect 501314 371052 501370 371086
rect 501404 371052 501460 371086
rect 501494 371052 501550 371086
rect 501584 371052 501640 371086
rect 501674 371052 501730 371086
rect 501764 371052 501820 371086
rect 501854 371052 501915 371086
rect 501221 371034 501915 371052
rect 501221 371000 501308 371034
rect 501342 371000 501408 371034
rect 501442 371000 501508 371034
rect 501542 371000 501608 371034
rect 501642 371000 501708 371034
rect 501742 371000 501808 371034
rect 501842 371000 501915 371034
rect 501221 370996 501915 371000
rect 501221 370962 501280 370996
rect 501314 370962 501370 370996
rect 501404 370962 501460 370996
rect 501494 370962 501550 370996
rect 501584 370962 501640 370996
rect 501674 370962 501730 370996
rect 501764 370962 501820 370996
rect 501854 370962 501915 370996
rect 501221 370934 501915 370962
rect 501221 370906 501308 370934
rect 501342 370906 501408 370934
rect 501221 370872 501280 370906
rect 501342 370900 501370 370906
rect 501314 370872 501370 370900
rect 501404 370900 501408 370906
rect 501442 370906 501508 370934
rect 501442 370900 501460 370906
rect 501404 370872 501460 370900
rect 501494 370900 501508 370906
rect 501542 370906 501608 370934
rect 501642 370906 501708 370934
rect 501742 370906 501808 370934
rect 501842 370906 501915 370934
rect 501542 370900 501550 370906
rect 501494 370872 501550 370900
rect 501584 370900 501608 370906
rect 501674 370900 501708 370906
rect 501764 370900 501808 370906
rect 501584 370872 501640 370900
rect 501674 370872 501730 370900
rect 501764 370872 501820 370900
rect 501854 370872 501915 370906
rect 501221 370813 501915 370872
rect 501977 371454 502049 371510
rect 501977 371420 501996 371454
rect 502030 371420 502049 371454
rect 501977 371364 502049 371420
rect 501977 371330 501996 371364
rect 502030 371330 502049 371364
rect 501977 371274 502049 371330
rect 501977 371240 501996 371274
rect 502030 371240 502049 371274
rect 501977 371184 502049 371240
rect 501977 371150 501996 371184
rect 502030 371150 502049 371184
rect 501977 371094 502049 371150
rect 501977 371060 501996 371094
rect 502030 371060 502049 371094
rect 501977 371004 502049 371060
rect 501977 370970 501996 371004
rect 502030 370970 502049 371004
rect 501977 370914 502049 370970
rect 501977 370880 501996 370914
rect 502030 370880 502049 370914
rect 501977 370824 502049 370880
rect 501087 370776 501104 370810
rect 501138 370790 501159 370810
rect 501087 370756 501106 370776
rect 501140 370756 501159 370790
rect 501087 370751 501159 370756
rect 501977 370790 501996 370824
rect 502030 370790 502049 370824
rect 501977 370751 502049 370790
rect 501087 370732 502049 370751
rect 501087 370720 501182 370732
rect 501087 370686 501104 370720
rect 501138 370698 501182 370720
rect 501216 370698 501272 370732
rect 501306 370698 501362 370732
rect 501396 370698 501452 370732
rect 501486 370698 501542 370732
rect 501576 370698 501632 370732
rect 501666 370698 501722 370732
rect 501756 370698 501812 370732
rect 501846 370698 501902 370732
rect 501936 370698 502049 370732
rect 501138 370686 502049 370698
rect 501087 370679 502049 370686
rect 502113 371640 502146 371674
rect 502180 371640 502212 371674
rect 502113 371584 502212 371640
rect 502113 371550 502146 371584
rect 502180 371550 502212 371584
rect 502113 371494 502212 371550
rect 502113 371460 502146 371494
rect 502180 371460 502212 371494
rect 502113 371404 502212 371460
rect 502113 371370 502146 371404
rect 502180 371370 502212 371404
rect 502113 371314 502212 371370
rect 502113 371280 502146 371314
rect 502180 371280 502212 371314
rect 502113 371224 502212 371280
rect 502113 371190 502146 371224
rect 502180 371190 502212 371224
rect 502113 371134 502212 371190
rect 502113 371100 502146 371134
rect 502180 371100 502212 371134
rect 502113 371044 502212 371100
rect 502113 371010 502146 371044
rect 502180 371010 502212 371044
rect 502113 370954 502212 371010
rect 502113 370920 502146 370954
rect 502180 370920 502212 370954
rect 502113 370864 502212 370920
rect 502113 370830 502146 370864
rect 502180 370830 502212 370864
rect 502113 370774 502212 370830
rect 502113 370740 502146 370774
rect 502180 370740 502212 370774
rect 502113 370684 502212 370740
rect 500924 370615 501023 370650
rect 502113 370650 502146 370684
rect 502180 370650 502212 370684
rect 502113 370615 502212 370650
rect 500924 370614 502212 370615
rect 500924 370580 500944 370614
rect 500978 370583 502212 370614
rect 500978 370580 500982 370583
rect 500924 370549 500982 370580
rect 501016 370549 501072 370583
rect 501106 370549 501162 370583
rect 501196 370549 501252 370583
rect 501286 370549 501342 370583
rect 501376 370549 501432 370583
rect 501466 370549 501522 370583
rect 501556 370549 501612 370583
rect 501646 370549 501702 370583
rect 501736 370549 501792 370583
rect 501826 370549 501882 370583
rect 501916 370549 501972 370583
rect 502006 370549 502062 370583
rect 502096 370549 502212 370583
rect 500924 370444 502212 370549
rect 500924 370410 500944 370444
rect 500978 370430 502212 370444
rect 500978 370410 500982 370430
rect 500924 370396 500982 370410
rect 501016 370396 501072 370430
rect 501106 370396 501162 370430
rect 501196 370396 501252 370430
rect 501286 370396 501342 370430
rect 501376 370396 501432 370430
rect 501466 370396 501522 370430
rect 501556 370396 501612 370430
rect 501646 370396 501702 370430
rect 501736 370396 501792 370430
rect 501826 370396 501882 370430
rect 501916 370396 501972 370430
rect 502006 370396 502062 370430
rect 502096 370396 502212 370430
rect 500924 370365 502212 370396
rect 500924 370354 501023 370365
rect 500924 370320 500944 370354
rect 500978 370334 501023 370354
rect 500924 370300 500959 370320
rect 500993 370300 501023 370334
rect 502113 370334 502212 370365
rect 500924 370264 501023 370300
rect 500924 370230 500944 370264
rect 500978 370244 501023 370264
rect 500924 370210 500959 370230
rect 500993 370210 501023 370244
rect 500924 370174 501023 370210
rect 500924 370140 500944 370174
rect 500978 370154 501023 370174
rect 500924 370120 500959 370140
rect 500993 370120 501023 370154
rect 500924 370084 501023 370120
rect 500924 370050 500944 370084
rect 500978 370064 501023 370084
rect 500924 370030 500959 370050
rect 500993 370030 501023 370064
rect 500924 369994 501023 370030
rect 500924 369960 500944 369994
rect 500978 369974 501023 369994
rect 500924 369940 500959 369960
rect 500993 369940 501023 369974
rect 500924 369904 501023 369940
rect 500924 369870 500944 369904
rect 500978 369884 501023 369904
rect 500924 369850 500959 369870
rect 500993 369850 501023 369884
rect 500924 369814 501023 369850
rect 500924 369780 500944 369814
rect 500978 369794 501023 369814
rect 500924 369760 500959 369780
rect 500993 369760 501023 369794
rect 500924 369724 501023 369760
rect 500924 369690 500944 369724
rect 500978 369704 501023 369724
rect 500924 369670 500959 369690
rect 500993 369670 501023 369704
rect 500924 369634 501023 369670
rect 500924 369600 500944 369634
rect 500978 369614 501023 369634
rect 500924 369580 500959 369600
rect 500993 369580 501023 369614
rect 500924 369544 501023 369580
rect 500924 369510 500944 369544
rect 500978 369524 501023 369544
rect 500924 369490 500959 369510
rect 500993 369490 501023 369524
rect 500924 369454 501023 369490
rect 500924 369420 500944 369454
rect 500978 369434 501023 369454
rect 500924 369400 500959 369420
rect 500993 369400 501023 369434
rect 500924 369364 501023 369400
rect 500924 369330 500944 369364
rect 500978 369344 501023 369364
rect 500924 369310 500959 369330
rect 500993 369310 501023 369344
rect 501087 370282 502049 370301
rect 501087 370280 501163 370282
rect 501087 370246 501104 370280
rect 501138 370248 501163 370280
rect 501197 370248 501253 370282
rect 501287 370248 501343 370282
rect 501377 370248 501433 370282
rect 501467 370248 501523 370282
rect 501557 370248 501613 370282
rect 501647 370248 501703 370282
rect 501737 370248 501793 370282
rect 501827 370248 501883 370282
rect 501917 370248 502049 370282
rect 501138 370246 502049 370248
rect 501087 370229 502049 370246
rect 501087 370190 501159 370229
rect 501087 370156 501104 370190
rect 501138 370170 501159 370190
rect 501087 370136 501106 370156
rect 501140 370136 501159 370170
rect 501977 370204 502049 370229
rect 501977 370170 501996 370204
rect 502030 370170 502049 370204
rect 501087 370100 501159 370136
rect 501087 370066 501104 370100
rect 501138 370080 501159 370100
rect 501087 370046 501106 370066
rect 501140 370046 501159 370080
rect 501087 370010 501159 370046
rect 501087 369976 501104 370010
rect 501138 369990 501159 370010
rect 501087 369956 501106 369976
rect 501140 369956 501159 369990
rect 501087 369920 501159 369956
rect 501087 369886 501104 369920
rect 501138 369900 501159 369920
rect 501087 369866 501106 369886
rect 501140 369866 501159 369900
rect 501087 369830 501159 369866
rect 501087 369796 501104 369830
rect 501138 369810 501159 369830
rect 501087 369776 501106 369796
rect 501140 369776 501159 369810
rect 501087 369740 501159 369776
rect 501087 369706 501104 369740
rect 501138 369720 501159 369740
rect 501087 369686 501106 369706
rect 501140 369686 501159 369720
rect 501087 369650 501159 369686
rect 501087 369616 501104 369650
rect 501138 369630 501159 369650
rect 501087 369596 501106 369616
rect 501140 369596 501159 369630
rect 501087 369560 501159 369596
rect 501087 369526 501104 369560
rect 501138 369540 501159 369560
rect 501087 369506 501106 369526
rect 501140 369506 501159 369540
rect 501087 369470 501159 369506
rect 501221 370106 501915 370167
rect 501221 370072 501280 370106
rect 501314 370094 501370 370106
rect 501342 370072 501370 370094
rect 501404 370094 501460 370106
rect 501404 370072 501408 370094
rect 501221 370060 501308 370072
rect 501342 370060 501408 370072
rect 501442 370072 501460 370094
rect 501494 370094 501550 370106
rect 501494 370072 501508 370094
rect 501442 370060 501508 370072
rect 501542 370072 501550 370094
rect 501584 370094 501640 370106
rect 501674 370094 501730 370106
rect 501764 370094 501820 370106
rect 501584 370072 501608 370094
rect 501674 370072 501708 370094
rect 501764 370072 501808 370094
rect 501854 370072 501915 370106
rect 501542 370060 501608 370072
rect 501642 370060 501708 370072
rect 501742 370060 501808 370072
rect 501842 370060 501915 370072
rect 501221 370016 501915 370060
rect 501221 369982 501280 370016
rect 501314 369994 501370 370016
rect 501342 369982 501370 369994
rect 501404 369994 501460 370016
rect 501404 369982 501408 369994
rect 501221 369960 501308 369982
rect 501342 369960 501408 369982
rect 501442 369982 501460 369994
rect 501494 369994 501550 370016
rect 501494 369982 501508 369994
rect 501442 369960 501508 369982
rect 501542 369982 501550 369994
rect 501584 369994 501640 370016
rect 501674 369994 501730 370016
rect 501764 369994 501820 370016
rect 501584 369982 501608 369994
rect 501674 369982 501708 369994
rect 501764 369982 501808 369994
rect 501854 369982 501915 370016
rect 501542 369960 501608 369982
rect 501642 369960 501708 369982
rect 501742 369960 501808 369982
rect 501842 369960 501915 369982
rect 501221 369926 501915 369960
rect 501221 369892 501280 369926
rect 501314 369894 501370 369926
rect 501342 369892 501370 369894
rect 501404 369894 501460 369926
rect 501404 369892 501408 369894
rect 501221 369860 501308 369892
rect 501342 369860 501408 369892
rect 501442 369892 501460 369894
rect 501494 369894 501550 369926
rect 501494 369892 501508 369894
rect 501442 369860 501508 369892
rect 501542 369892 501550 369894
rect 501584 369894 501640 369926
rect 501674 369894 501730 369926
rect 501764 369894 501820 369926
rect 501584 369892 501608 369894
rect 501674 369892 501708 369894
rect 501764 369892 501808 369894
rect 501854 369892 501915 369926
rect 501542 369860 501608 369892
rect 501642 369860 501708 369892
rect 501742 369860 501808 369892
rect 501842 369860 501915 369892
rect 501221 369836 501915 369860
rect 501221 369802 501280 369836
rect 501314 369802 501370 369836
rect 501404 369802 501460 369836
rect 501494 369802 501550 369836
rect 501584 369802 501640 369836
rect 501674 369802 501730 369836
rect 501764 369802 501820 369836
rect 501854 369802 501915 369836
rect 501221 369794 501915 369802
rect 501221 369760 501308 369794
rect 501342 369760 501408 369794
rect 501442 369760 501508 369794
rect 501542 369760 501608 369794
rect 501642 369760 501708 369794
rect 501742 369760 501808 369794
rect 501842 369760 501915 369794
rect 501221 369746 501915 369760
rect 501221 369712 501280 369746
rect 501314 369712 501370 369746
rect 501404 369712 501460 369746
rect 501494 369712 501550 369746
rect 501584 369712 501640 369746
rect 501674 369712 501730 369746
rect 501764 369712 501820 369746
rect 501854 369712 501915 369746
rect 501221 369694 501915 369712
rect 501221 369660 501308 369694
rect 501342 369660 501408 369694
rect 501442 369660 501508 369694
rect 501542 369660 501608 369694
rect 501642 369660 501708 369694
rect 501742 369660 501808 369694
rect 501842 369660 501915 369694
rect 501221 369656 501915 369660
rect 501221 369622 501280 369656
rect 501314 369622 501370 369656
rect 501404 369622 501460 369656
rect 501494 369622 501550 369656
rect 501584 369622 501640 369656
rect 501674 369622 501730 369656
rect 501764 369622 501820 369656
rect 501854 369622 501915 369656
rect 501221 369594 501915 369622
rect 501221 369566 501308 369594
rect 501342 369566 501408 369594
rect 501221 369532 501280 369566
rect 501342 369560 501370 369566
rect 501314 369532 501370 369560
rect 501404 369560 501408 369566
rect 501442 369566 501508 369594
rect 501442 369560 501460 369566
rect 501404 369532 501460 369560
rect 501494 369560 501508 369566
rect 501542 369566 501608 369594
rect 501642 369566 501708 369594
rect 501742 369566 501808 369594
rect 501842 369566 501915 369594
rect 501542 369560 501550 369566
rect 501494 369532 501550 369560
rect 501584 369560 501608 369566
rect 501674 369560 501708 369566
rect 501764 369560 501808 369566
rect 501584 369532 501640 369560
rect 501674 369532 501730 369560
rect 501764 369532 501820 369560
rect 501854 369532 501915 369566
rect 501221 369473 501915 369532
rect 501977 370114 502049 370170
rect 501977 370080 501996 370114
rect 502030 370080 502049 370114
rect 501977 370024 502049 370080
rect 501977 369990 501996 370024
rect 502030 369990 502049 370024
rect 501977 369934 502049 369990
rect 501977 369900 501996 369934
rect 502030 369900 502049 369934
rect 501977 369844 502049 369900
rect 501977 369810 501996 369844
rect 502030 369810 502049 369844
rect 501977 369754 502049 369810
rect 501977 369720 501996 369754
rect 502030 369720 502049 369754
rect 501977 369664 502049 369720
rect 501977 369630 501996 369664
rect 502030 369630 502049 369664
rect 501977 369574 502049 369630
rect 501977 369540 501996 369574
rect 502030 369540 502049 369574
rect 501977 369484 502049 369540
rect 501087 369436 501104 369470
rect 501138 369450 501159 369470
rect 501087 369416 501106 369436
rect 501140 369416 501159 369450
rect 501087 369411 501159 369416
rect 501977 369450 501996 369484
rect 502030 369450 502049 369484
rect 501977 369411 502049 369450
rect 501087 369392 502049 369411
rect 501087 369380 501182 369392
rect 501087 369346 501104 369380
rect 501138 369358 501182 369380
rect 501216 369358 501272 369392
rect 501306 369358 501362 369392
rect 501396 369358 501452 369392
rect 501486 369358 501542 369392
rect 501576 369358 501632 369392
rect 501666 369358 501722 369392
rect 501756 369358 501812 369392
rect 501846 369358 501902 369392
rect 501936 369358 502049 369392
rect 501138 369346 502049 369358
rect 501087 369339 502049 369346
rect 502113 370300 502146 370334
rect 502180 370300 502212 370334
rect 502113 370244 502212 370300
rect 502113 370210 502146 370244
rect 502180 370210 502212 370244
rect 502113 370154 502212 370210
rect 502113 370120 502146 370154
rect 502180 370120 502212 370154
rect 502113 370064 502212 370120
rect 502113 370030 502146 370064
rect 502180 370030 502212 370064
rect 502113 369974 502212 370030
rect 502113 369940 502146 369974
rect 502180 369940 502212 369974
rect 502113 369884 502212 369940
rect 502113 369850 502146 369884
rect 502180 369850 502212 369884
rect 502113 369794 502212 369850
rect 502113 369760 502146 369794
rect 502180 369760 502212 369794
rect 502113 369704 502212 369760
rect 502113 369670 502146 369704
rect 502180 369670 502212 369704
rect 502113 369614 502212 369670
rect 502113 369580 502146 369614
rect 502180 369580 502212 369614
rect 502113 369524 502212 369580
rect 502113 369490 502146 369524
rect 502180 369490 502212 369524
rect 502113 369434 502212 369490
rect 502113 369400 502146 369434
rect 502180 369400 502212 369434
rect 502113 369344 502212 369400
rect 500924 369275 501023 369310
rect 502113 369310 502146 369344
rect 502180 369310 502212 369344
rect 502113 369275 502212 369310
rect 500924 369274 502212 369275
rect 500924 369240 500944 369274
rect 500978 369243 502212 369274
rect 500978 369240 500982 369243
rect 500924 369209 500982 369240
rect 501016 369209 501072 369243
rect 501106 369209 501162 369243
rect 501196 369209 501252 369243
rect 501286 369209 501342 369243
rect 501376 369209 501432 369243
rect 501466 369209 501522 369243
rect 501556 369209 501612 369243
rect 501646 369209 501702 369243
rect 501736 369209 501792 369243
rect 501826 369209 501882 369243
rect 501916 369209 501972 369243
rect 502006 369209 502062 369243
rect 502096 369209 502212 369243
rect 500924 369104 502212 369209
rect 500924 369070 500944 369104
rect 500978 369090 502212 369104
rect 500978 369070 500982 369090
rect 500924 369056 500982 369070
rect 501016 369056 501072 369090
rect 501106 369056 501162 369090
rect 501196 369056 501252 369090
rect 501286 369056 501342 369090
rect 501376 369056 501432 369090
rect 501466 369056 501522 369090
rect 501556 369056 501612 369090
rect 501646 369056 501702 369090
rect 501736 369056 501792 369090
rect 501826 369056 501882 369090
rect 501916 369056 501972 369090
rect 502006 369056 502062 369090
rect 502096 369056 502212 369090
rect 500924 369025 502212 369056
rect 500924 369014 501023 369025
rect 500924 368980 500944 369014
rect 500978 368994 501023 369014
rect 500924 368960 500959 368980
rect 500993 368960 501023 368994
rect 502113 368994 502212 369025
rect 500924 368924 501023 368960
rect 500924 368890 500944 368924
rect 500978 368904 501023 368924
rect 500924 368870 500959 368890
rect 500993 368870 501023 368904
rect 500924 368834 501023 368870
rect 500924 368800 500944 368834
rect 500978 368814 501023 368834
rect 500924 368780 500959 368800
rect 500993 368780 501023 368814
rect 500924 368744 501023 368780
rect 500924 368710 500944 368744
rect 500978 368724 501023 368744
rect 500924 368690 500959 368710
rect 500993 368690 501023 368724
rect 500924 368654 501023 368690
rect 500924 368620 500944 368654
rect 500978 368634 501023 368654
rect 500924 368600 500959 368620
rect 500993 368600 501023 368634
rect 500924 368564 501023 368600
rect 500924 368530 500944 368564
rect 500978 368544 501023 368564
rect 500924 368510 500959 368530
rect 500993 368510 501023 368544
rect 500924 368474 501023 368510
rect 500924 368440 500944 368474
rect 500978 368454 501023 368474
rect 500924 368420 500959 368440
rect 500993 368420 501023 368454
rect 500924 368384 501023 368420
rect 500924 368350 500944 368384
rect 500978 368364 501023 368384
rect 500924 368330 500959 368350
rect 500993 368330 501023 368364
rect 500924 368294 501023 368330
rect 500924 368260 500944 368294
rect 500978 368274 501023 368294
rect 500924 368240 500959 368260
rect 500993 368240 501023 368274
rect 500924 368204 501023 368240
rect 500924 368170 500944 368204
rect 500978 368184 501023 368204
rect 500924 368150 500959 368170
rect 500993 368150 501023 368184
rect 500924 368114 501023 368150
rect 500924 368080 500944 368114
rect 500978 368094 501023 368114
rect 500924 368060 500959 368080
rect 500993 368060 501023 368094
rect 500924 368024 501023 368060
rect 500924 367990 500944 368024
rect 500978 368004 501023 368024
rect 500924 367970 500959 367990
rect 500993 367970 501023 368004
rect 501087 368942 502049 368961
rect 501087 368940 501163 368942
rect 501087 368906 501104 368940
rect 501138 368908 501163 368940
rect 501197 368908 501253 368942
rect 501287 368908 501343 368942
rect 501377 368908 501433 368942
rect 501467 368908 501523 368942
rect 501557 368908 501613 368942
rect 501647 368908 501703 368942
rect 501737 368908 501793 368942
rect 501827 368908 501883 368942
rect 501917 368908 502049 368942
rect 501138 368906 502049 368908
rect 501087 368889 502049 368906
rect 501087 368850 501159 368889
rect 501087 368816 501104 368850
rect 501138 368830 501159 368850
rect 501087 368796 501106 368816
rect 501140 368796 501159 368830
rect 501977 368864 502049 368889
rect 501977 368830 501996 368864
rect 502030 368830 502049 368864
rect 501087 368760 501159 368796
rect 501087 368726 501104 368760
rect 501138 368740 501159 368760
rect 501087 368706 501106 368726
rect 501140 368706 501159 368740
rect 501087 368670 501159 368706
rect 501087 368636 501104 368670
rect 501138 368650 501159 368670
rect 501087 368616 501106 368636
rect 501140 368616 501159 368650
rect 501087 368580 501159 368616
rect 501087 368546 501104 368580
rect 501138 368560 501159 368580
rect 501087 368526 501106 368546
rect 501140 368526 501159 368560
rect 501087 368490 501159 368526
rect 501087 368456 501104 368490
rect 501138 368470 501159 368490
rect 501087 368436 501106 368456
rect 501140 368436 501159 368470
rect 501087 368400 501159 368436
rect 501087 368366 501104 368400
rect 501138 368380 501159 368400
rect 501087 368346 501106 368366
rect 501140 368346 501159 368380
rect 501087 368310 501159 368346
rect 501087 368276 501104 368310
rect 501138 368290 501159 368310
rect 501087 368256 501106 368276
rect 501140 368256 501159 368290
rect 501087 368220 501159 368256
rect 501087 368186 501104 368220
rect 501138 368200 501159 368220
rect 501087 368166 501106 368186
rect 501140 368166 501159 368200
rect 501087 368130 501159 368166
rect 501221 368766 501915 368827
rect 501221 368732 501280 368766
rect 501314 368754 501370 368766
rect 501342 368732 501370 368754
rect 501404 368754 501460 368766
rect 501404 368732 501408 368754
rect 501221 368720 501308 368732
rect 501342 368720 501408 368732
rect 501442 368732 501460 368754
rect 501494 368754 501550 368766
rect 501494 368732 501508 368754
rect 501442 368720 501508 368732
rect 501542 368732 501550 368754
rect 501584 368754 501640 368766
rect 501674 368754 501730 368766
rect 501764 368754 501820 368766
rect 501584 368732 501608 368754
rect 501674 368732 501708 368754
rect 501764 368732 501808 368754
rect 501854 368732 501915 368766
rect 501542 368720 501608 368732
rect 501642 368720 501708 368732
rect 501742 368720 501808 368732
rect 501842 368720 501915 368732
rect 501221 368676 501915 368720
rect 501221 368642 501280 368676
rect 501314 368654 501370 368676
rect 501342 368642 501370 368654
rect 501404 368654 501460 368676
rect 501404 368642 501408 368654
rect 501221 368620 501308 368642
rect 501342 368620 501408 368642
rect 501442 368642 501460 368654
rect 501494 368654 501550 368676
rect 501494 368642 501508 368654
rect 501442 368620 501508 368642
rect 501542 368642 501550 368654
rect 501584 368654 501640 368676
rect 501674 368654 501730 368676
rect 501764 368654 501820 368676
rect 501584 368642 501608 368654
rect 501674 368642 501708 368654
rect 501764 368642 501808 368654
rect 501854 368642 501915 368676
rect 501542 368620 501608 368642
rect 501642 368620 501708 368642
rect 501742 368620 501808 368642
rect 501842 368620 501915 368642
rect 501221 368586 501915 368620
rect 501221 368552 501280 368586
rect 501314 368554 501370 368586
rect 501342 368552 501370 368554
rect 501404 368554 501460 368586
rect 501404 368552 501408 368554
rect 501221 368520 501308 368552
rect 501342 368520 501408 368552
rect 501442 368552 501460 368554
rect 501494 368554 501550 368586
rect 501494 368552 501508 368554
rect 501442 368520 501508 368552
rect 501542 368552 501550 368554
rect 501584 368554 501640 368586
rect 501674 368554 501730 368586
rect 501764 368554 501820 368586
rect 501584 368552 501608 368554
rect 501674 368552 501708 368554
rect 501764 368552 501808 368554
rect 501854 368552 501915 368586
rect 501542 368520 501608 368552
rect 501642 368520 501708 368552
rect 501742 368520 501808 368552
rect 501842 368520 501915 368552
rect 501221 368496 501915 368520
rect 501221 368462 501280 368496
rect 501314 368462 501370 368496
rect 501404 368462 501460 368496
rect 501494 368462 501550 368496
rect 501584 368462 501640 368496
rect 501674 368462 501730 368496
rect 501764 368462 501820 368496
rect 501854 368462 501915 368496
rect 501221 368454 501915 368462
rect 501221 368420 501308 368454
rect 501342 368420 501408 368454
rect 501442 368420 501508 368454
rect 501542 368420 501608 368454
rect 501642 368420 501708 368454
rect 501742 368420 501808 368454
rect 501842 368420 501915 368454
rect 501221 368406 501915 368420
rect 501221 368372 501280 368406
rect 501314 368372 501370 368406
rect 501404 368372 501460 368406
rect 501494 368372 501550 368406
rect 501584 368372 501640 368406
rect 501674 368372 501730 368406
rect 501764 368372 501820 368406
rect 501854 368372 501915 368406
rect 501221 368354 501915 368372
rect 501221 368320 501308 368354
rect 501342 368320 501408 368354
rect 501442 368320 501508 368354
rect 501542 368320 501608 368354
rect 501642 368320 501708 368354
rect 501742 368320 501808 368354
rect 501842 368320 501915 368354
rect 501221 368316 501915 368320
rect 501221 368282 501280 368316
rect 501314 368282 501370 368316
rect 501404 368282 501460 368316
rect 501494 368282 501550 368316
rect 501584 368282 501640 368316
rect 501674 368282 501730 368316
rect 501764 368282 501820 368316
rect 501854 368282 501915 368316
rect 501221 368254 501915 368282
rect 501221 368226 501308 368254
rect 501342 368226 501408 368254
rect 501221 368192 501280 368226
rect 501342 368220 501370 368226
rect 501314 368192 501370 368220
rect 501404 368220 501408 368226
rect 501442 368226 501508 368254
rect 501442 368220 501460 368226
rect 501404 368192 501460 368220
rect 501494 368220 501508 368226
rect 501542 368226 501608 368254
rect 501642 368226 501708 368254
rect 501742 368226 501808 368254
rect 501842 368226 501915 368254
rect 501542 368220 501550 368226
rect 501494 368192 501550 368220
rect 501584 368220 501608 368226
rect 501674 368220 501708 368226
rect 501764 368220 501808 368226
rect 501584 368192 501640 368220
rect 501674 368192 501730 368220
rect 501764 368192 501820 368220
rect 501854 368192 501915 368226
rect 501221 368133 501915 368192
rect 501977 368774 502049 368830
rect 501977 368740 501996 368774
rect 502030 368740 502049 368774
rect 501977 368684 502049 368740
rect 501977 368650 501996 368684
rect 502030 368650 502049 368684
rect 501977 368594 502049 368650
rect 501977 368560 501996 368594
rect 502030 368560 502049 368594
rect 501977 368504 502049 368560
rect 501977 368470 501996 368504
rect 502030 368470 502049 368504
rect 501977 368414 502049 368470
rect 501977 368380 501996 368414
rect 502030 368380 502049 368414
rect 501977 368324 502049 368380
rect 501977 368290 501996 368324
rect 502030 368290 502049 368324
rect 501977 368234 502049 368290
rect 501977 368200 501996 368234
rect 502030 368200 502049 368234
rect 501977 368144 502049 368200
rect 501087 368096 501104 368130
rect 501138 368110 501159 368130
rect 501087 368076 501106 368096
rect 501140 368076 501159 368110
rect 501087 368071 501159 368076
rect 501977 368110 501996 368144
rect 502030 368110 502049 368144
rect 501977 368071 502049 368110
rect 501087 368052 502049 368071
rect 501087 368040 501182 368052
rect 501087 368006 501104 368040
rect 501138 368018 501182 368040
rect 501216 368018 501272 368052
rect 501306 368018 501362 368052
rect 501396 368018 501452 368052
rect 501486 368018 501542 368052
rect 501576 368018 501632 368052
rect 501666 368018 501722 368052
rect 501756 368018 501812 368052
rect 501846 368018 501902 368052
rect 501936 368018 502049 368052
rect 501138 368006 502049 368018
rect 501087 367999 502049 368006
rect 502113 368960 502146 368994
rect 502180 368960 502212 368994
rect 502113 368904 502212 368960
rect 502113 368870 502146 368904
rect 502180 368870 502212 368904
rect 502113 368814 502212 368870
rect 502113 368780 502146 368814
rect 502180 368780 502212 368814
rect 502113 368724 502212 368780
rect 502113 368690 502146 368724
rect 502180 368690 502212 368724
rect 502113 368634 502212 368690
rect 502113 368600 502146 368634
rect 502180 368600 502212 368634
rect 502113 368544 502212 368600
rect 502113 368510 502146 368544
rect 502180 368510 502212 368544
rect 502113 368454 502212 368510
rect 502113 368420 502146 368454
rect 502180 368420 502212 368454
rect 502113 368364 502212 368420
rect 502113 368330 502146 368364
rect 502180 368330 502212 368364
rect 502113 368274 502212 368330
rect 502113 368240 502146 368274
rect 502180 368240 502212 368274
rect 502113 368184 502212 368240
rect 502113 368150 502146 368184
rect 502180 368150 502212 368184
rect 502113 368094 502212 368150
rect 502113 368060 502146 368094
rect 502180 368060 502212 368094
rect 502113 368004 502212 368060
rect 500924 367935 501023 367970
rect 502113 367970 502146 368004
rect 502180 367970 502212 368004
rect 502113 367935 502212 367970
rect 500924 367934 502212 367935
rect 500924 367900 500944 367934
rect 500978 367903 502212 367934
rect 500978 367900 500982 367903
rect 500924 367869 500982 367900
rect 501016 367869 501072 367903
rect 501106 367869 501162 367903
rect 501196 367869 501252 367903
rect 501286 367869 501342 367903
rect 501376 367869 501432 367903
rect 501466 367869 501522 367903
rect 501556 367869 501612 367903
rect 501646 367869 501702 367903
rect 501736 367869 501792 367903
rect 501826 367869 501882 367903
rect 501916 367869 501972 367903
rect 502006 367869 502062 367903
rect 502096 367869 502212 367903
rect 500924 367764 502212 367869
rect 500924 367730 500944 367764
rect 500978 367750 502212 367764
rect 500978 367730 500982 367750
rect 500924 367716 500982 367730
rect 501016 367716 501072 367750
rect 501106 367716 501162 367750
rect 501196 367716 501252 367750
rect 501286 367716 501342 367750
rect 501376 367716 501432 367750
rect 501466 367716 501522 367750
rect 501556 367716 501612 367750
rect 501646 367716 501702 367750
rect 501736 367716 501792 367750
rect 501826 367716 501882 367750
rect 501916 367716 501972 367750
rect 502006 367716 502062 367750
rect 502096 367716 502212 367750
rect 500924 367685 502212 367716
rect 500924 367674 501023 367685
rect 500924 367640 500944 367674
rect 500978 367654 501023 367674
rect 500924 367620 500959 367640
rect 500993 367620 501023 367654
rect 502113 367654 502212 367685
rect 500924 367584 501023 367620
rect 500924 367550 500944 367584
rect 500978 367564 501023 367584
rect 500924 367530 500959 367550
rect 500993 367530 501023 367564
rect 500924 367494 501023 367530
rect 500924 367460 500944 367494
rect 500978 367474 501023 367494
rect 500924 367440 500959 367460
rect 500993 367440 501023 367474
rect 500924 367404 501023 367440
rect 500924 367370 500944 367404
rect 500978 367384 501023 367404
rect 500924 367350 500959 367370
rect 500993 367350 501023 367384
rect 500924 367314 501023 367350
rect 500924 367280 500944 367314
rect 500978 367294 501023 367314
rect 500924 367260 500959 367280
rect 500993 367260 501023 367294
rect 500924 367224 501023 367260
rect 500924 367190 500944 367224
rect 500978 367204 501023 367224
rect 500924 367170 500959 367190
rect 500993 367170 501023 367204
rect 500924 367134 501023 367170
rect 500924 367100 500944 367134
rect 500978 367114 501023 367134
rect 500924 367080 500959 367100
rect 500993 367080 501023 367114
rect 500924 367044 501023 367080
rect 500924 367010 500944 367044
rect 500978 367024 501023 367044
rect 500924 366990 500959 367010
rect 500993 366990 501023 367024
rect 500924 366954 501023 366990
rect 500924 366920 500944 366954
rect 500978 366934 501023 366954
rect 500924 366900 500959 366920
rect 500993 366900 501023 366934
rect 500924 366864 501023 366900
rect 500924 366830 500944 366864
rect 500978 366844 501023 366864
rect 500924 366810 500959 366830
rect 500993 366810 501023 366844
rect 500924 366774 501023 366810
rect 500924 366740 500944 366774
rect 500978 366754 501023 366774
rect 500924 366720 500959 366740
rect 500993 366720 501023 366754
rect 500924 366684 501023 366720
rect 500924 366650 500944 366684
rect 500978 366664 501023 366684
rect 500924 366630 500959 366650
rect 500993 366630 501023 366664
rect 501087 367602 502049 367621
rect 501087 367600 501163 367602
rect 501087 367566 501104 367600
rect 501138 367568 501163 367600
rect 501197 367568 501253 367602
rect 501287 367568 501343 367602
rect 501377 367568 501433 367602
rect 501467 367568 501523 367602
rect 501557 367568 501613 367602
rect 501647 367568 501703 367602
rect 501737 367568 501793 367602
rect 501827 367568 501883 367602
rect 501917 367568 502049 367602
rect 501138 367566 502049 367568
rect 501087 367549 502049 367566
rect 501087 367510 501159 367549
rect 501087 367476 501104 367510
rect 501138 367490 501159 367510
rect 501087 367456 501106 367476
rect 501140 367456 501159 367490
rect 501977 367524 502049 367549
rect 501977 367490 501996 367524
rect 502030 367490 502049 367524
rect 501087 367420 501159 367456
rect 501087 367386 501104 367420
rect 501138 367400 501159 367420
rect 501087 367366 501106 367386
rect 501140 367366 501159 367400
rect 501087 367330 501159 367366
rect 501087 367296 501104 367330
rect 501138 367310 501159 367330
rect 501087 367276 501106 367296
rect 501140 367276 501159 367310
rect 501087 367240 501159 367276
rect 501087 367206 501104 367240
rect 501138 367220 501159 367240
rect 501087 367186 501106 367206
rect 501140 367186 501159 367220
rect 501087 367150 501159 367186
rect 501087 367116 501104 367150
rect 501138 367130 501159 367150
rect 501087 367096 501106 367116
rect 501140 367096 501159 367130
rect 501087 367060 501159 367096
rect 501087 367026 501104 367060
rect 501138 367040 501159 367060
rect 501087 367006 501106 367026
rect 501140 367006 501159 367040
rect 501087 366970 501159 367006
rect 501087 366936 501104 366970
rect 501138 366950 501159 366970
rect 501087 366916 501106 366936
rect 501140 366916 501159 366950
rect 501087 366880 501159 366916
rect 501087 366846 501104 366880
rect 501138 366860 501159 366880
rect 501087 366826 501106 366846
rect 501140 366826 501159 366860
rect 501087 366790 501159 366826
rect 501221 367426 501915 367487
rect 501221 367392 501280 367426
rect 501314 367414 501370 367426
rect 501342 367392 501370 367414
rect 501404 367414 501460 367426
rect 501404 367392 501408 367414
rect 501221 367380 501308 367392
rect 501342 367380 501408 367392
rect 501442 367392 501460 367414
rect 501494 367414 501550 367426
rect 501494 367392 501508 367414
rect 501442 367380 501508 367392
rect 501542 367392 501550 367414
rect 501584 367414 501640 367426
rect 501674 367414 501730 367426
rect 501764 367414 501820 367426
rect 501584 367392 501608 367414
rect 501674 367392 501708 367414
rect 501764 367392 501808 367414
rect 501854 367392 501915 367426
rect 501542 367380 501608 367392
rect 501642 367380 501708 367392
rect 501742 367380 501808 367392
rect 501842 367380 501915 367392
rect 501221 367336 501915 367380
rect 501221 367302 501280 367336
rect 501314 367314 501370 367336
rect 501342 367302 501370 367314
rect 501404 367314 501460 367336
rect 501404 367302 501408 367314
rect 501221 367280 501308 367302
rect 501342 367280 501408 367302
rect 501442 367302 501460 367314
rect 501494 367314 501550 367336
rect 501494 367302 501508 367314
rect 501442 367280 501508 367302
rect 501542 367302 501550 367314
rect 501584 367314 501640 367336
rect 501674 367314 501730 367336
rect 501764 367314 501820 367336
rect 501584 367302 501608 367314
rect 501674 367302 501708 367314
rect 501764 367302 501808 367314
rect 501854 367302 501915 367336
rect 501542 367280 501608 367302
rect 501642 367280 501708 367302
rect 501742 367280 501808 367302
rect 501842 367280 501915 367302
rect 501221 367246 501915 367280
rect 501221 367212 501280 367246
rect 501314 367214 501370 367246
rect 501342 367212 501370 367214
rect 501404 367214 501460 367246
rect 501404 367212 501408 367214
rect 501221 367180 501308 367212
rect 501342 367180 501408 367212
rect 501442 367212 501460 367214
rect 501494 367214 501550 367246
rect 501494 367212 501508 367214
rect 501442 367180 501508 367212
rect 501542 367212 501550 367214
rect 501584 367214 501640 367246
rect 501674 367214 501730 367246
rect 501764 367214 501820 367246
rect 501584 367212 501608 367214
rect 501674 367212 501708 367214
rect 501764 367212 501808 367214
rect 501854 367212 501915 367246
rect 501542 367180 501608 367212
rect 501642 367180 501708 367212
rect 501742 367180 501808 367212
rect 501842 367180 501915 367212
rect 501221 367156 501915 367180
rect 501221 367122 501280 367156
rect 501314 367122 501370 367156
rect 501404 367122 501460 367156
rect 501494 367122 501550 367156
rect 501584 367122 501640 367156
rect 501674 367122 501730 367156
rect 501764 367122 501820 367156
rect 501854 367122 501915 367156
rect 501221 367114 501915 367122
rect 501221 367080 501308 367114
rect 501342 367080 501408 367114
rect 501442 367080 501508 367114
rect 501542 367080 501608 367114
rect 501642 367080 501708 367114
rect 501742 367080 501808 367114
rect 501842 367080 501915 367114
rect 501221 367066 501915 367080
rect 501221 367032 501280 367066
rect 501314 367032 501370 367066
rect 501404 367032 501460 367066
rect 501494 367032 501550 367066
rect 501584 367032 501640 367066
rect 501674 367032 501730 367066
rect 501764 367032 501820 367066
rect 501854 367032 501915 367066
rect 501221 367014 501915 367032
rect 501221 366980 501308 367014
rect 501342 366980 501408 367014
rect 501442 366980 501508 367014
rect 501542 366980 501608 367014
rect 501642 366980 501708 367014
rect 501742 366980 501808 367014
rect 501842 366980 501915 367014
rect 501221 366976 501915 366980
rect 501221 366942 501280 366976
rect 501314 366942 501370 366976
rect 501404 366942 501460 366976
rect 501494 366942 501550 366976
rect 501584 366942 501640 366976
rect 501674 366942 501730 366976
rect 501764 366942 501820 366976
rect 501854 366942 501915 366976
rect 501221 366914 501915 366942
rect 501221 366886 501308 366914
rect 501342 366886 501408 366914
rect 501221 366852 501280 366886
rect 501342 366880 501370 366886
rect 501314 366852 501370 366880
rect 501404 366880 501408 366886
rect 501442 366886 501508 366914
rect 501442 366880 501460 366886
rect 501404 366852 501460 366880
rect 501494 366880 501508 366886
rect 501542 366886 501608 366914
rect 501642 366886 501708 366914
rect 501742 366886 501808 366914
rect 501842 366886 501915 366914
rect 501542 366880 501550 366886
rect 501494 366852 501550 366880
rect 501584 366880 501608 366886
rect 501674 366880 501708 366886
rect 501764 366880 501808 366886
rect 501584 366852 501640 366880
rect 501674 366852 501730 366880
rect 501764 366852 501820 366880
rect 501854 366852 501915 366886
rect 501221 366793 501915 366852
rect 501977 367434 502049 367490
rect 501977 367400 501996 367434
rect 502030 367400 502049 367434
rect 501977 367344 502049 367400
rect 501977 367310 501996 367344
rect 502030 367310 502049 367344
rect 501977 367254 502049 367310
rect 501977 367220 501996 367254
rect 502030 367220 502049 367254
rect 501977 367164 502049 367220
rect 501977 367130 501996 367164
rect 502030 367130 502049 367164
rect 501977 367074 502049 367130
rect 501977 367040 501996 367074
rect 502030 367040 502049 367074
rect 501977 366984 502049 367040
rect 501977 366950 501996 366984
rect 502030 366950 502049 366984
rect 501977 366894 502049 366950
rect 501977 366860 501996 366894
rect 502030 366860 502049 366894
rect 501977 366804 502049 366860
rect 501087 366756 501104 366790
rect 501138 366770 501159 366790
rect 501087 366736 501106 366756
rect 501140 366736 501159 366770
rect 501087 366731 501159 366736
rect 501977 366770 501996 366804
rect 502030 366770 502049 366804
rect 501977 366731 502049 366770
rect 501087 366712 502049 366731
rect 501087 366700 501182 366712
rect 501087 366666 501104 366700
rect 501138 366678 501182 366700
rect 501216 366678 501272 366712
rect 501306 366678 501362 366712
rect 501396 366678 501452 366712
rect 501486 366678 501542 366712
rect 501576 366678 501632 366712
rect 501666 366678 501722 366712
rect 501756 366678 501812 366712
rect 501846 366678 501902 366712
rect 501936 366678 502049 366712
rect 501138 366666 502049 366678
rect 501087 366659 502049 366666
rect 502113 367620 502146 367654
rect 502180 367620 502212 367654
rect 502113 367564 502212 367620
rect 502113 367530 502146 367564
rect 502180 367530 502212 367564
rect 502113 367474 502212 367530
rect 502113 367440 502146 367474
rect 502180 367440 502212 367474
rect 502113 367384 502212 367440
rect 502113 367350 502146 367384
rect 502180 367350 502212 367384
rect 502113 367294 502212 367350
rect 502113 367260 502146 367294
rect 502180 367260 502212 367294
rect 502113 367204 502212 367260
rect 502113 367170 502146 367204
rect 502180 367170 502212 367204
rect 502113 367114 502212 367170
rect 502113 367080 502146 367114
rect 502180 367080 502212 367114
rect 502113 367024 502212 367080
rect 502113 366990 502146 367024
rect 502180 366990 502212 367024
rect 502113 366934 502212 366990
rect 502113 366900 502146 366934
rect 502180 366900 502212 366934
rect 502113 366844 502212 366900
rect 502113 366810 502146 366844
rect 502180 366810 502212 366844
rect 502113 366754 502212 366810
rect 502113 366720 502146 366754
rect 502180 366720 502212 366754
rect 502113 366664 502212 366720
rect 500924 366595 501023 366630
rect 502113 366630 502146 366664
rect 502180 366630 502212 366664
rect 502113 366595 502212 366630
rect 500924 366594 502212 366595
rect 500924 366560 500944 366594
rect 500978 366563 502212 366594
rect 500978 366560 500982 366563
rect 500924 366529 500982 366560
rect 501016 366529 501072 366563
rect 501106 366529 501162 366563
rect 501196 366529 501252 366563
rect 501286 366529 501342 366563
rect 501376 366529 501432 366563
rect 501466 366529 501522 366563
rect 501556 366529 501612 366563
rect 501646 366529 501702 366563
rect 501736 366529 501792 366563
rect 501826 366529 501882 366563
rect 501916 366529 501972 366563
rect 502006 366529 502062 366563
rect 502096 366529 502212 366563
rect 500924 366424 502212 366529
rect 500924 366390 500944 366424
rect 500978 366410 502212 366424
rect 500978 366390 500982 366410
rect 500924 366376 500982 366390
rect 501016 366376 501072 366410
rect 501106 366376 501162 366410
rect 501196 366376 501252 366410
rect 501286 366376 501342 366410
rect 501376 366376 501432 366410
rect 501466 366376 501522 366410
rect 501556 366376 501612 366410
rect 501646 366376 501702 366410
rect 501736 366376 501792 366410
rect 501826 366376 501882 366410
rect 501916 366376 501972 366410
rect 502006 366376 502062 366410
rect 502096 366376 502212 366410
rect 500924 366345 502212 366376
rect 500924 366334 501023 366345
rect 500924 366300 500944 366334
rect 500978 366314 501023 366334
rect 500924 366280 500959 366300
rect 500993 366280 501023 366314
rect 502113 366314 502212 366345
rect 500924 366244 501023 366280
rect 500924 366210 500944 366244
rect 500978 366224 501023 366244
rect 500924 366190 500959 366210
rect 500993 366190 501023 366224
rect 500924 366154 501023 366190
rect 500924 366120 500944 366154
rect 500978 366134 501023 366154
rect 500924 366100 500959 366120
rect 500993 366100 501023 366134
rect 500924 366064 501023 366100
rect 500924 366030 500944 366064
rect 500978 366044 501023 366064
rect 500924 366010 500959 366030
rect 500993 366010 501023 366044
rect 500924 365974 501023 366010
rect 500924 365940 500944 365974
rect 500978 365954 501023 365974
rect 500924 365920 500959 365940
rect 500993 365920 501023 365954
rect 500924 365884 501023 365920
rect 500924 365850 500944 365884
rect 500978 365864 501023 365884
rect 500924 365830 500959 365850
rect 500993 365830 501023 365864
rect 500924 365794 501023 365830
rect 500924 365760 500944 365794
rect 500978 365774 501023 365794
rect 500924 365740 500959 365760
rect 500993 365740 501023 365774
rect 500924 365704 501023 365740
rect 500924 365670 500944 365704
rect 500978 365684 501023 365704
rect 500924 365650 500959 365670
rect 500993 365650 501023 365684
rect 500924 365614 501023 365650
rect 500924 365580 500944 365614
rect 500978 365594 501023 365614
rect 500924 365560 500959 365580
rect 500993 365560 501023 365594
rect 500924 365524 501023 365560
rect 500924 365490 500944 365524
rect 500978 365504 501023 365524
rect 500924 365470 500959 365490
rect 500993 365470 501023 365504
rect 500924 365434 501023 365470
rect 500924 365400 500944 365434
rect 500978 365414 501023 365434
rect 500924 365380 500959 365400
rect 500993 365380 501023 365414
rect 500924 365344 501023 365380
rect 500924 365310 500944 365344
rect 500978 365324 501023 365344
rect 500924 365290 500959 365310
rect 500993 365290 501023 365324
rect 501087 366262 502049 366281
rect 501087 366260 501163 366262
rect 501087 366226 501104 366260
rect 501138 366228 501163 366260
rect 501197 366228 501253 366262
rect 501287 366228 501343 366262
rect 501377 366228 501433 366262
rect 501467 366228 501523 366262
rect 501557 366228 501613 366262
rect 501647 366228 501703 366262
rect 501737 366228 501793 366262
rect 501827 366228 501883 366262
rect 501917 366228 502049 366262
rect 501138 366226 502049 366228
rect 501087 366209 502049 366226
rect 501087 366170 501159 366209
rect 501087 366136 501104 366170
rect 501138 366150 501159 366170
rect 501087 366116 501106 366136
rect 501140 366116 501159 366150
rect 501977 366184 502049 366209
rect 501977 366150 501996 366184
rect 502030 366150 502049 366184
rect 501087 366080 501159 366116
rect 501087 366046 501104 366080
rect 501138 366060 501159 366080
rect 501087 366026 501106 366046
rect 501140 366026 501159 366060
rect 501087 365990 501159 366026
rect 501087 365956 501104 365990
rect 501138 365970 501159 365990
rect 501087 365936 501106 365956
rect 501140 365936 501159 365970
rect 501087 365900 501159 365936
rect 501087 365866 501104 365900
rect 501138 365880 501159 365900
rect 501087 365846 501106 365866
rect 501140 365846 501159 365880
rect 501087 365810 501159 365846
rect 501087 365776 501104 365810
rect 501138 365790 501159 365810
rect 501087 365756 501106 365776
rect 501140 365756 501159 365790
rect 501087 365720 501159 365756
rect 501087 365686 501104 365720
rect 501138 365700 501159 365720
rect 501087 365666 501106 365686
rect 501140 365666 501159 365700
rect 501087 365630 501159 365666
rect 501087 365596 501104 365630
rect 501138 365610 501159 365630
rect 501087 365576 501106 365596
rect 501140 365576 501159 365610
rect 501087 365540 501159 365576
rect 501087 365506 501104 365540
rect 501138 365520 501159 365540
rect 501087 365486 501106 365506
rect 501140 365486 501159 365520
rect 501087 365450 501159 365486
rect 501221 366086 501915 366147
rect 501221 366052 501280 366086
rect 501314 366074 501370 366086
rect 501342 366052 501370 366074
rect 501404 366074 501460 366086
rect 501404 366052 501408 366074
rect 501221 366040 501308 366052
rect 501342 366040 501408 366052
rect 501442 366052 501460 366074
rect 501494 366074 501550 366086
rect 501494 366052 501508 366074
rect 501442 366040 501508 366052
rect 501542 366052 501550 366074
rect 501584 366074 501640 366086
rect 501674 366074 501730 366086
rect 501764 366074 501820 366086
rect 501584 366052 501608 366074
rect 501674 366052 501708 366074
rect 501764 366052 501808 366074
rect 501854 366052 501915 366086
rect 501542 366040 501608 366052
rect 501642 366040 501708 366052
rect 501742 366040 501808 366052
rect 501842 366040 501915 366052
rect 501221 365996 501915 366040
rect 501221 365962 501280 365996
rect 501314 365974 501370 365996
rect 501342 365962 501370 365974
rect 501404 365974 501460 365996
rect 501404 365962 501408 365974
rect 501221 365940 501308 365962
rect 501342 365940 501408 365962
rect 501442 365962 501460 365974
rect 501494 365974 501550 365996
rect 501494 365962 501508 365974
rect 501442 365940 501508 365962
rect 501542 365962 501550 365974
rect 501584 365974 501640 365996
rect 501674 365974 501730 365996
rect 501764 365974 501820 365996
rect 501584 365962 501608 365974
rect 501674 365962 501708 365974
rect 501764 365962 501808 365974
rect 501854 365962 501915 365996
rect 501542 365940 501608 365962
rect 501642 365940 501708 365962
rect 501742 365940 501808 365962
rect 501842 365940 501915 365962
rect 501221 365906 501915 365940
rect 501221 365872 501280 365906
rect 501314 365874 501370 365906
rect 501342 365872 501370 365874
rect 501404 365874 501460 365906
rect 501404 365872 501408 365874
rect 501221 365840 501308 365872
rect 501342 365840 501408 365872
rect 501442 365872 501460 365874
rect 501494 365874 501550 365906
rect 501494 365872 501508 365874
rect 501442 365840 501508 365872
rect 501542 365872 501550 365874
rect 501584 365874 501640 365906
rect 501674 365874 501730 365906
rect 501764 365874 501820 365906
rect 501584 365872 501608 365874
rect 501674 365872 501708 365874
rect 501764 365872 501808 365874
rect 501854 365872 501915 365906
rect 501542 365840 501608 365872
rect 501642 365840 501708 365872
rect 501742 365840 501808 365872
rect 501842 365840 501915 365872
rect 501221 365816 501915 365840
rect 501221 365782 501280 365816
rect 501314 365782 501370 365816
rect 501404 365782 501460 365816
rect 501494 365782 501550 365816
rect 501584 365782 501640 365816
rect 501674 365782 501730 365816
rect 501764 365782 501820 365816
rect 501854 365782 501915 365816
rect 501221 365774 501915 365782
rect 501221 365740 501308 365774
rect 501342 365740 501408 365774
rect 501442 365740 501508 365774
rect 501542 365740 501608 365774
rect 501642 365740 501708 365774
rect 501742 365740 501808 365774
rect 501842 365740 501915 365774
rect 501221 365726 501915 365740
rect 501221 365692 501280 365726
rect 501314 365692 501370 365726
rect 501404 365692 501460 365726
rect 501494 365692 501550 365726
rect 501584 365692 501640 365726
rect 501674 365692 501730 365726
rect 501764 365692 501820 365726
rect 501854 365692 501915 365726
rect 501221 365674 501915 365692
rect 501221 365640 501308 365674
rect 501342 365640 501408 365674
rect 501442 365640 501508 365674
rect 501542 365640 501608 365674
rect 501642 365640 501708 365674
rect 501742 365640 501808 365674
rect 501842 365640 501915 365674
rect 501221 365636 501915 365640
rect 501221 365602 501280 365636
rect 501314 365602 501370 365636
rect 501404 365602 501460 365636
rect 501494 365602 501550 365636
rect 501584 365602 501640 365636
rect 501674 365602 501730 365636
rect 501764 365602 501820 365636
rect 501854 365602 501915 365636
rect 501221 365574 501915 365602
rect 501221 365546 501308 365574
rect 501342 365546 501408 365574
rect 501221 365512 501280 365546
rect 501342 365540 501370 365546
rect 501314 365512 501370 365540
rect 501404 365540 501408 365546
rect 501442 365546 501508 365574
rect 501442 365540 501460 365546
rect 501404 365512 501460 365540
rect 501494 365540 501508 365546
rect 501542 365546 501608 365574
rect 501642 365546 501708 365574
rect 501742 365546 501808 365574
rect 501842 365546 501915 365574
rect 501542 365540 501550 365546
rect 501494 365512 501550 365540
rect 501584 365540 501608 365546
rect 501674 365540 501708 365546
rect 501764 365540 501808 365546
rect 501584 365512 501640 365540
rect 501674 365512 501730 365540
rect 501764 365512 501820 365540
rect 501854 365512 501915 365546
rect 501221 365453 501915 365512
rect 501977 366094 502049 366150
rect 501977 366060 501996 366094
rect 502030 366060 502049 366094
rect 501977 366004 502049 366060
rect 501977 365970 501996 366004
rect 502030 365970 502049 366004
rect 501977 365914 502049 365970
rect 501977 365880 501996 365914
rect 502030 365880 502049 365914
rect 501977 365824 502049 365880
rect 501977 365790 501996 365824
rect 502030 365790 502049 365824
rect 501977 365734 502049 365790
rect 501977 365700 501996 365734
rect 502030 365700 502049 365734
rect 501977 365644 502049 365700
rect 501977 365610 501996 365644
rect 502030 365610 502049 365644
rect 501977 365554 502049 365610
rect 501977 365520 501996 365554
rect 502030 365520 502049 365554
rect 501977 365464 502049 365520
rect 501087 365416 501104 365450
rect 501138 365430 501159 365450
rect 501087 365396 501106 365416
rect 501140 365396 501159 365430
rect 501087 365391 501159 365396
rect 501977 365430 501996 365464
rect 502030 365430 502049 365464
rect 501977 365391 502049 365430
rect 501087 365372 502049 365391
rect 501087 365360 501182 365372
rect 501087 365326 501104 365360
rect 501138 365338 501182 365360
rect 501216 365338 501272 365372
rect 501306 365338 501362 365372
rect 501396 365338 501452 365372
rect 501486 365338 501542 365372
rect 501576 365338 501632 365372
rect 501666 365338 501722 365372
rect 501756 365338 501812 365372
rect 501846 365338 501902 365372
rect 501936 365338 502049 365372
rect 501138 365326 502049 365338
rect 501087 365319 502049 365326
rect 502113 366280 502146 366314
rect 502180 366280 502212 366314
rect 502113 366224 502212 366280
rect 502113 366190 502146 366224
rect 502180 366190 502212 366224
rect 502113 366134 502212 366190
rect 502113 366100 502146 366134
rect 502180 366100 502212 366134
rect 502113 366044 502212 366100
rect 502113 366010 502146 366044
rect 502180 366010 502212 366044
rect 502113 365954 502212 366010
rect 502113 365920 502146 365954
rect 502180 365920 502212 365954
rect 502113 365864 502212 365920
rect 502113 365830 502146 365864
rect 502180 365830 502212 365864
rect 502113 365774 502212 365830
rect 502113 365740 502146 365774
rect 502180 365740 502212 365774
rect 502113 365684 502212 365740
rect 502113 365650 502146 365684
rect 502180 365650 502212 365684
rect 502113 365594 502212 365650
rect 502113 365560 502146 365594
rect 502180 365560 502212 365594
rect 502113 365504 502212 365560
rect 502113 365470 502146 365504
rect 502180 365470 502212 365504
rect 502113 365414 502212 365470
rect 502113 365380 502146 365414
rect 502180 365380 502212 365414
rect 502113 365324 502212 365380
rect 500924 365255 501023 365290
rect 502113 365290 502146 365324
rect 502180 365290 502212 365324
rect 502113 365255 502212 365290
rect 500924 365254 502212 365255
rect 500924 365220 500944 365254
rect 500978 365223 502212 365254
rect 500978 365220 500982 365223
rect 500924 365189 500982 365220
rect 501016 365189 501072 365223
rect 501106 365189 501162 365223
rect 501196 365189 501252 365223
rect 501286 365189 501342 365223
rect 501376 365189 501432 365223
rect 501466 365189 501522 365223
rect 501556 365189 501612 365223
rect 501646 365189 501702 365223
rect 501736 365189 501792 365223
rect 501826 365189 501882 365223
rect 501916 365189 501972 365223
rect 502006 365189 502062 365223
rect 502096 365189 502212 365223
rect 500924 365084 502212 365189
rect 500924 365050 500944 365084
rect 500978 365070 502212 365084
rect 500978 365050 500982 365070
rect 500924 365036 500982 365050
rect 501016 365036 501072 365070
rect 501106 365036 501162 365070
rect 501196 365036 501252 365070
rect 501286 365036 501342 365070
rect 501376 365036 501432 365070
rect 501466 365036 501522 365070
rect 501556 365036 501612 365070
rect 501646 365036 501702 365070
rect 501736 365036 501792 365070
rect 501826 365036 501882 365070
rect 501916 365036 501972 365070
rect 502006 365036 502062 365070
rect 502096 365036 502212 365070
rect 500924 365005 502212 365036
rect 500924 364994 501023 365005
rect 500924 364960 500944 364994
rect 500978 364974 501023 364994
rect 500924 364940 500959 364960
rect 500993 364940 501023 364974
rect 502113 364974 502212 365005
rect 500924 364904 501023 364940
rect 500924 364870 500944 364904
rect 500978 364884 501023 364904
rect 500924 364850 500959 364870
rect 500993 364850 501023 364884
rect 500924 364814 501023 364850
rect 500924 364780 500944 364814
rect 500978 364794 501023 364814
rect 500924 364760 500959 364780
rect 500993 364760 501023 364794
rect 500924 364724 501023 364760
rect 500924 364690 500944 364724
rect 500978 364704 501023 364724
rect 500924 364670 500959 364690
rect 500993 364670 501023 364704
rect 500924 364634 501023 364670
rect 500924 364600 500944 364634
rect 500978 364614 501023 364634
rect 500924 364580 500959 364600
rect 500993 364580 501023 364614
rect 500924 364544 501023 364580
rect 500924 364510 500944 364544
rect 500978 364524 501023 364544
rect 500924 364490 500959 364510
rect 500993 364490 501023 364524
rect 500924 364454 501023 364490
rect 500924 364420 500944 364454
rect 500978 364434 501023 364454
rect 500924 364400 500959 364420
rect 500993 364400 501023 364434
rect 500924 364364 501023 364400
rect 500924 364330 500944 364364
rect 500978 364344 501023 364364
rect 500924 364310 500959 364330
rect 500993 364310 501023 364344
rect 500924 364274 501023 364310
rect 500924 364240 500944 364274
rect 500978 364254 501023 364274
rect 500924 364220 500959 364240
rect 500993 364220 501023 364254
rect 500924 364184 501023 364220
rect 500924 364150 500944 364184
rect 500978 364164 501023 364184
rect 500924 364130 500959 364150
rect 500993 364130 501023 364164
rect 500924 364094 501023 364130
rect 500924 364060 500944 364094
rect 500978 364074 501023 364094
rect 500924 364040 500959 364060
rect 500993 364040 501023 364074
rect 500924 364004 501023 364040
rect 500924 363970 500944 364004
rect 500978 363984 501023 364004
rect 500924 363950 500959 363970
rect 500993 363950 501023 363984
rect 501087 364922 502049 364941
rect 501087 364920 501163 364922
rect 501087 364886 501104 364920
rect 501138 364888 501163 364920
rect 501197 364888 501253 364922
rect 501287 364888 501343 364922
rect 501377 364888 501433 364922
rect 501467 364888 501523 364922
rect 501557 364888 501613 364922
rect 501647 364888 501703 364922
rect 501737 364888 501793 364922
rect 501827 364888 501883 364922
rect 501917 364888 502049 364922
rect 501138 364886 502049 364888
rect 501087 364869 502049 364886
rect 501087 364830 501159 364869
rect 501087 364796 501104 364830
rect 501138 364810 501159 364830
rect 501087 364776 501106 364796
rect 501140 364776 501159 364810
rect 501977 364844 502049 364869
rect 501977 364810 501996 364844
rect 502030 364810 502049 364844
rect 501087 364740 501159 364776
rect 501087 364706 501104 364740
rect 501138 364720 501159 364740
rect 501087 364686 501106 364706
rect 501140 364686 501159 364720
rect 501087 364650 501159 364686
rect 501087 364616 501104 364650
rect 501138 364630 501159 364650
rect 501087 364596 501106 364616
rect 501140 364596 501159 364630
rect 501087 364560 501159 364596
rect 501087 364526 501104 364560
rect 501138 364540 501159 364560
rect 501087 364506 501106 364526
rect 501140 364506 501159 364540
rect 501087 364470 501159 364506
rect 501087 364436 501104 364470
rect 501138 364450 501159 364470
rect 501087 364416 501106 364436
rect 501140 364416 501159 364450
rect 501087 364380 501159 364416
rect 501087 364346 501104 364380
rect 501138 364360 501159 364380
rect 501087 364326 501106 364346
rect 501140 364326 501159 364360
rect 501087 364290 501159 364326
rect 501087 364256 501104 364290
rect 501138 364270 501159 364290
rect 501087 364236 501106 364256
rect 501140 364236 501159 364270
rect 501087 364200 501159 364236
rect 501087 364166 501104 364200
rect 501138 364180 501159 364200
rect 501087 364146 501106 364166
rect 501140 364146 501159 364180
rect 501087 364110 501159 364146
rect 501221 364746 501915 364807
rect 501221 364712 501280 364746
rect 501314 364734 501370 364746
rect 501342 364712 501370 364734
rect 501404 364734 501460 364746
rect 501404 364712 501408 364734
rect 501221 364700 501308 364712
rect 501342 364700 501408 364712
rect 501442 364712 501460 364734
rect 501494 364734 501550 364746
rect 501494 364712 501508 364734
rect 501442 364700 501508 364712
rect 501542 364712 501550 364734
rect 501584 364734 501640 364746
rect 501674 364734 501730 364746
rect 501764 364734 501820 364746
rect 501584 364712 501608 364734
rect 501674 364712 501708 364734
rect 501764 364712 501808 364734
rect 501854 364712 501915 364746
rect 501542 364700 501608 364712
rect 501642 364700 501708 364712
rect 501742 364700 501808 364712
rect 501842 364700 501915 364712
rect 501221 364656 501915 364700
rect 501221 364622 501280 364656
rect 501314 364634 501370 364656
rect 501342 364622 501370 364634
rect 501404 364634 501460 364656
rect 501404 364622 501408 364634
rect 501221 364600 501308 364622
rect 501342 364600 501408 364622
rect 501442 364622 501460 364634
rect 501494 364634 501550 364656
rect 501494 364622 501508 364634
rect 501442 364600 501508 364622
rect 501542 364622 501550 364634
rect 501584 364634 501640 364656
rect 501674 364634 501730 364656
rect 501764 364634 501820 364656
rect 501584 364622 501608 364634
rect 501674 364622 501708 364634
rect 501764 364622 501808 364634
rect 501854 364622 501915 364656
rect 501542 364600 501608 364622
rect 501642 364600 501708 364622
rect 501742 364600 501808 364622
rect 501842 364600 501915 364622
rect 501221 364566 501915 364600
rect 501221 364532 501280 364566
rect 501314 364534 501370 364566
rect 501342 364532 501370 364534
rect 501404 364534 501460 364566
rect 501404 364532 501408 364534
rect 501221 364500 501308 364532
rect 501342 364500 501408 364532
rect 501442 364532 501460 364534
rect 501494 364534 501550 364566
rect 501494 364532 501508 364534
rect 501442 364500 501508 364532
rect 501542 364532 501550 364534
rect 501584 364534 501640 364566
rect 501674 364534 501730 364566
rect 501764 364534 501820 364566
rect 501584 364532 501608 364534
rect 501674 364532 501708 364534
rect 501764 364532 501808 364534
rect 501854 364532 501915 364566
rect 501542 364500 501608 364532
rect 501642 364500 501708 364532
rect 501742 364500 501808 364532
rect 501842 364500 501915 364532
rect 501221 364476 501915 364500
rect 501221 364442 501280 364476
rect 501314 364442 501370 364476
rect 501404 364442 501460 364476
rect 501494 364442 501550 364476
rect 501584 364442 501640 364476
rect 501674 364442 501730 364476
rect 501764 364442 501820 364476
rect 501854 364442 501915 364476
rect 501221 364434 501915 364442
rect 501221 364400 501308 364434
rect 501342 364400 501408 364434
rect 501442 364400 501508 364434
rect 501542 364400 501608 364434
rect 501642 364400 501708 364434
rect 501742 364400 501808 364434
rect 501842 364400 501915 364434
rect 501221 364386 501915 364400
rect 501221 364352 501280 364386
rect 501314 364352 501370 364386
rect 501404 364352 501460 364386
rect 501494 364352 501550 364386
rect 501584 364352 501640 364386
rect 501674 364352 501730 364386
rect 501764 364352 501820 364386
rect 501854 364352 501915 364386
rect 501221 364334 501915 364352
rect 501221 364300 501308 364334
rect 501342 364300 501408 364334
rect 501442 364300 501508 364334
rect 501542 364300 501608 364334
rect 501642 364300 501708 364334
rect 501742 364300 501808 364334
rect 501842 364300 501915 364334
rect 501221 364296 501915 364300
rect 501221 364262 501280 364296
rect 501314 364262 501370 364296
rect 501404 364262 501460 364296
rect 501494 364262 501550 364296
rect 501584 364262 501640 364296
rect 501674 364262 501730 364296
rect 501764 364262 501820 364296
rect 501854 364262 501915 364296
rect 501221 364234 501915 364262
rect 501221 364206 501308 364234
rect 501342 364206 501408 364234
rect 501221 364172 501280 364206
rect 501342 364200 501370 364206
rect 501314 364172 501370 364200
rect 501404 364200 501408 364206
rect 501442 364206 501508 364234
rect 501442 364200 501460 364206
rect 501404 364172 501460 364200
rect 501494 364200 501508 364206
rect 501542 364206 501608 364234
rect 501642 364206 501708 364234
rect 501742 364206 501808 364234
rect 501842 364206 501915 364234
rect 501542 364200 501550 364206
rect 501494 364172 501550 364200
rect 501584 364200 501608 364206
rect 501674 364200 501708 364206
rect 501764 364200 501808 364206
rect 501584 364172 501640 364200
rect 501674 364172 501730 364200
rect 501764 364172 501820 364200
rect 501854 364172 501915 364206
rect 501221 364113 501915 364172
rect 501977 364754 502049 364810
rect 501977 364720 501996 364754
rect 502030 364720 502049 364754
rect 501977 364664 502049 364720
rect 501977 364630 501996 364664
rect 502030 364630 502049 364664
rect 501977 364574 502049 364630
rect 501977 364540 501996 364574
rect 502030 364540 502049 364574
rect 501977 364484 502049 364540
rect 501977 364450 501996 364484
rect 502030 364450 502049 364484
rect 501977 364394 502049 364450
rect 501977 364360 501996 364394
rect 502030 364360 502049 364394
rect 501977 364304 502049 364360
rect 501977 364270 501996 364304
rect 502030 364270 502049 364304
rect 501977 364214 502049 364270
rect 501977 364180 501996 364214
rect 502030 364180 502049 364214
rect 501977 364124 502049 364180
rect 501087 364076 501104 364110
rect 501138 364090 501159 364110
rect 501087 364056 501106 364076
rect 501140 364056 501159 364090
rect 501087 364051 501159 364056
rect 501977 364090 501996 364124
rect 502030 364090 502049 364124
rect 501977 364051 502049 364090
rect 501087 364032 502049 364051
rect 501087 364020 501182 364032
rect 501087 363986 501104 364020
rect 501138 363998 501182 364020
rect 501216 363998 501272 364032
rect 501306 363998 501362 364032
rect 501396 363998 501452 364032
rect 501486 363998 501542 364032
rect 501576 363998 501632 364032
rect 501666 363998 501722 364032
rect 501756 363998 501812 364032
rect 501846 363998 501902 364032
rect 501936 363998 502049 364032
rect 501138 363986 502049 363998
rect 501087 363979 502049 363986
rect 502113 364940 502146 364974
rect 502180 364940 502212 364974
rect 502113 364884 502212 364940
rect 502113 364850 502146 364884
rect 502180 364850 502212 364884
rect 502113 364794 502212 364850
rect 502113 364760 502146 364794
rect 502180 364760 502212 364794
rect 502113 364704 502212 364760
rect 502113 364670 502146 364704
rect 502180 364670 502212 364704
rect 502113 364614 502212 364670
rect 502113 364580 502146 364614
rect 502180 364580 502212 364614
rect 502113 364524 502212 364580
rect 502113 364490 502146 364524
rect 502180 364490 502212 364524
rect 502113 364434 502212 364490
rect 502113 364400 502146 364434
rect 502180 364400 502212 364434
rect 502113 364344 502212 364400
rect 502113 364310 502146 364344
rect 502180 364310 502212 364344
rect 502113 364254 502212 364310
rect 502113 364220 502146 364254
rect 502180 364220 502212 364254
rect 502113 364164 502212 364220
rect 502113 364130 502146 364164
rect 502180 364130 502212 364164
rect 502113 364074 502212 364130
rect 502113 364040 502146 364074
rect 502180 364040 502212 364074
rect 502113 363984 502212 364040
rect 500924 363915 501023 363950
rect 502113 363950 502146 363984
rect 502180 363950 502212 363984
rect 502113 363915 502212 363950
rect 500924 363914 502212 363915
rect 500924 363880 500944 363914
rect 500978 363883 502212 363914
rect 500978 363880 500982 363883
rect 500924 363849 500982 363880
rect 501016 363849 501072 363883
rect 501106 363849 501162 363883
rect 501196 363849 501252 363883
rect 501286 363849 501342 363883
rect 501376 363849 501432 363883
rect 501466 363849 501522 363883
rect 501556 363849 501612 363883
rect 501646 363849 501702 363883
rect 501736 363849 501792 363883
rect 501826 363849 501882 363883
rect 501916 363849 501972 363883
rect 502006 363849 502062 363883
rect 502096 363849 502212 363883
rect 500924 363744 502212 363849
rect 500924 363710 500944 363744
rect 500978 363730 502212 363744
rect 500978 363710 500982 363730
rect 500924 363696 500982 363710
rect 501016 363696 501072 363730
rect 501106 363696 501162 363730
rect 501196 363696 501252 363730
rect 501286 363696 501342 363730
rect 501376 363696 501432 363730
rect 501466 363696 501522 363730
rect 501556 363696 501612 363730
rect 501646 363696 501702 363730
rect 501736 363696 501792 363730
rect 501826 363696 501882 363730
rect 501916 363696 501972 363730
rect 502006 363696 502062 363730
rect 502096 363696 502212 363730
rect 500924 363665 502212 363696
rect 500924 363654 501023 363665
rect 500924 363620 500944 363654
rect 500978 363634 501023 363654
rect 500924 363600 500959 363620
rect 500993 363600 501023 363634
rect 502113 363634 502212 363665
rect 500924 363564 501023 363600
rect 500924 363530 500944 363564
rect 500978 363544 501023 363564
rect 500924 363510 500959 363530
rect 500993 363510 501023 363544
rect 500924 363474 501023 363510
rect 500924 363440 500944 363474
rect 500978 363454 501023 363474
rect 500924 363420 500959 363440
rect 500993 363420 501023 363454
rect 500924 363384 501023 363420
rect 500924 363350 500944 363384
rect 500978 363364 501023 363384
rect 500924 363330 500959 363350
rect 500993 363330 501023 363364
rect 500924 363294 501023 363330
rect 500924 363260 500944 363294
rect 500978 363274 501023 363294
rect 500924 363240 500959 363260
rect 500993 363240 501023 363274
rect 500924 363204 501023 363240
rect 500924 363170 500944 363204
rect 500978 363184 501023 363204
rect 500924 363150 500959 363170
rect 500993 363150 501023 363184
rect 500924 363114 501023 363150
rect 500924 363080 500944 363114
rect 500978 363094 501023 363114
rect 500924 363060 500959 363080
rect 500993 363060 501023 363094
rect 500924 363024 501023 363060
rect 500924 362990 500944 363024
rect 500978 363004 501023 363024
rect 500924 362970 500959 362990
rect 500993 362970 501023 363004
rect 500924 362934 501023 362970
rect 500924 362900 500944 362934
rect 500978 362914 501023 362934
rect 500924 362880 500959 362900
rect 500993 362880 501023 362914
rect 500924 362844 501023 362880
rect 500924 362810 500944 362844
rect 500978 362824 501023 362844
rect 500924 362790 500959 362810
rect 500993 362790 501023 362824
rect 500924 362754 501023 362790
rect 500924 362720 500944 362754
rect 500978 362734 501023 362754
rect 500924 362700 500959 362720
rect 500993 362700 501023 362734
rect 500924 362664 501023 362700
rect 500924 362630 500944 362664
rect 500978 362644 501023 362664
rect 500924 362610 500959 362630
rect 500993 362610 501023 362644
rect 501087 363582 502049 363601
rect 501087 363580 501163 363582
rect 501087 363546 501104 363580
rect 501138 363548 501163 363580
rect 501197 363548 501253 363582
rect 501287 363548 501343 363582
rect 501377 363548 501433 363582
rect 501467 363548 501523 363582
rect 501557 363548 501613 363582
rect 501647 363548 501703 363582
rect 501737 363548 501793 363582
rect 501827 363548 501883 363582
rect 501917 363548 502049 363582
rect 501138 363546 502049 363548
rect 501087 363529 502049 363546
rect 501087 363490 501159 363529
rect 501087 363456 501104 363490
rect 501138 363470 501159 363490
rect 501087 363436 501106 363456
rect 501140 363436 501159 363470
rect 501977 363504 502049 363529
rect 501977 363470 501996 363504
rect 502030 363470 502049 363504
rect 501087 363400 501159 363436
rect 501087 363366 501104 363400
rect 501138 363380 501159 363400
rect 501087 363346 501106 363366
rect 501140 363346 501159 363380
rect 501087 363310 501159 363346
rect 501087 363276 501104 363310
rect 501138 363290 501159 363310
rect 501087 363256 501106 363276
rect 501140 363256 501159 363290
rect 501087 363220 501159 363256
rect 501087 363186 501104 363220
rect 501138 363200 501159 363220
rect 501087 363166 501106 363186
rect 501140 363166 501159 363200
rect 501087 363130 501159 363166
rect 501087 363096 501104 363130
rect 501138 363110 501159 363130
rect 501087 363076 501106 363096
rect 501140 363076 501159 363110
rect 501087 363040 501159 363076
rect 501087 363006 501104 363040
rect 501138 363020 501159 363040
rect 501087 362986 501106 363006
rect 501140 362986 501159 363020
rect 501087 362950 501159 362986
rect 501087 362916 501104 362950
rect 501138 362930 501159 362950
rect 501087 362896 501106 362916
rect 501140 362896 501159 362930
rect 501087 362860 501159 362896
rect 501087 362826 501104 362860
rect 501138 362840 501159 362860
rect 501087 362806 501106 362826
rect 501140 362806 501159 362840
rect 501087 362770 501159 362806
rect 501221 363406 501915 363467
rect 501221 363372 501280 363406
rect 501314 363394 501370 363406
rect 501342 363372 501370 363394
rect 501404 363394 501460 363406
rect 501404 363372 501408 363394
rect 501221 363360 501308 363372
rect 501342 363360 501408 363372
rect 501442 363372 501460 363394
rect 501494 363394 501550 363406
rect 501494 363372 501508 363394
rect 501442 363360 501508 363372
rect 501542 363372 501550 363394
rect 501584 363394 501640 363406
rect 501674 363394 501730 363406
rect 501764 363394 501820 363406
rect 501584 363372 501608 363394
rect 501674 363372 501708 363394
rect 501764 363372 501808 363394
rect 501854 363372 501915 363406
rect 501542 363360 501608 363372
rect 501642 363360 501708 363372
rect 501742 363360 501808 363372
rect 501842 363360 501915 363372
rect 501221 363316 501915 363360
rect 501221 363282 501280 363316
rect 501314 363294 501370 363316
rect 501342 363282 501370 363294
rect 501404 363294 501460 363316
rect 501404 363282 501408 363294
rect 501221 363260 501308 363282
rect 501342 363260 501408 363282
rect 501442 363282 501460 363294
rect 501494 363294 501550 363316
rect 501494 363282 501508 363294
rect 501442 363260 501508 363282
rect 501542 363282 501550 363294
rect 501584 363294 501640 363316
rect 501674 363294 501730 363316
rect 501764 363294 501820 363316
rect 501584 363282 501608 363294
rect 501674 363282 501708 363294
rect 501764 363282 501808 363294
rect 501854 363282 501915 363316
rect 501542 363260 501608 363282
rect 501642 363260 501708 363282
rect 501742 363260 501808 363282
rect 501842 363260 501915 363282
rect 501221 363226 501915 363260
rect 501221 363192 501280 363226
rect 501314 363194 501370 363226
rect 501342 363192 501370 363194
rect 501404 363194 501460 363226
rect 501404 363192 501408 363194
rect 501221 363160 501308 363192
rect 501342 363160 501408 363192
rect 501442 363192 501460 363194
rect 501494 363194 501550 363226
rect 501494 363192 501508 363194
rect 501442 363160 501508 363192
rect 501542 363192 501550 363194
rect 501584 363194 501640 363226
rect 501674 363194 501730 363226
rect 501764 363194 501820 363226
rect 501584 363192 501608 363194
rect 501674 363192 501708 363194
rect 501764 363192 501808 363194
rect 501854 363192 501915 363226
rect 501542 363160 501608 363192
rect 501642 363160 501708 363192
rect 501742 363160 501808 363192
rect 501842 363160 501915 363192
rect 501221 363136 501915 363160
rect 501221 363102 501280 363136
rect 501314 363102 501370 363136
rect 501404 363102 501460 363136
rect 501494 363102 501550 363136
rect 501584 363102 501640 363136
rect 501674 363102 501730 363136
rect 501764 363102 501820 363136
rect 501854 363102 501915 363136
rect 501221 363094 501915 363102
rect 501221 363060 501308 363094
rect 501342 363060 501408 363094
rect 501442 363060 501508 363094
rect 501542 363060 501608 363094
rect 501642 363060 501708 363094
rect 501742 363060 501808 363094
rect 501842 363060 501915 363094
rect 501221 363046 501915 363060
rect 501221 363012 501280 363046
rect 501314 363012 501370 363046
rect 501404 363012 501460 363046
rect 501494 363012 501550 363046
rect 501584 363012 501640 363046
rect 501674 363012 501730 363046
rect 501764 363012 501820 363046
rect 501854 363012 501915 363046
rect 501221 362994 501915 363012
rect 501221 362960 501308 362994
rect 501342 362960 501408 362994
rect 501442 362960 501508 362994
rect 501542 362960 501608 362994
rect 501642 362960 501708 362994
rect 501742 362960 501808 362994
rect 501842 362960 501915 362994
rect 501221 362956 501915 362960
rect 501221 362922 501280 362956
rect 501314 362922 501370 362956
rect 501404 362922 501460 362956
rect 501494 362922 501550 362956
rect 501584 362922 501640 362956
rect 501674 362922 501730 362956
rect 501764 362922 501820 362956
rect 501854 362922 501915 362956
rect 501221 362894 501915 362922
rect 501221 362866 501308 362894
rect 501342 362866 501408 362894
rect 501221 362832 501280 362866
rect 501342 362860 501370 362866
rect 501314 362832 501370 362860
rect 501404 362860 501408 362866
rect 501442 362866 501508 362894
rect 501442 362860 501460 362866
rect 501404 362832 501460 362860
rect 501494 362860 501508 362866
rect 501542 362866 501608 362894
rect 501642 362866 501708 362894
rect 501742 362866 501808 362894
rect 501842 362866 501915 362894
rect 501542 362860 501550 362866
rect 501494 362832 501550 362860
rect 501584 362860 501608 362866
rect 501674 362860 501708 362866
rect 501764 362860 501808 362866
rect 501584 362832 501640 362860
rect 501674 362832 501730 362860
rect 501764 362832 501820 362860
rect 501854 362832 501915 362866
rect 501221 362773 501915 362832
rect 501977 363414 502049 363470
rect 501977 363380 501996 363414
rect 502030 363380 502049 363414
rect 501977 363324 502049 363380
rect 501977 363290 501996 363324
rect 502030 363290 502049 363324
rect 501977 363234 502049 363290
rect 501977 363200 501996 363234
rect 502030 363200 502049 363234
rect 501977 363144 502049 363200
rect 501977 363110 501996 363144
rect 502030 363110 502049 363144
rect 501977 363054 502049 363110
rect 501977 363020 501996 363054
rect 502030 363020 502049 363054
rect 501977 362964 502049 363020
rect 501977 362930 501996 362964
rect 502030 362930 502049 362964
rect 501977 362874 502049 362930
rect 501977 362840 501996 362874
rect 502030 362840 502049 362874
rect 501977 362784 502049 362840
rect 501087 362736 501104 362770
rect 501138 362750 501159 362770
rect 501087 362716 501106 362736
rect 501140 362716 501159 362750
rect 501087 362711 501159 362716
rect 501977 362750 501996 362784
rect 502030 362750 502049 362784
rect 501977 362711 502049 362750
rect 501087 362692 502049 362711
rect 501087 362680 501182 362692
rect 501087 362646 501104 362680
rect 501138 362658 501182 362680
rect 501216 362658 501272 362692
rect 501306 362658 501362 362692
rect 501396 362658 501452 362692
rect 501486 362658 501542 362692
rect 501576 362658 501632 362692
rect 501666 362658 501722 362692
rect 501756 362658 501812 362692
rect 501846 362658 501902 362692
rect 501936 362658 502049 362692
rect 501138 362646 502049 362658
rect 501087 362639 502049 362646
rect 502113 363600 502146 363634
rect 502180 363600 502212 363634
rect 502113 363544 502212 363600
rect 502113 363510 502146 363544
rect 502180 363510 502212 363544
rect 502113 363454 502212 363510
rect 502113 363420 502146 363454
rect 502180 363420 502212 363454
rect 502113 363364 502212 363420
rect 502113 363330 502146 363364
rect 502180 363330 502212 363364
rect 502113 363274 502212 363330
rect 502113 363240 502146 363274
rect 502180 363240 502212 363274
rect 502113 363184 502212 363240
rect 502113 363150 502146 363184
rect 502180 363150 502212 363184
rect 502113 363094 502212 363150
rect 502113 363060 502146 363094
rect 502180 363060 502212 363094
rect 502113 363004 502212 363060
rect 502113 362970 502146 363004
rect 502180 362970 502212 363004
rect 502113 362914 502212 362970
rect 502113 362880 502146 362914
rect 502180 362880 502212 362914
rect 502113 362824 502212 362880
rect 502113 362790 502146 362824
rect 502180 362790 502212 362824
rect 502113 362734 502212 362790
rect 502113 362700 502146 362734
rect 502180 362700 502212 362734
rect 502113 362644 502212 362700
rect 500924 362575 501023 362610
rect 502113 362610 502146 362644
rect 502180 362610 502212 362644
rect 502113 362575 502212 362610
rect 500924 362574 502212 362575
rect 500924 362540 500944 362574
rect 500978 362543 502212 362574
rect 500978 362540 500982 362543
rect 500924 362509 500982 362540
rect 501016 362509 501072 362543
rect 501106 362509 501162 362543
rect 501196 362509 501252 362543
rect 501286 362509 501342 362543
rect 501376 362509 501432 362543
rect 501466 362509 501522 362543
rect 501556 362509 501612 362543
rect 501646 362509 501702 362543
rect 501736 362509 501792 362543
rect 501826 362509 501882 362543
rect 501916 362509 501972 362543
rect 502006 362509 502062 362543
rect 502096 362509 502212 362543
rect 500924 362476 502212 362509
rect 502478 372987 502538 373170
rect 502478 372953 502491 372987
rect 502525 372953 502538 372987
rect 502478 372787 502538 372953
rect 502478 372753 502491 372787
rect 502525 372753 502538 372787
rect 502478 372587 502538 372753
rect 502478 372553 502491 372587
rect 502525 372553 502538 372587
rect 502478 372387 502538 372553
rect 502478 372353 502491 372387
rect 502525 372353 502538 372387
rect 502478 372187 502538 372353
rect 502478 372153 502491 372187
rect 502525 372153 502538 372187
rect 502478 371987 502538 372153
rect 502478 371953 502491 371987
rect 502525 371953 502538 371987
rect 502478 371787 502538 371953
rect 502478 371753 502491 371787
rect 502525 371753 502538 371787
rect 502478 371587 502538 371753
rect 502478 371553 502491 371587
rect 502525 371553 502538 371587
rect 502478 371387 502538 371553
rect 502478 371353 502491 371387
rect 502525 371353 502538 371387
rect 502478 371187 502538 371353
rect 502478 371153 502491 371187
rect 502525 371153 502538 371187
rect 502478 370987 502538 371153
rect 502478 370953 502491 370987
rect 502525 370953 502538 370987
rect 502478 370787 502538 370953
rect 502478 370753 502491 370787
rect 502525 370753 502538 370787
rect 502478 370587 502538 370753
rect 502478 370553 502491 370587
rect 502525 370553 502538 370587
rect 502478 370387 502538 370553
rect 502478 370353 502491 370387
rect 502525 370353 502538 370387
rect 502478 370187 502538 370353
rect 502478 370153 502491 370187
rect 502525 370153 502538 370187
rect 502478 369987 502538 370153
rect 502478 369953 502491 369987
rect 502525 369953 502538 369987
rect 502478 369787 502538 369953
rect 502478 369753 502491 369787
rect 502525 369753 502538 369787
rect 502478 369587 502538 369753
rect 502478 369553 502491 369587
rect 502525 369553 502538 369587
rect 502478 369387 502538 369553
rect 502478 369353 502491 369387
rect 502525 369353 502538 369387
rect 502478 369187 502538 369353
rect 502478 369153 502491 369187
rect 502525 369153 502538 369187
rect 502478 368987 502538 369153
rect 502478 368953 502491 368987
rect 502525 368953 502538 368987
rect 502478 368787 502538 368953
rect 502478 368753 502491 368787
rect 502525 368753 502538 368787
rect 502478 368587 502538 368753
rect 502478 368553 502491 368587
rect 502525 368553 502538 368587
rect 502478 368387 502538 368553
rect 502478 368353 502491 368387
rect 502525 368353 502538 368387
rect 502478 368187 502538 368353
rect 502478 368153 502491 368187
rect 502525 368153 502538 368187
rect 502478 367987 502538 368153
rect 502478 367953 502491 367987
rect 502525 367953 502538 367987
rect 502478 367787 502538 367953
rect 502478 367753 502491 367787
rect 502525 367753 502538 367787
rect 502478 367587 502538 367753
rect 502478 367553 502491 367587
rect 502525 367553 502538 367587
rect 502478 367387 502538 367553
rect 502478 367353 502491 367387
rect 502525 367353 502538 367387
rect 502478 367187 502538 367353
rect 502478 367153 502491 367187
rect 502525 367153 502538 367187
rect 502478 366987 502538 367153
rect 502478 366953 502491 366987
rect 502525 366953 502538 366987
rect 502478 366787 502538 366953
rect 502478 366753 502491 366787
rect 502525 366753 502538 366787
rect 502478 366587 502538 366753
rect 502478 366553 502491 366587
rect 502525 366553 502538 366587
rect 502478 366387 502538 366553
rect 502478 366353 502491 366387
rect 502525 366353 502538 366387
rect 502478 366187 502538 366353
rect 502478 366153 502491 366187
rect 502525 366153 502538 366187
rect 502478 365987 502538 366153
rect 502478 365953 502491 365987
rect 502525 365953 502538 365987
rect 502478 365787 502538 365953
rect 502478 365753 502491 365787
rect 502525 365753 502538 365787
rect 502478 365587 502538 365753
rect 502478 365553 502491 365587
rect 502525 365553 502538 365587
rect 502478 365387 502538 365553
rect 502478 365353 502491 365387
rect 502525 365353 502538 365387
rect 502478 365187 502538 365353
rect 502478 365153 502491 365187
rect 502525 365153 502538 365187
rect 502478 364987 502538 365153
rect 502478 364953 502491 364987
rect 502525 364953 502538 364987
rect 502478 364787 502538 364953
rect 502478 364753 502491 364787
rect 502525 364753 502538 364787
rect 502478 364587 502538 364753
rect 502478 364553 502491 364587
rect 502525 364553 502538 364587
rect 502478 364387 502538 364553
rect 502478 364353 502491 364387
rect 502525 364353 502538 364387
rect 502478 364187 502538 364353
rect 502478 364153 502491 364187
rect 502525 364153 502538 364187
rect 502478 363987 502538 364153
rect 502478 363953 502491 363987
rect 502525 363953 502538 363987
rect 502478 363787 502538 363953
rect 502478 363753 502491 363787
rect 502525 363753 502538 363787
rect 502478 363587 502538 363753
rect 502478 363553 502491 363587
rect 502525 363553 502538 363587
rect 502478 363387 502538 363553
rect 502478 363353 502491 363387
rect 502525 363353 502538 363387
rect 502478 363187 502538 363353
rect 502478 363153 502491 363187
rect 502525 363153 502538 363187
rect 502478 362987 502538 363153
rect 502478 362953 502491 362987
rect 502525 362953 502538 362987
rect 502478 362787 502538 362953
rect 502478 362753 502491 362787
rect 502525 362753 502538 362787
rect 502478 362587 502538 362753
rect 502478 362553 502491 362587
rect 502525 362553 502538 362587
rect 502478 362450 502538 362553
rect 504358 372987 504418 373170
rect 504358 372953 504371 372987
rect 504405 372953 504418 372987
rect 504358 372787 504418 372953
rect 504358 372753 504371 372787
rect 504405 372753 504418 372787
rect 504358 372587 504418 372753
rect 504358 372553 504371 372587
rect 504405 372553 504418 372587
rect 504358 372387 504418 372553
rect 504358 372353 504371 372387
rect 504405 372353 504418 372387
rect 504358 372187 504418 372353
rect 504358 372153 504371 372187
rect 504405 372153 504418 372187
rect 504358 371987 504418 372153
rect 504358 371953 504371 371987
rect 504405 371953 504418 371987
rect 504358 371787 504418 371953
rect 504358 371753 504371 371787
rect 504405 371753 504418 371787
rect 504358 371587 504418 371753
rect 504358 371553 504371 371587
rect 504405 371553 504418 371587
rect 504358 371387 504418 371553
rect 504358 371353 504371 371387
rect 504405 371353 504418 371387
rect 504358 371187 504418 371353
rect 504358 371153 504371 371187
rect 504405 371153 504418 371187
rect 504358 370987 504418 371153
rect 504358 370953 504371 370987
rect 504405 370953 504418 370987
rect 504358 370787 504418 370953
rect 504358 370753 504371 370787
rect 504405 370753 504418 370787
rect 504358 370587 504418 370753
rect 504358 370553 504371 370587
rect 504405 370553 504418 370587
rect 504358 370387 504418 370553
rect 504358 370353 504371 370387
rect 504405 370353 504418 370387
rect 504358 370187 504418 370353
rect 504358 370153 504371 370187
rect 504405 370153 504418 370187
rect 504358 369987 504418 370153
rect 504358 369953 504371 369987
rect 504405 369953 504418 369987
rect 504358 369787 504418 369953
rect 504358 369753 504371 369787
rect 504405 369753 504418 369787
rect 504358 369587 504418 369753
rect 504358 369553 504371 369587
rect 504405 369553 504418 369587
rect 504358 369387 504418 369553
rect 504358 369353 504371 369387
rect 504405 369353 504418 369387
rect 504358 369187 504418 369353
rect 504358 369153 504371 369187
rect 504405 369153 504418 369187
rect 504358 368987 504418 369153
rect 504358 368953 504371 368987
rect 504405 368953 504418 368987
rect 504358 368787 504418 368953
rect 504358 368753 504371 368787
rect 504405 368753 504418 368787
rect 504358 368587 504418 368753
rect 504358 368553 504371 368587
rect 504405 368553 504418 368587
rect 504358 368387 504418 368553
rect 504358 368353 504371 368387
rect 504405 368353 504418 368387
rect 504358 368187 504418 368353
rect 504358 368153 504371 368187
rect 504405 368153 504418 368187
rect 504358 367987 504418 368153
rect 504358 367953 504371 367987
rect 504405 367953 504418 367987
rect 504358 367787 504418 367953
rect 504358 367753 504371 367787
rect 504405 367753 504418 367787
rect 504358 367587 504418 367753
rect 504358 367553 504371 367587
rect 504405 367553 504418 367587
rect 504358 367387 504418 367553
rect 504358 367353 504371 367387
rect 504405 367353 504418 367387
rect 504358 367187 504418 367353
rect 504358 367153 504371 367187
rect 504405 367153 504418 367187
rect 504358 366987 504418 367153
rect 504358 366953 504371 366987
rect 504405 366953 504418 366987
rect 504358 366787 504418 366953
rect 504358 366753 504371 366787
rect 504405 366753 504418 366787
rect 504358 366587 504418 366753
rect 504358 366553 504371 366587
rect 504405 366553 504418 366587
rect 504358 366387 504418 366553
rect 504358 366353 504371 366387
rect 504405 366353 504418 366387
rect 504358 366187 504418 366353
rect 504358 366153 504371 366187
rect 504405 366153 504418 366187
rect 504358 365987 504418 366153
rect 504358 365953 504371 365987
rect 504405 365953 504418 365987
rect 504358 365787 504418 365953
rect 504358 365753 504371 365787
rect 504405 365753 504418 365787
rect 504358 365587 504418 365753
rect 504358 365553 504371 365587
rect 504405 365553 504418 365587
rect 504358 365387 504418 365553
rect 504358 365353 504371 365387
rect 504405 365353 504418 365387
rect 504358 365187 504418 365353
rect 504358 365153 504371 365187
rect 504405 365153 504418 365187
rect 504358 364987 504418 365153
rect 504358 364953 504371 364987
rect 504405 364953 504418 364987
rect 504358 364787 504418 364953
rect 504358 364753 504371 364787
rect 504405 364753 504418 364787
rect 504358 364587 504418 364753
rect 504358 364553 504371 364587
rect 504405 364553 504418 364587
rect 504358 364387 504418 364553
rect 504358 364353 504371 364387
rect 504405 364353 504418 364387
rect 504358 364187 504418 364353
rect 504358 364153 504371 364187
rect 504405 364153 504418 364187
rect 504358 363987 504418 364153
rect 504358 363953 504371 363987
rect 504405 363953 504418 363987
rect 504358 363787 504418 363953
rect 504358 363753 504371 363787
rect 504405 363753 504418 363787
rect 504358 363587 504418 363753
rect 504358 363553 504371 363587
rect 504405 363553 504418 363587
rect 504358 363387 504418 363553
rect 504358 363353 504371 363387
rect 504405 363353 504418 363387
rect 504358 363187 504418 363353
rect 504358 363153 504371 363187
rect 504405 363153 504418 363187
rect 504358 362987 504418 363153
rect 504358 362953 504371 362987
rect 504405 362953 504418 362987
rect 504358 362787 504418 362953
rect 504358 362753 504371 362787
rect 504405 362753 504418 362787
rect 504358 362587 504418 362753
rect 504358 362553 504371 362587
rect 504405 362553 504418 362587
rect 504358 362450 504418 362553
rect 504684 373124 505972 373144
rect 504684 373090 504704 373124
rect 504738 373110 505972 373124
rect 504738 373090 504742 373110
rect 504684 373076 504742 373090
rect 504776 373076 504832 373110
rect 504866 373076 504922 373110
rect 504956 373076 505012 373110
rect 505046 373076 505102 373110
rect 505136 373076 505192 373110
rect 505226 373076 505282 373110
rect 505316 373076 505372 373110
rect 505406 373076 505462 373110
rect 505496 373076 505552 373110
rect 505586 373076 505642 373110
rect 505676 373076 505732 373110
rect 505766 373076 505822 373110
rect 505856 373076 505972 373110
rect 504684 373045 505972 373076
rect 504684 373034 504783 373045
rect 504684 373000 504704 373034
rect 504738 373014 504783 373034
rect 504684 372980 504719 373000
rect 504753 372980 504783 373014
rect 505873 373014 505972 373045
rect 504684 372944 504783 372980
rect 504684 372910 504704 372944
rect 504738 372924 504783 372944
rect 504684 372890 504719 372910
rect 504753 372890 504783 372924
rect 504684 372854 504783 372890
rect 504684 372820 504704 372854
rect 504738 372834 504783 372854
rect 504684 372800 504719 372820
rect 504753 372800 504783 372834
rect 504684 372764 504783 372800
rect 504684 372730 504704 372764
rect 504738 372744 504783 372764
rect 504684 372710 504719 372730
rect 504753 372710 504783 372744
rect 504684 372674 504783 372710
rect 504684 372640 504704 372674
rect 504738 372654 504783 372674
rect 504684 372620 504719 372640
rect 504753 372620 504783 372654
rect 504684 372584 504783 372620
rect 504684 372550 504704 372584
rect 504738 372564 504783 372584
rect 504684 372530 504719 372550
rect 504753 372530 504783 372564
rect 504684 372494 504783 372530
rect 504684 372460 504704 372494
rect 504738 372474 504783 372494
rect 504684 372440 504719 372460
rect 504753 372440 504783 372474
rect 504684 372404 504783 372440
rect 504684 372370 504704 372404
rect 504738 372384 504783 372404
rect 504684 372350 504719 372370
rect 504753 372350 504783 372384
rect 504684 372314 504783 372350
rect 504684 372280 504704 372314
rect 504738 372294 504783 372314
rect 504684 372260 504719 372280
rect 504753 372260 504783 372294
rect 504684 372224 504783 372260
rect 504684 372190 504704 372224
rect 504738 372204 504783 372224
rect 504684 372170 504719 372190
rect 504753 372170 504783 372204
rect 504684 372134 504783 372170
rect 504684 372100 504704 372134
rect 504738 372114 504783 372134
rect 504684 372080 504719 372100
rect 504753 372080 504783 372114
rect 504684 372044 504783 372080
rect 504684 372010 504704 372044
rect 504738 372024 504783 372044
rect 504684 371990 504719 372010
rect 504753 371990 504783 372024
rect 504847 372962 505809 372981
rect 504847 372960 504923 372962
rect 504847 372926 504864 372960
rect 504898 372928 504923 372960
rect 504957 372928 505013 372962
rect 505047 372928 505103 372962
rect 505137 372928 505193 372962
rect 505227 372928 505283 372962
rect 505317 372928 505373 372962
rect 505407 372928 505463 372962
rect 505497 372928 505553 372962
rect 505587 372928 505643 372962
rect 505677 372928 505809 372962
rect 504898 372926 505809 372928
rect 504847 372909 505809 372926
rect 504847 372870 504919 372909
rect 504847 372836 504864 372870
rect 504898 372850 504919 372870
rect 504847 372816 504866 372836
rect 504900 372816 504919 372850
rect 505737 372884 505809 372909
rect 505737 372850 505756 372884
rect 505790 372850 505809 372884
rect 504847 372780 504919 372816
rect 504847 372746 504864 372780
rect 504898 372760 504919 372780
rect 504847 372726 504866 372746
rect 504900 372726 504919 372760
rect 504847 372690 504919 372726
rect 504847 372656 504864 372690
rect 504898 372670 504919 372690
rect 504847 372636 504866 372656
rect 504900 372636 504919 372670
rect 504847 372600 504919 372636
rect 504847 372566 504864 372600
rect 504898 372580 504919 372600
rect 504847 372546 504866 372566
rect 504900 372546 504919 372580
rect 504847 372510 504919 372546
rect 504847 372476 504864 372510
rect 504898 372490 504919 372510
rect 504847 372456 504866 372476
rect 504900 372456 504919 372490
rect 504847 372420 504919 372456
rect 504847 372386 504864 372420
rect 504898 372400 504919 372420
rect 504847 372366 504866 372386
rect 504900 372366 504919 372400
rect 504847 372330 504919 372366
rect 504847 372296 504864 372330
rect 504898 372310 504919 372330
rect 504847 372276 504866 372296
rect 504900 372276 504919 372310
rect 504847 372240 504919 372276
rect 504847 372206 504864 372240
rect 504898 372220 504919 372240
rect 504847 372186 504866 372206
rect 504900 372186 504919 372220
rect 504847 372150 504919 372186
rect 504981 372786 505675 372847
rect 504981 372752 505040 372786
rect 505074 372774 505130 372786
rect 505102 372752 505130 372774
rect 505164 372774 505220 372786
rect 505164 372752 505168 372774
rect 504981 372740 505068 372752
rect 505102 372740 505168 372752
rect 505202 372752 505220 372774
rect 505254 372774 505310 372786
rect 505254 372752 505268 372774
rect 505202 372740 505268 372752
rect 505302 372752 505310 372774
rect 505344 372774 505400 372786
rect 505434 372774 505490 372786
rect 505524 372774 505580 372786
rect 505344 372752 505368 372774
rect 505434 372752 505468 372774
rect 505524 372752 505568 372774
rect 505614 372752 505675 372786
rect 505302 372740 505368 372752
rect 505402 372740 505468 372752
rect 505502 372740 505568 372752
rect 505602 372740 505675 372752
rect 504981 372696 505675 372740
rect 504981 372662 505040 372696
rect 505074 372674 505130 372696
rect 505102 372662 505130 372674
rect 505164 372674 505220 372696
rect 505164 372662 505168 372674
rect 504981 372640 505068 372662
rect 505102 372640 505168 372662
rect 505202 372662 505220 372674
rect 505254 372674 505310 372696
rect 505254 372662 505268 372674
rect 505202 372640 505268 372662
rect 505302 372662 505310 372674
rect 505344 372674 505400 372696
rect 505434 372674 505490 372696
rect 505524 372674 505580 372696
rect 505344 372662 505368 372674
rect 505434 372662 505468 372674
rect 505524 372662 505568 372674
rect 505614 372662 505675 372696
rect 505302 372640 505368 372662
rect 505402 372640 505468 372662
rect 505502 372640 505568 372662
rect 505602 372640 505675 372662
rect 504981 372606 505675 372640
rect 504981 372572 505040 372606
rect 505074 372574 505130 372606
rect 505102 372572 505130 372574
rect 505164 372574 505220 372606
rect 505164 372572 505168 372574
rect 504981 372540 505068 372572
rect 505102 372540 505168 372572
rect 505202 372572 505220 372574
rect 505254 372574 505310 372606
rect 505254 372572 505268 372574
rect 505202 372540 505268 372572
rect 505302 372572 505310 372574
rect 505344 372574 505400 372606
rect 505434 372574 505490 372606
rect 505524 372574 505580 372606
rect 505344 372572 505368 372574
rect 505434 372572 505468 372574
rect 505524 372572 505568 372574
rect 505614 372572 505675 372606
rect 505302 372540 505368 372572
rect 505402 372540 505468 372572
rect 505502 372540 505568 372572
rect 505602 372540 505675 372572
rect 504981 372516 505675 372540
rect 504981 372482 505040 372516
rect 505074 372482 505130 372516
rect 505164 372482 505220 372516
rect 505254 372482 505310 372516
rect 505344 372482 505400 372516
rect 505434 372482 505490 372516
rect 505524 372482 505580 372516
rect 505614 372482 505675 372516
rect 504981 372474 505675 372482
rect 504981 372440 505068 372474
rect 505102 372440 505168 372474
rect 505202 372440 505268 372474
rect 505302 372440 505368 372474
rect 505402 372440 505468 372474
rect 505502 372440 505568 372474
rect 505602 372440 505675 372474
rect 504981 372426 505675 372440
rect 504981 372392 505040 372426
rect 505074 372392 505130 372426
rect 505164 372392 505220 372426
rect 505254 372392 505310 372426
rect 505344 372392 505400 372426
rect 505434 372392 505490 372426
rect 505524 372392 505580 372426
rect 505614 372392 505675 372426
rect 504981 372374 505675 372392
rect 504981 372340 505068 372374
rect 505102 372340 505168 372374
rect 505202 372340 505268 372374
rect 505302 372340 505368 372374
rect 505402 372340 505468 372374
rect 505502 372340 505568 372374
rect 505602 372340 505675 372374
rect 504981 372336 505675 372340
rect 504981 372302 505040 372336
rect 505074 372302 505130 372336
rect 505164 372302 505220 372336
rect 505254 372302 505310 372336
rect 505344 372302 505400 372336
rect 505434 372302 505490 372336
rect 505524 372302 505580 372336
rect 505614 372302 505675 372336
rect 504981 372274 505675 372302
rect 504981 372246 505068 372274
rect 505102 372246 505168 372274
rect 504981 372212 505040 372246
rect 505102 372240 505130 372246
rect 505074 372212 505130 372240
rect 505164 372240 505168 372246
rect 505202 372246 505268 372274
rect 505202 372240 505220 372246
rect 505164 372212 505220 372240
rect 505254 372240 505268 372246
rect 505302 372246 505368 372274
rect 505402 372246 505468 372274
rect 505502 372246 505568 372274
rect 505602 372246 505675 372274
rect 505302 372240 505310 372246
rect 505254 372212 505310 372240
rect 505344 372240 505368 372246
rect 505434 372240 505468 372246
rect 505524 372240 505568 372246
rect 505344 372212 505400 372240
rect 505434 372212 505490 372240
rect 505524 372212 505580 372240
rect 505614 372212 505675 372246
rect 504981 372153 505675 372212
rect 505737 372794 505809 372850
rect 505737 372760 505756 372794
rect 505790 372760 505809 372794
rect 505737 372704 505809 372760
rect 505737 372670 505756 372704
rect 505790 372670 505809 372704
rect 505737 372614 505809 372670
rect 505737 372580 505756 372614
rect 505790 372580 505809 372614
rect 505737 372524 505809 372580
rect 505737 372490 505756 372524
rect 505790 372490 505809 372524
rect 505737 372434 505809 372490
rect 505737 372400 505756 372434
rect 505790 372400 505809 372434
rect 505737 372344 505809 372400
rect 505737 372310 505756 372344
rect 505790 372310 505809 372344
rect 505737 372254 505809 372310
rect 505737 372220 505756 372254
rect 505790 372220 505809 372254
rect 505737 372164 505809 372220
rect 504847 372116 504864 372150
rect 504898 372130 504919 372150
rect 504847 372096 504866 372116
rect 504900 372096 504919 372130
rect 504847 372091 504919 372096
rect 505737 372130 505756 372164
rect 505790 372130 505809 372164
rect 505737 372091 505809 372130
rect 504847 372072 505809 372091
rect 504847 372060 504942 372072
rect 504847 372026 504864 372060
rect 504898 372038 504942 372060
rect 504976 372038 505032 372072
rect 505066 372038 505122 372072
rect 505156 372038 505212 372072
rect 505246 372038 505302 372072
rect 505336 372038 505392 372072
rect 505426 372038 505482 372072
rect 505516 372038 505572 372072
rect 505606 372038 505662 372072
rect 505696 372038 505809 372072
rect 504898 372026 505809 372038
rect 504847 372019 505809 372026
rect 505873 372980 505906 373014
rect 505940 372980 505972 373014
rect 505873 372924 505972 372980
rect 505873 372890 505906 372924
rect 505940 372890 505972 372924
rect 505873 372834 505972 372890
rect 505873 372800 505906 372834
rect 505940 372800 505972 372834
rect 505873 372744 505972 372800
rect 505873 372710 505906 372744
rect 505940 372710 505972 372744
rect 505873 372654 505972 372710
rect 505873 372620 505906 372654
rect 505940 372620 505972 372654
rect 505873 372564 505972 372620
rect 505873 372530 505906 372564
rect 505940 372530 505972 372564
rect 505873 372474 505972 372530
rect 505873 372440 505906 372474
rect 505940 372440 505972 372474
rect 505873 372384 505972 372440
rect 505873 372350 505906 372384
rect 505940 372350 505972 372384
rect 505873 372294 505972 372350
rect 505873 372260 505906 372294
rect 505940 372260 505972 372294
rect 505873 372204 505972 372260
rect 505873 372170 505906 372204
rect 505940 372170 505972 372204
rect 505873 372114 505972 372170
rect 505873 372080 505906 372114
rect 505940 372080 505972 372114
rect 505873 372024 505972 372080
rect 504684 371955 504783 371990
rect 505873 371990 505906 372024
rect 505940 371990 505972 372024
rect 505873 371955 505972 371990
rect 504684 371954 505972 371955
rect 504684 371920 504704 371954
rect 504738 371923 505972 371954
rect 504738 371920 504742 371923
rect 504684 371889 504742 371920
rect 504776 371889 504832 371923
rect 504866 371889 504922 371923
rect 504956 371889 505012 371923
rect 505046 371889 505102 371923
rect 505136 371889 505192 371923
rect 505226 371889 505282 371923
rect 505316 371889 505372 371923
rect 505406 371889 505462 371923
rect 505496 371889 505552 371923
rect 505586 371889 505642 371923
rect 505676 371889 505732 371923
rect 505766 371889 505822 371923
rect 505856 371889 505972 371923
rect 504684 371784 505972 371889
rect 504684 371750 504704 371784
rect 504738 371770 505972 371784
rect 504738 371750 504742 371770
rect 504684 371736 504742 371750
rect 504776 371736 504832 371770
rect 504866 371736 504922 371770
rect 504956 371736 505012 371770
rect 505046 371736 505102 371770
rect 505136 371736 505192 371770
rect 505226 371736 505282 371770
rect 505316 371736 505372 371770
rect 505406 371736 505462 371770
rect 505496 371736 505552 371770
rect 505586 371736 505642 371770
rect 505676 371736 505732 371770
rect 505766 371736 505822 371770
rect 505856 371736 505972 371770
rect 504684 371705 505972 371736
rect 504684 371694 504783 371705
rect 504684 371660 504704 371694
rect 504738 371674 504783 371694
rect 504684 371640 504719 371660
rect 504753 371640 504783 371674
rect 505873 371674 505972 371705
rect 504684 371604 504783 371640
rect 504684 371570 504704 371604
rect 504738 371584 504783 371604
rect 504684 371550 504719 371570
rect 504753 371550 504783 371584
rect 504684 371514 504783 371550
rect 504684 371480 504704 371514
rect 504738 371494 504783 371514
rect 504684 371460 504719 371480
rect 504753 371460 504783 371494
rect 504684 371424 504783 371460
rect 504684 371390 504704 371424
rect 504738 371404 504783 371424
rect 504684 371370 504719 371390
rect 504753 371370 504783 371404
rect 504684 371334 504783 371370
rect 504684 371300 504704 371334
rect 504738 371314 504783 371334
rect 504684 371280 504719 371300
rect 504753 371280 504783 371314
rect 504684 371244 504783 371280
rect 504684 371210 504704 371244
rect 504738 371224 504783 371244
rect 504684 371190 504719 371210
rect 504753 371190 504783 371224
rect 504684 371154 504783 371190
rect 504684 371120 504704 371154
rect 504738 371134 504783 371154
rect 504684 371100 504719 371120
rect 504753 371100 504783 371134
rect 504684 371064 504783 371100
rect 504684 371030 504704 371064
rect 504738 371044 504783 371064
rect 504684 371010 504719 371030
rect 504753 371010 504783 371044
rect 504684 370974 504783 371010
rect 504684 370940 504704 370974
rect 504738 370954 504783 370974
rect 504684 370920 504719 370940
rect 504753 370920 504783 370954
rect 504684 370884 504783 370920
rect 504684 370850 504704 370884
rect 504738 370864 504783 370884
rect 504684 370830 504719 370850
rect 504753 370830 504783 370864
rect 504684 370794 504783 370830
rect 504684 370760 504704 370794
rect 504738 370774 504783 370794
rect 504684 370740 504719 370760
rect 504753 370740 504783 370774
rect 504684 370704 504783 370740
rect 504684 370670 504704 370704
rect 504738 370684 504783 370704
rect 504684 370650 504719 370670
rect 504753 370650 504783 370684
rect 504847 371622 505809 371641
rect 504847 371620 504923 371622
rect 504847 371586 504864 371620
rect 504898 371588 504923 371620
rect 504957 371588 505013 371622
rect 505047 371588 505103 371622
rect 505137 371588 505193 371622
rect 505227 371588 505283 371622
rect 505317 371588 505373 371622
rect 505407 371588 505463 371622
rect 505497 371588 505553 371622
rect 505587 371588 505643 371622
rect 505677 371588 505809 371622
rect 504898 371586 505809 371588
rect 504847 371569 505809 371586
rect 504847 371530 504919 371569
rect 504847 371496 504864 371530
rect 504898 371510 504919 371530
rect 504847 371476 504866 371496
rect 504900 371476 504919 371510
rect 505737 371544 505809 371569
rect 505737 371510 505756 371544
rect 505790 371510 505809 371544
rect 504847 371440 504919 371476
rect 504847 371406 504864 371440
rect 504898 371420 504919 371440
rect 504847 371386 504866 371406
rect 504900 371386 504919 371420
rect 504847 371350 504919 371386
rect 504847 371316 504864 371350
rect 504898 371330 504919 371350
rect 504847 371296 504866 371316
rect 504900 371296 504919 371330
rect 504847 371260 504919 371296
rect 504847 371226 504864 371260
rect 504898 371240 504919 371260
rect 504847 371206 504866 371226
rect 504900 371206 504919 371240
rect 504847 371170 504919 371206
rect 504847 371136 504864 371170
rect 504898 371150 504919 371170
rect 504847 371116 504866 371136
rect 504900 371116 504919 371150
rect 504847 371080 504919 371116
rect 504847 371046 504864 371080
rect 504898 371060 504919 371080
rect 504847 371026 504866 371046
rect 504900 371026 504919 371060
rect 504847 370990 504919 371026
rect 504847 370956 504864 370990
rect 504898 370970 504919 370990
rect 504847 370936 504866 370956
rect 504900 370936 504919 370970
rect 504847 370900 504919 370936
rect 504847 370866 504864 370900
rect 504898 370880 504919 370900
rect 504847 370846 504866 370866
rect 504900 370846 504919 370880
rect 504847 370810 504919 370846
rect 504981 371446 505675 371507
rect 504981 371412 505040 371446
rect 505074 371434 505130 371446
rect 505102 371412 505130 371434
rect 505164 371434 505220 371446
rect 505164 371412 505168 371434
rect 504981 371400 505068 371412
rect 505102 371400 505168 371412
rect 505202 371412 505220 371434
rect 505254 371434 505310 371446
rect 505254 371412 505268 371434
rect 505202 371400 505268 371412
rect 505302 371412 505310 371434
rect 505344 371434 505400 371446
rect 505434 371434 505490 371446
rect 505524 371434 505580 371446
rect 505344 371412 505368 371434
rect 505434 371412 505468 371434
rect 505524 371412 505568 371434
rect 505614 371412 505675 371446
rect 505302 371400 505368 371412
rect 505402 371400 505468 371412
rect 505502 371400 505568 371412
rect 505602 371400 505675 371412
rect 504981 371356 505675 371400
rect 504981 371322 505040 371356
rect 505074 371334 505130 371356
rect 505102 371322 505130 371334
rect 505164 371334 505220 371356
rect 505164 371322 505168 371334
rect 504981 371300 505068 371322
rect 505102 371300 505168 371322
rect 505202 371322 505220 371334
rect 505254 371334 505310 371356
rect 505254 371322 505268 371334
rect 505202 371300 505268 371322
rect 505302 371322 505310 371334
rect 505344 371334 505400 371356
rect 505434 371334 505490 371356
rect 505524 371334 505580 371356
rect 505344 371322 505368 371334
rect 505434 371322 505468 371334
rect 505524 371322 505568 371334
rect 505614 371322 505675 371356
rect 505302 371300 505368 371322
rect 505402 371300 505468 371322
rect 505502 371300 505568 371322
rect 505602 371300 505675 371322
rect 504981 371266 505675 371300
rect 504981 371232 505040 371266
rect 505074 371234 505130 371266
rect 505102 371232 505130 371234
rect 505164 371234 505220 371266
rect 505164 371232 505168 371234
rect 504981 371200 505068 371232
rect 505102 371200 505168 371232
rect 505202 371232 505220 371234
rect 505254 371234 505310 371266
rect 505254 371232 505268 371234
rect 505202 371200 505268 371232
rect 505302 371232 505310 371234
rect 505344 371234 505400 371266
rect 505434 371234 505490 371266
rect 505524 371234 505580 371266
rect 505344 371232 505368 371234
rect 505434 371232 505468 371234
rect 505524 371232 505568 371234
rect 505614 371232 505675 371266
rect 505302 371200 505368 371232
rect 505402 371200 505468 371232
rect 505502 371200 505568 371232
rect 505602 371200 505675 371232
rect 504981 371176 505675 371200
rect 504981 371142 505040 371176
rect 505074 371142 505130 371176
rect 505164 371142 505220 371176
rect 505254 371142 505310 371176
rect 505344 371142 505400 371176
rect 505434 371142 505490 371176
rect 505524 371142 505580 371176
rect 505614 371142 505675 371176
rect 504981 371134 505675 371142
rect 504981 371100 505068 371134
rect 505102 371100 505168 371134
rect 505202 371100 505268 371134
rect 505302 371100 505368 371134
rect 505402 371100 505468 371134
rect 505502 371100 505568 371134
rect 505602 371100 505675 371134
rect 504981 371086 505675 371100
rect 504981 371052 505040 371086
rect 505074 371052 505130 371086
rect 505164 371052 505220 371086
rect 505254 371052 505310 371086
rect 505344 371052 505400 371086
rect 505434 371052 505490 371086
rect 505524 371052 505580 371086
rect 505614 371052 505675 371086
rect 504981 371034 505675 371052
rect 504981 371000 505068 371034
rect 505102 371000 505168 371034
rect 505202 371000 505268 371034
rect 505302 371000 505368 371034
rect 505402 371000 505468 371034
rect 505502 371000 505568 371034
rect 505602 371000 505675 371034
rect 504981 370996 505675 371000
rect 504981 370962 505040 370996
rect 505074 370962 505130 370996
rect 505164 370962 505220 370996
rect 505254 370962 505310 370996
rect 505344 370962 505400 370996
rect 505434 370962 505490 370996
rect 505524 370962 505580 370996
rect 505614 370962 505675 370996
rect 504981 370934 505675 370962
rect 504981 370906 505068 370934
rect 505102 370906 505168 370934
rect 504981 370872 505040 370906
rect 505102 370900 505130 370906
rect 505074 370872 505130 370900
rect 505164 370900 505168 370906
rect 505202 370906 505268 370934
rect 505202 370900 505220 370906
rect 505164 370872 505220 370900
rect 505254 370900 505268 370906
rect 505302 370906 505368 370934
rect 505402 370906 505468 370934
rect 505502 370906 505568 370934
rect 505602 370906 505675 370934
rect 505302 370900 505310 370906
rect 505254 370872 505310 370900
rect 505344 370900 505368 370906
rect 505434 370900 505468 370906
rect 505524 370900 505568 370906
rect 505344 370872 505400 370900
rect 505434 370872 505490 370900
rect 505524 370872 505580 370900
rect 505614 370872 505675 370906
rect 504981 370813 505675 370872
rect 505737 371454 505809 371510
rect 505737 371420 505756 371454
rect 505790 371420 505809 371454
rect 505737 371364 505809 371420
rect 505737 371330 505756 371364
rect 505790 371330 505809 371364
rect 505737 371274 505809 371330
rect 505737 371240 505756 371274
rect 505790 371240 505809 371274
rect 505737 371184 505809 371240
rect 505737 371150 505756 371184
rect 505790 371150 505809 371184
rect 505737 371094 505809 371150
rect 505737 371060 505756 371094
rect 505790 371060 505809 371094
rect 505737 371004 505809 371060
rect 505737 370970 505756 371004
rect 505790 370970 505809 371004
rect 505737 370914 505809 370970
rect 505737 370880 505756 370914
rect 505790 370880 505809 370914
rect 505737 370824 505809 370880
rect 504847 370776 504864 370810
rect 504898 370790 504919 370810
rect 504847 370756 504866 370776
rect 504900 370756 504919 370790
rect 504847 370751 504919 370756
rect 505737 370790 505756 370824
rect 505790 370790 505809 370824
rect 505737 370751 505809 370790
rect 504847 370732 505809 370751
rect 504847 370720 504942 370732
rect 504847 370686 504864 370720
rect 504898 370698 504942 370720
rect 504976 370698 505032 370732
rect 505066 370698 505122 370732
rect 505156 370698 505212 370732
rect 505246 370698 505302 370732
rect 505336 370698 505392 370732
rect 505426 370698 505482 370732
rect 505516 370698 505572 370732
rect 505606 370698 505662 370732
rect 505696 370698 505809 370732
rect 504898 370686 505809 370698
rect 504847 370679 505809 370686
rect 505873 371640 505906 371674
rect 505940 371640 505972 371674
rect 505873 371584 505972 371640
rect 505873 371550 505906 371584
rect 505940 371550 505972 371584
rect 505873 371494 505972 371550
rect 505873 371460 505906 371494
rect 505940 371460 505972 371494
rect 505873 371404 505972 371460
rect 505873 371370 505906 371404
rect 505940 371370 505972 371404
rect 505873 371314 505972 371370
rect 505873 371280 505906 371314
rect 505940 371280 505972 371314
rect 505873 371224 505972 371280
rect 505873 371190 505906 371224
rect 505940 371190 505972 371224
rect 505873 371134 505972 371190
rect 505873 371100 505906 371134
rect 505940 371100 505972 371134
rect 505873 371044 505972 371100
rect 505873 371010 505906 371044
rect 505940 371010 505972 371044
rect 505873 370954 505972 371010
rect 505873 370920 505906 370954
rect 505940 370920 505972 370954
rect 505873 370864 505972 370920
rect 505873 370830 505906 370864
rect 505940 370830 505972 370864
rect 505873 370774 505972 370830
rect 505873 370740 505906 370774
rect 505940 370740 505972 370774
rect 505873 370684 505972 370740
rect 504684 370615 504783 370650
rect 505873 370650 505906 370684
rect 505940 370650 505972 370684
rect 505873 370615 505972 370650
rect 504684 370614 505972 370615
rect 504684 370580 504704 370614
rect 504738 370583 505972 370614
rect 504738 370580 504742 370583
rect 504684 370549 504742 370580
rect 504776 370549 504832 370583
rect 504866 370549 504922 370583
rect 504956 370549 505012 370583
rect 505046 370549 505102 370583
rect 505136 370549 505192 370583
rect 505226 370549 505282 370583
rect 505316 370549 505372 370583
rect 505406 370549 505462 370583
rect 505496 370549 505552 370583
rect 505586 370549 505642 370583
rect 505676 370549 505732 370583
rect 505766 370549 505822 370583
rect 505856 370549 505972 370583
rect 504684 370444 505972 370549
rect 504684 370410 504704 370444
rect 504738 370430 505972 370444
rect 504738 370410 504742 370430
rect 504684 370396 504742 370410
rect 504776 370396 504832 370430
rect 504866 370396 504922 370430
rect 504956 370396 505012 370430
rect 505046 370396 505102 370430
rect 505136 370396 505192 370430
rect 505226 370396 505282 370430
rect 505316 370396 505372 370430
rect 505406 370396 505462 370430
rect 505496 370396 505552 370430
rect 505586 370396 505642 370430
rect 505676 370396 505732 370430
rect 505766 370396 505822 370430
rect 505856 370396 505972 370430
rect 504684 370365 505972 370396
rect 504684 370354 504783 370365
rect 504684 370320 504704 370354
rect 504738 370334 504783 370354
rect 504684 370300 504719 370320
rect 504753 370300 504783 370334
rect 505873 370334 505972 370365
rect 504684 370264 504783 370300
rect 504684 370230 504704 370264
rect 504738 370244 504783 370264
rect 504684 370210 504719 370230
rect 504753 370210 504783 370244
rect 504684 370174 504783 370210
rect 504684 370140 504704 370174
rect 504738 370154 504783 370174
rect 504684 370120 504719 370140
rect 504753 370120 504783 370154
rect 504684 370084 504783 370120
rect 504684 370050 504704 370084
rect 504738 370064 504783 370084
rect 504684 370030 504719 370050
rect 504753 370030 504783 370064
rect 504684 369994 504783 370030
rect 504684 369960 504704 369994
rect 504738 369974 504783 369994
rect 504684 369940 504719 369960
rect 504753 369940 504783 369974
rect 504684 369904 504783 369940
rect 504684 369870 504704 369904
rect 504738 369884 504783 369904
rect 504684 369850 504719 369870
rect 504753 369850 504783 369884
rect 504684 369814 504783 369850
rect 504684 369780 504704 369814
rect 504738 369794 504783 369814
rect 504684 369760 504719 369780
rect 504753 369760 504783 369794
rect 504684 369724 504783 369760
rect 504684 369690 504704 369724
rect 504738 369704 504783 369724
rect 504684 369670 504719 369690
rect 504753 369670 504783 369704
rect 504684 369634 504783 369670
rect 504684 369600 504704 369634
rect 504738 369614 504783 369634
rect 504684 369580 504719 369600
rect 504753 369580 504783 369614
rect 504684 369544 504783 369580
rect 504684 369510 504704 369544
rect 504738 369524 504783 369544
rect 504684 369490 504719 369510
rect 504753 369490 504783 369524
rect 504684 369454 504783 369490
rect 504684 369420 504704 369454
rect 504738 369434 504783 369454
rect 504684 369400 504719 369420
rect 504753 369400 504783 369434
rect 504684 369364 504783 369400
rect 504684 369330 504704 369364
rect 504738 369344 504783 369364
rect 504684 369310 504719 369330
rect 504753 369310 504783 369344
rect 504847 370282 505809 370301
rect 504847 370280 504923 370282
rect 504847 370246 504864 370280
rect 504898 370248 504923 370280
rect 504957 370248 505013 370282
rect 505047 370248 505103 370282
rect 505137 370248 505193 370282
rect 505227 370248 505283 370282
rect 505317 370248 505373 370282
rect 505407 370248 505463 370282
rect 505497 370248 505553 370282
rect 505587 370248 505643 370282
rect 505677 370248 505809 370282
rect 504898 370246 505809 370248
rect 504847 370229 505809 370246
rect 504847 370190 504919 370229
rect 504847 370156 504864 370190
rect 504898 370170 504919 370190
rect 504847 370136 504866 370156
rect 504900 370136 504919 370170
rect 505737 370204 505809 370229
rect 505737 370170 505756 370204
rect 505790 370170 505809 370204
rect 504847 370100 504919 370136
rect 504847 370066 504864 370100
rect 504898 370080 504919 370100
rect 504847 370046 504866 370066
rect 504900 370046 504919 370080
rect 504847 370010 504919 370046
rect 504847 369976 504864 370010
rect 504898 369990 504919 370010
rect 504847 369956 504866 369976
rect 504900 369956 504919 369990
rect 504847 369920 504919 369956
rect 504847 369886 504864 369920
rect 504898 369900 504919 369920
rect 504847 369866 504866 369886
rect 504900 369866 504919 369900
rect 504847 369830 504919 369866
rect 504847 369796 504864 369830
rect 504898 369810 504919 369830
rect 504847 369776 504866 369796
rect 504900 369776 504919 369810
rect 504847 369740 504919 369776
rect 504847 369706 504864 369740
rect 504898 369720 504919 369740
rect 504847 369686 504866 369706
rect 504900 369686 504919 369720
rect 504847 369650 504919 369686
rect 504847 369616 504864 369650
rect 504898 369630 504919 369650
rect 504847 369596 504866 369616
rect 504900 369596 504919 369630
rect 504847 369560 504919 369596
rect 504847 369526 504864 369560
rect 504898 369540 504919 369560
rect 504847 369506 504866 369526
rect 504900 369506 504919 369540
rect 504847 369470 504919 369506
rect 504981 370106 505675 370167
rect 504981 370072 505040 370106
rect 505074 370094 505130 370106
rect 505102 370072 505130 370094
rect 505164 370094 505220 370106
rect 505164 370072 505168 370094
rect 504981 370060 505068 370072
rect 505102 370060 505168 370072
rect 505202 370072 505220 370094
rect 505254 370094 505310 370106
rect 505254 370072 505268 370094
rect 505202 370060 505268 370072
rect 505302 370072 505310 370094
rect 505344 370094 505400 370106
rect 505434 370094 505490 370106
rect 505524 370094 505580 370106
rect 505344 370072 505368 370094
rect 505434 370072 505468 370094
rect 505524 370072 505568 370094
rect 505614 370072 505675 370106
rect 505302 370060 505368 370072
rect 505402 370060 505468 370072
rect 505502 370060 505568 370072
rect 505602 370060 505675 370072
rect 504981 370016 505675 370060
rect 504981 369982 505040 370016
rect 505074 369994 505130 370016
rect 505102 369982 505130 369994
rect 505164 369994 505220 370016
rect 505164 369982 505168 369994
rect 504981 369960 505068 369982
rect 505102 369960 505168 369982
rect 505202 369982 505220 369994
rect 505254 369994 505310 370016
rect 505254 369982 505268 369994
rect 505202 369960 505268 369982
rect 505302 369982 505310 369994
rect 505344 369994 505400 370016
rect 505434 369994 505490 370016
rect 505524 369994 505580 370016
rect 505344 369982 505368 369994
rect 505434 369982 505468 369994
rect 505524 369982 505568 369994
rect 505614 369982 505675 370016
rect 505302 369960 505368 369982
rect 505402 369960 505468 369982
rect 505502 369960 505568 369982
rect 505602 369960 505675 369982
rect 504981 369926 505675 369960
rect 504981 369892 505040 369926
rect 505074 369894 505130 369926
rect 505102 369892 505130 369894
rect 505164 369894 505220 369926
rect 505164 369892 505168 369894
rect 504981 369860 505068 369892
rect 505102 369860 505168 369892
rect 505202 369892 505220 369894
rect 505254 369894 505310 369926
rect 505254 369892 505268 369894
rect 505202 369860 505268 369892
rect 505302 369892 505310 369894
rect 505344 369894 505400 369926
rect 505434 369894 505490 369926
rect 505524 369894 505580 369926
rect 505344 369892 505368 369894
rect 505434 369892 505468 369894
rect 505524 369892 505568 369894
rect 505614 369892 505675 369926
rect 505302 369860 505368 369892
rect 505402 369860 505468 369892
rect 505502 369860 505568 369892
rect 505602 369860 505675 369892
rect 504981 369836 505675 369860
rect 504981 369802 505040 369836
rect 505074 369802 505130 369836
rect 505164 369802 505220 369836
rect 505254 369802 505310 369836
rect 505344 369802 505400 369836
rect 505434 369802 505490 369836
rect 505524 369802 505580 369836
rect 505614 369802 505675 369836
rect 504981 369794 505675 369802
rect 504981 369760 505068 369794
rect 505102 369760 505168 369794
rect 505202 369760 505268 369794
rect 505302 369760 505368 369794
rect 505402 369760 505468 369794
rect 505502 369760 505568 369794
rect 505602 369760 505675 369794
rect 504981 369746 505675 369760
rect 504981 369712 505040 369746
rect 505074 369712 505130 369746
rect 505164 369712 505220 369746
rect 505254 369712 505310 369746
rect 505344 369712 505400 369746
rect 505434 369712 505490 369746
rect 505524 369712 505580 369746
rect 505614 369712 505675 369746
rect 504981 369694 505675 369712
rect 504981 369660 505068 369694
rect 505102 369660 505168 369694
rect 505202 369660 505268 369694
rect 505302 369660 505368 369694
rect 505402 369660 505468 369694
rect 505502 369660 505568 369694
rect 505602 369660 505675 369694
rect 504981 369656 505675 369660
rect 504981 369622 505040 369656
rect 505074 369622 505130 369656
rect 505164 369622 505220 369656
rect 505254 369622 505310 369656
rect 505344 369622 505400 369656
rect 505434 369622 505490 369656
rect 505524 369622 505580 369656
rect 505614 369622 505675 369656
rect 504981 369594 505675 369622
rect 504981 369566 505068 369594
rect 505102 369566 505168 369594
rect 504981 369532 505040 369566
rect 505102 369560 505130 369566
rect 505074 369532 505130 369560
rect 505164 369560 505168 369566
rect 505202 369566 505268 369594
rect 505202 369560 505220 369566
rect 505164 369532 505220 369560
rect 505254 369560 505268 369566
rect 505302 369566 505368 369594
rect 505402 369566 505468 369594
rect 505502 369566 505568 369594
rect 505602 369566 505675 369594
rect 505302 369560 505310 369566
rect 505254 369532 505310 369560
rect 505344 369560 505368 369566
rect 505434 369560 505468 369566
rect 505524 369560 505568 369566
rect 505344 369532 505400 369560
rect 505434 369532 505490 369560
rect 505524 369532 505580 369560
rect 505614 369532 505675 369566
rect 504981 369473 505675 369532
rect 505737 370114 505809 370170
rect 505737 370080 505756 370114
rect 505790 370080 505809 370114
rect 505737 370024 505809 370080
rect 505737 369990 505756 370024
rect 505790 369990 505809 370024
rect 505737 369934 505809 369990
rect 505737 369900 505756 369934
rect 505790 369900 505809 369934
rect 505737 369844 505809 369900
rect 505737 369810 505756 369844
rect 505790 369810 505809 369844
rect 505737 369754 505809 369810
rect 505737 369720 505756 369754
rect 505790 369720 505809 369754
rect 505737 369664 505809 369720
rect 505737 369630 505756 369664
rect 505790 369630 505809 369664
rect 505737 369574 505809 369630
rect 505737 369540 505756 369574
rect 505790 369540 505809 369574
rect 505737 369484 505809 369540
rect 504847 369436 504864 369470
rect 504898 369450 504919 369470
rect 504847 369416 504866 369436
rect 504900 369416 504919 369450
rect 504847 369411 504919 369416
rect 505737 369450 505756 369484
rect 505790 369450 505809 369484
rect 505737 369411 505809 369450
rect 504847 369392 505809 369411
rect 504847 369380 504942 369392
rect 504847 369346 504864 369380
rect 504898 369358 504942 369380
rect 504976 369358 505032 369392
rect 505066 369358 505122 369392
rect 505156 369358 505212 369392
rect 505246 369358 505302 369392
rect 505336 369358 505392 369392
rect 505426 369358 505482 369392
rect 505516 369358 505572 369392
rect 505606 369358 505662 369392
rect 505696 369358 505809 369392
rect 504898 369346 505809 369358
rect 504847 369339 505809 369346
rect 505873 370300 505906 370334
rect 505940 370300 505972 370334
rect 505873 370244 505972 370300
rect 505873 370210 505906 370244
rect 505940 370210 505972 370244
rect 505873 370154 505972 370210
rect 505873 370120 505906 370154
rect 505940 370120 505972 370154
rect 505873 370064 505972 370120
rect 505873 370030 505906 370064
rect 505940 370030 505972 370064
rect 505873 369974 505972 370030
rect 505873 369940 505906 369974
rect 505940 369940 505972 369974
rect 505873 369884 505972 369940
rect 505873 369850 505906 369884
rect 505940 369850 505972 369884
rect 505873 369794 505972 369850
rect 505873 369760 505906 369794
rect 505940 369760 505972 369794
rect 505873 369704 505972 369760
rect 505873 369670 505906 369704
rect 505940 369670 505972 369704
rect 505873 369614 505972 369670
rect 505873 369580 505906 369614
rect 505940 369580 505972 369614
rect 505873 369524 505972 369580
rect 505873 369490 505906 369524
rect 505940 369490 505972 369524
rect 505873 369434 505972 369490
rect 505873 369400 505906 369434
rect 505940 369400 505972 369434
rect 505873 369344 505972 369400
rect 504684 369275 504783 369310
rect 505873 369310 505906 369344
rect 505940 369310 505972 369344
rect 505873 369275 505972 369310
rect 504684 369274 505972 369275
rect 504684 369240 504704 369274
rect 504738 369243 505972 369274
rect 504738 369240 504742 369243
rect 504684 369209 504742 369240
rect 504776 369209 504832 369243
rect 504866 369209 504922 369243
rect 504956 369209 505012 369243
rect 505046 369209 505102 369243
rect 505136 369209 505192 369243
rect 505226 369209 505282 369243
rect 505316 369209 505372 369243
rect 505406 369209 505462 369243
rect 505496 369209 505552 369243
rect 505586 369209 505642 369243
rect 505676 369209 505732 369243
rect 505766 369209 505822 369243
rect 505856 369209 505972 369243
rect 504684 369104 505972 369209
rect 504684 369070 504704 369104
rect 504738 369090 505972 369104
rect 504738 369070 504742 369090
rect 504684 369056 504742 369070
rect 504776 369056 504832 369090
rect 504866 369056 504922 369090
rect 504956 369056 505012 369090
rect 505046 369056 505102 369090
rect 505136 369056 505192 369090
rect 505226 369056 505282 369090
rect 505316 369056 505372 369090
rect 505406 369056 505462 369090
rect 505496 369056 505552 369090
rect 505586 369056 505642 369090
rect 505676 369056 505732 369090
rect 505766 369056 505822 369090
rect 505856 369056 505972 369090
rect 504684 369025 505972 369056
rect 504684 369014 504783 369025
rect 504684 368980 504704 369014
rect 504738 368994 504783 369014
rect 504684 368960 504719 368980
rect 504753 368960 504783 368994
rect 505873 368994 505972 369025
rect 504684 368924 504783 368960
rect 504684 368890 504704 368924
rect 504738 368904 504783 368924
rect 504684 368870 504719 368890
rect 504753 368870 504783 368904
rect 504684 368834 504783 368870
rect 504684 368800 504704 368834
rect 504738 368814 504783 368834
rect 504684 368780 504719 368800
rect 504753 368780 504783 368814
rect 504684 368744 504783 368780
rect 504684 368710 504704 368744
rect 504738 368724 504783 368744
rect 504684 368690 504719 368710
rect 504753 368690 504783 368724
rect 504684 368654 504783 368690
rect 504684 368620 504704 368654
rect 504738 368634 504783 368654
rect 504684 368600 504719 368620
rect 504753 368600 504783 368634
rect 504684 368564 504783 368600
rect 504684 368530 504704 368564
rect 504738 368544 504783 368564
rect 504684 368510 504719 368530
rect 504753 368510 504783 368544
rect 504684 368474 504783 368510
rect 504684 368440 504704 368474
rect 504738 368454 504783 368474
rect 504684 368420 504719 368440
rect 504753 368420 504783 368454
rect 504684 368384 504783 368420
rect 504684 368350 504704 368384
rect 504738 368364 504783 368384
rect 504684 368330 504719 368350
rect 504753 368330 504783 368364
rect 504684 368294 504783 368330
rect 504684 368260 504704 368294
rect 504738 368274 504783 368294
rect 504684 368240 504719 368260
rect 504753 368240 504783 368274
rect 504684 368204 504783 368240
rect 504684 368170 504704 368204
rect 504738 368184 504783 368204
rect 504684 368150 504719 368170
rect 504753 368150 504783 368184
rect 504684 368114 504783 368150
rect 504684 368080 504704 368114
rect 504738 368094 504783 368114
rect 504684 368060 504719 368080
rect 504753 368060 504783 368094
rect 504684 368024 504783 368060
rect 504684 367990 504704 368024
rect 504738 368004 504783 368024
rect 504684 367970 504719 367990
rect 504753 367970 504783 368004
rect 504847 368942 505809 368961
rect 504847 368940 504923 368942
rect 504847 368906 504864 368940
rect 504898 368908 504923 368940
rect 504957 368908 505013 368942
rect 505047 368908 505103 368942
rect 505137 368908 505193 368942
rect 505227 368908 505283 368942
rect 505317 368908 505373 368942
rect 505407 368908 505463 368942
rect 505497 368908 505553 368942
rect 505587 368908 505643 368942
rect 505677 368908 505809 368942
rect 504898 368906 505809 368908
rect 504847 368889 505809 368906
rect 504847 368850 504919 368889
rect 504847 368816 504864 368850
rect 504898 368830 504919 368850
rect 504847 368796 504866 368816
rect 504900 368796 504919 368830
rect 505737 368864 505809 368889
rect 505737 368830 505756 368864
rect 505790 368830 505809 368864
rect 504847 368760 504919 368796
rect 504847 368726 504864 368760
rect 504898 368740 504919 368760
rect 504847 368706 504866 368726
rect 504900 368706 504919 368740
rect 504847 368670 504919 368706
rect 504847 368636 504864 368670
rect 504898 368650 504919 368670
rect 504847 368616 504866 368636
rect 504900 368616 504919 368650
rect 504847 368580 504919 368616
rect 504847 368546 504864 368580
rect 504898 368560 504919 368580
rect 504847 368526 504866 368546
rect 504900 368526 504919 368560
rect 504847 368490 504919 368526
rect 504847 368456 504864 368490
rect 504898 368470 504919 368490
rect 504847 368436 504866 368456
rect 504900 368436 504919 368470
rect 504847 368400 504919 368436
rect 504847 368366 504864 368400
rect 504898 368380 504919 368400
rect 504847 368346 504866 368366
rect 504900 368346 504919 368380
rect 504847 368310 504919 368346
rect 504847 368276 504864 368310
rect 504898 368290 504919 368310
rect 504847 368256 504866 368276
rect 504900 368256 504919 368290
rect 504847 368220 504919 368256
rect 504847 368186 504864 368220
rect 504898 368200 504919 368220
rect 504847 368166 504866 368186
rect 504900 368166 504919 368200
rect 504847 368130 504919 368166
rect 504981 368766 505675 368827
rect 504981 368732 505040 368766
rect 505074 368754 505130 368766
rect 505102 368732 505130 368754
rect 505164 368754 505220 368766
rect 505164 368732 505168 368754
rect 504981 368720 505068 368732
rect 505102 368720 505168 368732
rect 505202 368732 505220 368754
rect 505254 368754 505310 368766
rect 505254 368732 505268 368754
rect 505202 368720 505268 368732
rect 505302 368732 505310 368754
rect 505344 368754 505400 368766
rect 505434 368754 505490 368766
rect 505524 368754 505580 368766
rect 505344 368732 505368 368754
rect 505434 368732 505468 368754
rect 505524 368732 505568 368754
rect 505614 368732 505675 368766
rect 505302 368720 505368 368732
rect 505402 368720 505468 368732
rect 505502 368720 505568 368732
rect 505602 368720 505675 368732
rect 504981 368676 505675 368720
rect 504981 368642 505040 368676
rect 505074 368654 505130 368676
rect 505102 368642 505130 368654
rect 505164 368654 505220 368676
rect 505164 368642 505168 368654
rect 504981 368620 505068 368642
rect 505102 368620 505168 368642
rect 505202 368642 505220 368654
rect 505254 368654 505310 368676
rect 505254 368642 505268 368654
rect 505202 368620 505268 368642
rect 505302 368642 505310 368654
rect 505344 368654 505400 368676
rect 505434 368654 505490 368676
rect 505524 368654 505580 368676
rect 505344 368642 505368 368654
rect 505434 368642 505468 368654
rect 505524 368642 505568 368654
rect 505614 368642 505675 368676
rect 505302 368620 505368 368642
rect 505402 368620 505468 368642
rect 505502 368620 505568 368642
rect 505602 368620 505675 368642
rect 504981 368586 505675 368620
rect 504981 368552 505040 368586
rect 505074 368554 505130 368586
rect 505102 368552 505130 368554
rect 505164 368554 505220 368586
rect 505164 368552 505168 368554
rect 504981 368520 505068 368552
rect 505102 368520 505168 368552
rect 505202 368552 505220 368554
rect 505254 368554 505310 368586
rect 505254 368552 505268 368554
rect 505202 368520 505268 368552
rect 505302 368552 505310 368554
rect 505344 368554 505400 368586
rect 505434 368554 505490 368586
rect 505524 368554 505580 368586
rect 505344 368552 505368 368554
rect 505434 368552 505468 368554
rect 505524 368552 505568 368554
rect 505614 368552 505675 368586
rect 505302 368520 505368 368552
rect 505402 368520 505468 368552
rect 505502 368520 505568 368552
rect 505602 368520 505675 368552
rect 504981 368496 505675 368520
rect 504981 368462 505040 368496
rect 505074 368462 505130 368496
rect 505164 368462 505220 368496
rect 505254 368462 505310 368496
rect 505344 368462 505400 368496
rect 505434 368462 505490 368496
rect 505524 368462 505580 368496
rect 505614 368462 505675 368496
rect 504981 368454 505675 368462
rect 504981 368420 505068 368454
rect 505102 368420 505168 368454
rect 505202 368420 505268 368454
rect 505302 368420 505368 368454
rect 505402 368420 505468 368454
rect 505502 368420 505568 368454
rect 505602 368420 505675 368454
rect 504981 368406 505675 368420
rect 504981 368372 505040 368406
rect 505074 368372 505130 368406
rect 505164 368372 505220 368406
rect 505254 368372 505310 368406
rect 505344 368372 505400 368406
rect 505434 368372 505490 368406
rect 505524 368372 505580 368406
rect 505614 368372 505675 368406
rect 504981 368354 505675 368372
rect 504981 368320 505068 368354
rect 505102 368320 505168 368354
rect 505202 368320 505268 368354
rect 505302 368320 505368 368354
rect 505402 368320 505468 368354
rect 505502 368320 505568 368354
rect 505602 368320 505675 368354
rect 504981 368316 505675 368320
rect 504981 368282 505040 368316
rect 505074 368282 505130 368316
rect 505164 368282 505220 368316
rect 505254 368282 505310 368316
rect 505344 368282 505400 368316
rect 505434 368282 505490 368316
rect 505524 368282 505580 368316
rect 505614 368282 505675 368316
rect 504981 368254 505675 368282
rect 504981 368226 505068 368254
rect 505102 368226 505168 368254
rect 504981 368192 505040 368226
rect 505102 368220 505130 368226
rect 505074 368192 505130 368220
rect 505164 368220 505168 368226
rect 505202 368226 505268 368254
rect 505202 368220 505220 368226
rect 505164 368192 505220 368220
rect 505254 368220 505268 368226
rect 505302 368226 505368 368254
rect 505402 368226 505468 368254
rect 505502 368226 505568 368254
rect 505602 368226 505675 368254
rect 505302 368220 505310 368226
rect 505254 368192 505310 368220
rect 505344 368220 505368 368226
rect 505434 368220 505468 368226
rect 505524 368220 505568 368226
rect 505344 368192 505400 368220
rect 505434 368192 505490 368220
rect 505524 368192 505580 368220
rect 505614 368192 505675 368226
rect 504981 368133 505675 368192
rect 505737 368774 505809 368830
rect 505737 368740 505756 368774
rect 505790 368740 505809 368774
rect 505737 368684 505809 368740
rect 505737 368650 505756 368684
rect 505790 368650 505809 368684
rect 505737 368594 505809 368650
rect 505737 368560 505756 368594
rect 505790 368560 505809 368594
rect 505737 368504 505809 368560
rect 505737 368470 505756 368504
rect 505790 368470 505809 368504
rect 505737 368414 505809 368470
rect 505737 368380 505756 368414
rect 505790 368380 505809 368414
rect 505737 368324 505809 368380
rect 505737 368290 505756 368324
rect 505790 368290 505809 368324
rect 505737 368234 505809 368290
rect 505737 368200 505756 368234
rect 505790 368200 505809 368234
rect 505737 368144 505809 368200
rect 504847 368096 504864 368130
rect 504898 368110 504919 368130
rect 504847 368076 504866 368096
rect 504900 368076 504919 368110
rect 504847 368071 504919 368076
rect 505737 368110 505756 368144
rect 505790 368110 505809 368144
rect 505737 368071 505809 368110
rect 504847 368052 505809 368071
rect 504847 368040 504942 368052
rect 504847 368006 504864 368040
rect 504898 368018 504942 368040
rect 504976 368018 505032 368052
rect 505066 368018 505122 368052
rect 505156 368018 505212 368052
rect 505246 368018 505302 368052
rect 505336 368018 505392 368052
rect 505426 368018 505482 368052
rect 505516 368018 505572 368052
rect 505606 368018 505662 368052
rect 505696 368018 505809 368052
rect 504898 368006 505809 368018
rect 504847 367999 505809 368006
rect 505873 368960 505906 368994
rect 505940 368960 505972 368994
rect 505873 368904 505972 368960
rect 505873 368870 505906 368904
rect 505940 368870 505972 368904
rect 505873 368814 505972 368870
rect 505873 368780 505906 368814
rect 505940 368780 505972 368814
rect 505873 368724 505972 368780
rect 505873 368690 505906 368724
rect 505940 368690 505972 368724
rect 505873 368634 505972 368690
rect 505873 368600 505906 368634
rect 505940 368600 505972 368634
rect 505873 368544 505972 368600
rect 505873 368510 505906 368544
rect 505940 368510 505972 368544
rect 505873 368454 505972 368510
rect 505873 368420 505906 368454
rect 505940 368420 505972 368454
rect 505873 368364 505972 368420
rect 505873 368330 505906 368364
rect 505940 368330 505972 368364
rect 505873 368274 505972 368330
rect 505873 368240 505906 368274
rect 505940 368240 505972 368274
rect 505873 368184 505972 368240
rect 505873 368150 505906 368184
rect 505940 368150 505972 368184
rect 505873 368094 505972 368150
rect 505873 368060 505906 368094
rect 505940 368060 505972 368094
rect 505873 368004 505972 368060
rect 504684 367935 504783 367970
rect 505873 367970 505906 368004
rect 505940 367970 505972 368004
rect 505873 367935 505972 367970
rect 504684 367934 505972 367935
rect 504684 367900 504704 367934
rect 504738 367903 505972 367934
rect 504738 367900 504742 367903
rect 504684 367869 504742 367900
rect 504776 367869 504832 367903
rect 504866 367869 504922 367903
rect 504956 367869 505012 367903
rect 505046 367869 505102 367903
rect 505136 367869 505192 367903
rect 505226 367869 505282 367903
rect 505316 367869 505372 367903
rect 505406 367869 505462 367903
rect 505496 367869 505552 367903
rect 505586 367869 505642 367903
rect 505676 367869 505732 367903
rect 505766 367869 505822 367903
rect 505856 367869 505972 367903
rect 504684 367764 505972 367869
rect 504684 367730 504704 367764
rect 504738 367750 505972 367764
rect 504738 367730 504742 367750
rect 504684 367716 504742 367730
rect 504776 367716 504832 367750
rect 504866 367716 504922 367750
rect 504956 367716 505012 367750
rect 505046 367716 505102 367750
rect 505136 367716 505192 367750
rect 505226 367716 505282 367750
rect 505316 367716 505372 367750
rect 505406 367716 505462 367750
rect 505496 367716 505552 367750
rect 505586 367716 505642 367750
rect 505676 367716 505732 367750
rect 505766 367716 505822 367750
rect 505856 367716 505972 367750
rect 504684 367685 505972 367716
rect 504684 367674 504783 367685
rect 504684 367640 504704 367674
rect 504738 367654 504783 367674
rect 504684 367620 504719 367640
rect 504753 367620 504783 367654
rect 505873 367654 505972 367685
rect 504684 367584 504783 367620
rect 504684 367550 504704 367584
rect 504738 367564 504783 367584
rect 504684 367530 504719 367550
rect 504753 367530 504783 367564
rect 504684 367494 504783 367530
rect 504684 367460 504704 367494
rect 504738 367474 504783 367494
rect 504684 367440 504719 367460
rect 504753 367440 504783 367474
rect 504684 367404 504783 367440
rect 504684 367370 504704 367404
rect 504738 367384 504783 367404
rect 504684 367350 504719 367370
rect 504753 367350 504783 367384
rect 504684 367314 504783 367350
rect 504684 367280 504704 367314
rect 504738 367294 504783 367314
rect 504684 367260 504719 367280
rect 504753 367260 504783 367294
rect 504684 367224 504783 367260
rect 504684 367190 504704 367224
rect 504738 367204 504783 367224
rect 504684 367170 504719 367190
rect 504753 367170 504783 367204
rect 504684 367134 504783 367170
rect 504684 367100 504704 367134
rect 504738 367114 504783 367134
rect 504684 367080 504719 367100
rect 504753 367080 504783 367114
rect 504684 367044 504783 367080
rect 504684 367010 504704 367044
rect 504738 367024 504783 367044
rect 504684 366990 504719 367010
rect 504753 366990 504783 367024
rect 504684 366954 504783 366990
rect 504684 366920 504704 366954
rect 504738 366934 504783 366954
rect 504684 366900 504719 366920
rect 504753 366900 504783 366934
rect 504684 366864 504783 366900
rect 504684 366830 504704 366864
rect 504738 366844 504783 366864
rect 504684 366810 504719 366830
rect 504753 366810 504783 366844
rect 504684 366774 504783 366810
rect 504684 366740 504704 366774
rect 504738 366754 504783 366774
rect 504684 366720 504719 366740
rect 504753 366720 504783 366754
rect 504684 366684 504783 366720
rect 504684 366650 504704 366684
rect 504738 366664 504783 366684
rect 504684 366630 504719 366650
rect 504753 366630 504783 366664
rect 504847 367602 505809 367621
rect 504847 367600 504923 367602
rect 504847 367566 504864 367600
rect 504898 367568 504923 367600
rect 504957 367568 505013 367602
rect 505047 367568 505103 367602
rect 505137 367568 505193 367602
rect 505227 367568 505283 367602
rect 505317 367568 505373 367602
rect 505407 367568 505463 367602
rect 505497 367568 505553 367602
rect 505587 367568 505643 367602
rect 505677 367568 505809 367602
rect 504898 367566 505809 367568
rect 504847 367549 505809 367566
rect 504847 367510 504919 367549
rect 504847 367476 504864 367510
rect 504898 367490 504919 367510
rect 504847 367456 504866 367476
rect 504900 367456 504919 367490
rect 505737 367524 505809 367549
rect 505737 367490 505756 367524
rect 505790 367490 505809 367524
rect 504847 367420 504919 367456
rect 504847 367386 504864 367420
rect 504898 367400 504919 367420
rect 504847 367366 504866 367386
rect 504900 367366 504919 367400
rect 504847 367330 504919 367366
rect 504847 367296 504864 367330
rect 504898 367310 504919 367330
rect 504847 367276 504866 367296
rect 504900 367276 504919 367310
rect 504847 367240 504919 367276
rect 504847 367206 504864 367240
rect 504898 367220 504919 367240
rect 504847 367186 504866 367206
rect 504900 367186 504919 367220
rect 504847 367150 504919 367186
rect 504847 367116 504864 367150
rect 504898 367130 504919 367150
rect 504847 367096 504866 367116
rect 504900 367096 504919 367130
rect 504847 367060 504919 367096
rect 504847 367026 504864 367060
rect 504898 367040 504919 367060
rect 504847 367006 504866 367026
rect 504900 367006 504919 367040
rect 504847 366970 504919 367006
rect 504847 366936 504864 366970
rect 504898 366950 504919 366970
rect 504847 366916 504866 366936
rect 504900 366916 504919 366950
rect 504847 366880 504919 366916
rect 504847 366846 504864 366880
rect 504898 366860 504919 366880
rect 504847 366826 504866 366846
rect 504900 366826 504919 366860
rect 504847 366790 504919 366826
rect 504981 367426 505675 367487
rect 504981 367392 505040 367426
rect 505074 367414 505130 367426
rect 505102 367392 505130 367414
rect 505164 367414 505220 367426
rect 505164 367392 505168 367414
rect 504981 367380 505068 367392
rect 505102 367380 505168 367392
rect 505202 367392 505220 367414
rect 505254 367414 505310 367426
rect 505254 367392 505268 367414
rect 505202 367380 505268 367392
rect 505302 367392 505310 367414
rect 505344 367414 505400 367426
rect 505434 367414 505490 367426
rect 505524 367414 505580 367426
rect 505344 367392 505368 367414
rect 505434 367392 505468 367414
rect 505524 367392 505568 367414
rect 505614 367392 505675 367426
rect 505302 367380 505368 367392
rect 505402 367380 505468 367392
rect 505502 367380 505568 367392
rect 505602 367380 505675 367392
rect 504981 367336 505675 367380
rect 504981 367302 505040 367336
rect 505074 367314 505130 367336
rect 505102 367302 505130 367314
rect 505164 367314 505220 367336
rect 505164 367302 505168 367314
rect 504981 367280 505068 367302
rect 505102 367280 505168 367302
rect 505202 367302 505220 367314
rect 505254 367314 505310 367336
rect 505254 367302 505268 367314
rect 505202 367280 505268 367302
rect 505302 367302 505310 367314
rect 505344 367314 505400 367336
rect 505434 367314 505490 367336
rect 505524 367314 505580 367336
rect 505344 367302 505368 367314
rect 505434 367302 505468 367314
rect 505524 367302 505568 367314
rect 505614 367302 505675 367336
rect 505302 367280 505368 367302
rect 505402 367280 505468 367302
rect 505502 367280 505568 367302
rect 505602 367280 505675 367302
rect 504981 367246 505675 367280
rect 504981 367212 505040 367246
rect 505074 367214 505130 367246
rect 505102 367212 505130 367214
rect 505164 367214 505220 367246
rect 505164 367212 505168 367214
rect 504981 367180 505068 367212
rect 505102 367180 505168 367212
rect 505202 367212 505220 367214
rect 505254 367214 505310 367246
rect 505254 367212 505268 367214
rect 505202 367180 505268 367212
rect 505302 367212 505310 367214
rect 505344 367214 505400 367246
rect 505434 367214 505490 367246
rect 505524 367214 505580 367246
rect 505344 367212 505368 367214
rect 505434 367212 505468 367214
rect 505524 367212 505568 367214
rect 505614 367212 505675 367246
rect 505302 367180 505368 367212
rect 505402 367180 505468 367212
rect 505502 367180 505568 367212
rect 505602 367180 505675 367212
rect 504981 367156 505675 367180
rect 504981 367122 505040 367156
rect 505074 367122 505130 367156
rect 505164 367122 505220 367156
rect 505254 367122 505310 367156
rect 505344 367122 505400 367156
rect 505434 367122 505490 367156
rect 505524 367122 505580 367156
rect 505614 367122 505675 367156
rect 504981 367114 505675 367122
rect 504981 367080 505068 367114
rect 505102 367080 505168 367114
rect 505202 367080 505268 367114
rect 505302 367080 505368 367114
rect 505402 367080 505468 367114
rect 505502 367080 505568 367114
rect 505602 367080 505675 367114
rect 504981 367066 505675 367080
rect 504981 367032 505040 367066
rect 505074 367032 505130 367066
rect 505164 367032 505220 367066
rect 505254 367032 505310 367066
rect 505344 367032 505400 367066
rect 505434 367032 505490 367066
rect 505524 367032 505580 367066
rect 505614 367032 505675 367066
rect 504981 367014 505675 367032
rect 504981 366980 505068 367014
rect 505102 366980 505168 367014
rect 505202 366980 505268 367014
rect 505302 366980 505368 367014
rect 505402 366980 505468 367014
rect 505502 366980 505568 367014
rect 505602 366980 505675 367014
rect 504981 366976 505675 366980
rect 504981 366942 505040 366976
rect 505074 366942 505130 366976
rect 505164 366942 505220 366976
rect 505254 366942 505310 366976
rect 505344 366942 505400 366976
rect 505434 366942 505490 366976
rect 505524 366942 505580 366976
rect 505614 366942 505675 366976
rect 504981 366914 505675 366942
rect 504981 366886 505068 366914
rect 505102 366886 505168 366914
rect 504981 366852 505040 366886
rect 505102 366880 505130 366886
rect 505074 366852 505130 366880
rect 505164 366880 505168 366886
rect 505202 366886 505268 366914
rect 505202 366880 505220 366886
rect 505164 366852 505220 366880
rect 505254 366880 505268 366886
rect 505302 366886 505368 366914
rect 505402 366886 505468 366914
rect 505502 366886 505568 366914
rect 505602 366886 505675 366914
rect 505302 366880 505310 366886
rect 505254 366852 505310 366880
rect 505344 366880 505368 366886
rect 505434 366880 505468 366886
rect 505524 366880 505568 366886
rect 505344 366852 505400 366880
rect 505434 366852 505490 366880
rect 505524 366852 505580 366880
rect 505614 366852 505675 366886
rect 504981 366793 505675 366852
rect 505737 367434 505809 367490
rect 505737 367400 505756 367434
rect 505790 367400 505809 367434
rect 505737 367344 505809 367400
rect 505737 367310 505756 367344
rect 505790 367310 505809 367344
rect 505737 367254 505809 367310
rect 505737 367220 505756 367254
rect 505790 367220 505809 367254
rect 505737 367164 505809 367220
rect 505737 367130 505756 367164
rect 505790 367130 505809 367164
rect 505737 367074 505809 367130
rect 505737 367040 505756 367074
rect 505790 367040 505809 367074
rect 505737 366984 505809 367040
rect 505737 366950 505756 366984
rect 505790 366950 505809 366984
rect 505737 366894 505809 366950
rect 505737 366860 505756 366894
rect 505790 366860 505809 366894
rect 505737 366804 505809 366860
rect 504847 366756 504864 366790
rect 504898 366770 504919 366790
rect 504847 366736 504866 366756
rect 504900 366736 504919 366770
rect 504847 366731 504919 366736
rect 505737 366770 505756 366804
rect 505790 366770 505809 366804
rect 505737 366731 505809 366770
rect 504847 366712 505809 366731
rect 504847 366700 504942 366712
rect 504847 366666 504864 366700
rect 504898 366678 504942 366700
rect 504976 366678 505032 366712
rect 505066 366678 505122 366712
rect 505156 366678 505212 366712
rect 505246 366678 505302 366712
rect 505336 366678 505392 366712
rect 505426 366678 505482 366712
rect 505516 366678 505572 366712
rect 505606 366678 505662 366712
rect 505696 366678 505809 366712
rect 504898 366666 505809 366678
rect 504847 366659 505809 366666
rect 505873 367620 505906 367654
rect 505940 367620 505972 367654
rect 505873 367564 505972 367620
rect 505873 367530 505906 367564
rect 505940 367530 505972 367564
rect 505873 367474 505972 367530
rect 505873 367440 505906 367474
rect 505940 367440 505972 367474
rect 505873 367384 505972 367440
rect 505873 367350 505906 367384
rect 505940 367350 505972 367384
rect 505873 367294 505972 367350
rect 505873 367260 505906 367294
rect 505940 367260 505972 367294
rect 505873 367204 505972 367260
rect 505873 367170 505906 367204
rect 505940 367170 505972 367204
rect 505873 367114 505972 367170
rect 505873 367080 505906 367114
rect 505940 367080 505972 367114
rect 505873 367024 505972 367080
rect 505873 366990 505906 367024
rect 505940 366990 505972 367024
rect 505873 366934 505972 366990
rect 505873 366900 505906 366934
rect 505940 366900 505972 366934
rect 505873 366844 505972 366900
rect 505873 366810 505906 366844
rect 505940 366810 505972 366844
rect 505873 366754 505972 366810
rect 505873 366720 505906 366754
rect 505940 366720 505972 366754
rect 505873 366664 505972 366720
rect 504684 366595 504783 366630
rect 505873 366630 505906 366664
rect 505940 366630 505972 366664
rect 505873 366595 505972 366630
rect 504684 366594 505972 366595
rect 504684 366560 504704 366594
rect 504738 366563 505972 366594
rect 504738 366560 504742 366563
rect 504684 366529 504742 366560
rect 504776 366529 504832 366563
rect 504866 366529 504922 366563
rect 504956 366529 505012 366563
rect 505046 366529 505102 366563
rect 505136 366529 505192 366563
rect 505226 366529 505282 366563
rect 505316 366529 505372 366563
rect 505406 366529 505462 366563
rect 505496 366529 505552 366563
rect 505586 366529 505642 366563
rect 505676 366529 505732 366563
rect 505766 366529 505822 366563
rect 505856 366529 505972 366563
rect 504684 366424 505972 366529
rect 504684 366390 504704 366424
rect 504738 366410 505972 366424
rect 504738 366390 504742 366410
rect 504684 366376 504742 366390
rect 504776 366376 504832 366410
rect 504866 366376 504922 366410
rect 504956 366376 505012 366410
rect 505046 366376 505102 366410
rect 505136 366376 505192 366410
rect 505226 366376 505282 366410
rect 505316 366376 505372 366410
rect 505406 366376 505462 366410
rect 505496 366376 505552 366410
rect 505586 366376 505642 366410
rect 505676 366376 505732 366410
rect 505766 366376 505822 366410
rect 505856 366376 505972 366410
rect 504684 366345 505972 366376
rect 504684 366334 504783 366345
rect 504684 366300 504704 366334
rect 504738 366314 504783 366334
rect 504684 366280 504719 366300
rect 504753 366280 504783 366314
rect 505873 366314 505972 366345
rect 504684 366244 504783 366280
rect 504684 366210 504704 366244
rect 504738 366224 504783 366244
rect 504684 366190 504719 366210
rect 504753 366190 504783 366224
rect 504684 366154 504783 366190
rect 504684 366120 504704 366154
rect 504738 366134 504783 366154
rect 504684 366100 504719 366120
rect 504753 366100 504783 366134
rect 504684 366064 504783 366100
rect 504684 366030 504704 366064
rect 504738 366044 504783 366064
rect 504684 366010 504719 366030
rect 504753 366010 504783 366044
rect 504684 365974 504783 366010
rect 504684 365940 504704 365974
rect 504738 365954 504783 365974
rect 504684 365920 504719 365940
rect 504753 365920 504783 365954
rect 504684 365884 504783 365920
rect 504684 365850 504704 365884
rect 504738 365864 504783 365884
rect 504684 365830 504719 365850
rect 504753 365830 504783 365864
rect 504684 365794 504783 365830
rect 504684 365760 504704 365794
rect 504738 365774 504783 365794
rect 504684 365740 504719 365760
rect 504753 365740 504783 365774
rect 504684 365704 504783 365740
rect 504684 365670 504704 365704
rect 504738 365684 504783 365704
rect 504684 365650 504719 365670
rect 504753 365650 504783 365684
rect 504684 365614 504783 365650
rect 504684 365580 504704 365614
rect 504738 365594 504783 365614
rect 504684 365560 504719 365580
rect 504753 365560 504783 365594
rect 504684 365524 504783 365560
rect 504684 365490 504704 365524
rect 504738 365504 504783 365524
rect 504684 365470 504719 365490
rect 504753 365470 504783 365504
rect 504684 365434 504783 365470
rect 504684 365400 504704 365434
rect 504738 365414 504783 365434
rect 504684 365380 504719 365400
rect 504753 365380 504783 365414
rect 504684 365344 504783 365380
rect 504684 365310 504704 365344
rect 504738 365324 504783 365344
rect 504684 365290 504719 365310
rect 504753 365290 504783 365324
rect 504847 366262 505809 366281
rect 504847 366260 504923 366262
rect 504847 366226 504864 366260
rect 504898 366228 504923 366260
rect 504957 366228 505013 366262
rect 505047 366228 505103 366262
rect 505137 366228 505193 366262
rect 505227 366228 505283 366262
rect 505317 366228 505373 366262
rect 505407 366228 505463 366262
rect 505497 366228 505553 366262
rect 505587 366228 505643 366262
rect 505677 366228 505809 366262
rect 504898 366226 505809 366228
rect 504847 366209 505809 366226
rect 504847 366170 504919 366209
rect 504847 366136 504864 366170
rect 504898 366150 504919 366170
rect 504847 366116 504866 366136
rect 504900 366116 504919 366150
rect 505737 366184 505809 366209
rect 505737 366150 505756 366184
rect 505790 366150 505809 366184
rect 504847 366080 504919 366116
rect 504847 366046 504864 366080
rect 504898 366060 504919 366080
rect 504847 366026 504866 366046
rect 504900 366026 504919 366060
rect 504847 365990 504919 366026
rect 504847 365956 504864 365990
rect 504898 365970 504919 365990
rect 504847 365936 504866 365956
rect 504900 365936 504919 365970
rect 504847 365900 504919 365936
rect 504847 365866 504864 365900
rect 504898 365880 504919 365900
rect 504847 365846 504866 365866
rect 504900 365846 504919 365880
rect 504847 365810 504919 365846
rect 504847 365776 504864 365810
rect 504898 365790 504919 365810
rect 504847 365756 504866 365776
rect 504900 365756 504919 365790
rect 504847 365720 504919 365756
rect 504847 365686 504864 365720
rect 504898 365700 504919 365720
rect 504847 365666 504866 365686
rect 504900 365666 504919 365700
rect 504847 365630 504919 365666
rect 504847 365596 504864 365630
rect 504898 365610 504919 365630
rect 504847 365576 504866 365596
rect 504900 365576 504919 365610
rect 504847 365540 504919 365576
rect 504847 365506 504864 365540
rect 504898 365520 504919 365540
rect 504847 365486 504866 365506
rect 504900 365486 504919 365520
rect 504847 365450 504919 365486
rect 504981 366086 505675 366147
rect 504981 366052 505040 366086
rect 505074 366074 505130 366086
rect 505102 366052 505130 366074
rect 505164 366074 505220 366086
rect 505164 366052 505168 366074
rect 504981 366040 505068 366052
rect 505102 366040 505168 366052
rect 505202 366052 505220 366074
rect 505254 366074 505310 366086
rect 505254 366052 505268 366074
rect 505202 366040 505268 366052
rect 505302 366052 505310 366074
rect 505344 366074 505400 366086
rect 505434 366074 505490 366086
rect 505524 366074 505580 366086
rect 505344 366052 505368 366074
rect 505434 366052 505468 366074
rect 505524 366052 505568 366074
rect 505614 366052 505675 366086
rect 505302 366040 505368 366052
rect 505402 366040 505468 366052
rect 505502 366040 505568 366052
rect 505602 366040 505675 366052
rect 504981 365996 505675 366040
rect 504981 365962 505040 365996
rect 505074 365974 505130 365996
rect 505102 365962 505130 365974
rect 505164 365974 505220 365996
rect 505164 365962 505168 365974
rect 504981 365940 505068 365962
rect 505102 365940 505168 365962
rect 505202 365962 505220 365974
rect 505254 365974 505310 365996
rect 505254 365962 505268 365974
rect 505202 365940 505268 365962
rect 505302 365962 505310 365974
rect 505344 365974 505400 365996
rect 505434 365974 505490 365996
rect 505524 365974 505580 365996
rect 505344 365962 505368 365974
rect 505434 365962 505468 365974
rect 505524 365962 505568 365974
rect 505614 365962 505675 365996
rect 505302 365940 505368 365962
rect 505402 365940 505468 365962
rect 505502 365940 505568 365962
rect 505602 365940 505675 365962
rect 504981 365906 505675 365940
rect 504981 365872 505040 365906
rect 505074 365874 505130 365906
rect 505102 365872 505130 365874
rect 505164 365874 505220 365906
rect 505164 365872 505168 365874
rect 504981 365840 505068 365872
rect 505102 365840 505168 365872
rect 505202 365872 505220 365874
rect 505254 365874 505310 365906
rect 505254 365872 505268 365874
rect 505202 365840 505268 365872
rect 505302 365872 505310 365874
rect 505344 365874 505400 365906
rect 505434 365874 505490 365906
rect 505524 365874 505580 365906
rect 505344 365872 505368 365874
rect 505434 365872 505468 365874
rect 505524 365872 505568 365874
rect 505614 365872 505675 365906
rect 505302 365840 505368 365872
rect 505402 365840 505468 365872
rect 505502 365840 505568 365872
rect 505602 365840 505675 365872
rect 504981 365816 505675 365840
rect 504981 365782 505040 365816
rect 505074 365782 505130 365816
rect 505164 365782 505220 365816
rect 505254 365782 505310 365816
rect 505344 365782 505400 365816
rect 505434 365782 505490 365816
rect 505524 365782 505580 365816
rect 505614 365782 505675 365816
rect 504981 365774 505675 365782
rect 504981 365740 505068 365774
rect 505102 365740 505168 365774
rect 505202 365740 505268 365774
rect 505302 365740 505368 365774
rect 505402 365740 505468 365774
rect 505502 365740 505568 365774
rect 505602 365740 505675 365774
rect 504981 365726 505675 365740
rect 504981 365692 505040 365726
rect 505074 365692 505130 365726
rect 505164 365692 505220 365726
rect 505254 365692 505310 365726
rect 505344 365692 505400 365726
rect 505434 365692 505490 365726
rect 505524 365692 505580 365726
rect 505614 365692 505675 365726
rect 504981 365674 505675 365692
rect 504981 365640 505068 365674
rect 505102 365640 505168 365674
rect 505202 365640 505268 365674
rect 505302 365640 505368 365674
rect 505402 365640 505468 365674
rect 505502 365640 505568 365674
rect 505602 365640 505675 365674
rect 504981 365636 505675 365640
rect 504981 365602 505040 365636
rect 505074 365602 505130 365636
rect 505164 365602 505220 365636
rect 505254 365602 505310 365636
rect 505344 365602 505400 365636
rect 505434 365602 505490 365636
rect 505524 365602 505580 365636
rect 505614 365602 505675 365636
rect 504981 365574 505675 365602
rect 504981 365546 505068 365574
rect 505102 365546 505168 365574
rect 504981 365512 505040 365546
rect 505102 365540 505130 365546
rect 505074 365512 505130 365540
rect 505164 365540 505168 365546
rect 505202 365546 505268 365574
rect 505202 365540 505220 365546
rect 505164 365512 505220 365540
rect 505254 365540 505268 365546
rect 505302 365546 505368 365574
rect 505402 365546 505468 365574
rect 505502 365546 505568 365574
rect 505602 365546 505675 365574
rect 505302 365540 505310 365546
rect 505254 365512 505310 365540
rect 505344 365540 505368 365546
rect 505434 365540 505468 365546
rect 505524 365540 505568 365546
rect 505344 365512 505400 365540
rect 505434 365512 505490 365540
rect 505524 365512 505580 365540
rect 505614 365512 505675 365546
rect 504981 365453 505675 365512
rect 505737 366094 505809 366150
rect 505737 366060 505756 366094
rect 505790 366060 505809 366094
rect 505737 366004 505809 366060
rect 505737 365970 505756 366004
rect 505790 365970 505809 366004
rect 505737 365914 505809 365970
rect 505737 365880 505756 365914
rect 505790 365880 505809 365914
rect 505737 365824 505809 365880
rect 505737 365790 505756 365824
rect 505790 365790 505809 365824
rect 505737 365734 505809 365790
rect 505737 365700 505756 365734
rect 505790 365700 505809 365734
rect 505737 365644 505809 365700
rect 505737 365610 505756 365644
rect 505790 365610 505809 365644
rect 505737 365554 505809 365610
rect 505737 365520 505756 365554
rect 505790 365520 505809 365554
rect 505737 365464 505809 365520
rect 504847 365416 504864 365450
rect 504898 365430 504919 365450
rect 504847 365396 504866 365416
rect 504900 365396 504919 365430
rect 504847 365391 504919 365396
rect 505737 365430 505756 365464
rect 505790 365430 505809 365464
rect 505737 365391 505809 365430
rect 504847 365372 505809 365391
rect 504847 365360 504942 365372
rect 504847 365326 504864 365360
rect 504898 365338 504942 365360
rect 504976 365338 505032 365372
rect 505066 365338 505122 365372
rect 505156 365338 505212 365372
rect 505246 365338 505302 365372
rect 505336 365338 505392 365372
rect 505426 365338 505482 365372
rect 505516 365338 505572 365372
rect 505606 365338 505662 365372
rect 505696 365338 505809 365372
rect 504898 365326 505809 365338
rect 504847 365319 505809 365326
rect 505873 366280 505906 366314
rect 505940 366280 505972 366314
rect 505873 366224 505972 366280
rect 505873 366190 505906 366224
rect 505940 366190 505972 366224
rect 505873 366134 505972 366190
rect 505873 366100 505906 366134
rect 505940 366100 505972 366134
rect 505873 366044 505972 366100
rect 505873 366010 505906 366044
rect 505940 366010 505972 366044
rect 505873 365954 505972 366010
rect 505873 365920 505906 365954
rect 505940 365920 505972 365954
rect 505873 365864 505972 365920
rect 505873 365830 505906 365864
rect 505940 365830 505972 365864
rect 505873 365774 505972 365830
rect 505873 365740 505906 365774
rect 505940 365740 505972 365774
rect 505873 365684 505972 365740
rect 505873 365650 505906 365684
rect 505940 365650 505972 365684
rect 505873 365594 505972 365650
rect 505873 365560 505906 365594
rect 505940 365560 505972 365594
rect 505873 365504 505972 365560
rect 505873 365470 505906 365504
rect 505940 365470 505972 365504
rect 505873 365414 505972 365470
rect 505873 365380 505906 365414
rect 505940 365380 505972 365414
rect 505873 365324 505972 365380
rect 504684 365255 504783 365290
rect 505873 365290 505906 365324
rect 505940 365290 505972 365324
rect 505873 365255 505972 365290
rect 504684 365254 505972 365255
rect 504684 365220 504704 365254
rect 504738 365223 505972 365254
rect 504738 365220 504742 365223
rect 504684 365189 504742 365220
rect 504776 365189 504832 365223
rect 504866 365189 504922 365223
rect 504956 365189 505012 365223
rect 505046 365189 505102 365223
rect 505136 365189 505192 365223
rect 505226 365189 505282 365223
rect 505316 365189 505372 365223
rect 505406 365189 505462 365223
rect 505496 365189 505552 365223
rect 505586 365189 505642 365223
rect 505676 365189 505732 365223
rect 505766 365189 505822 365223
rect 505856 365189 505972 365223
rect 504684 365084 505972 365189
rect 504684 365050 504704 365084
rect 504738 365070 505972 365084
rect 504738 365050 504742 365070
rect 504684 365036 504742 365050
rect 504776 365036 504832 365070
rect 504866 365036 504922 365070
rect 504956 365036 505012 365070
rect 505046 365036 505102 365070
rect 505136 365036 505192 365070
rect 505226 365036 505282 365070
rect 505316 365036 505372 365070
rect 505406 365036 505462 365070
rect 505496 365036 505552 365070
rect 505586 365036 505642 365070
rect 505676 365036 505732 365070
rect 505766 365036 505822 365070
rect 505856 365036 505972 365070
rect 504684 365005 505972 365036
rect 504684 364994 504783 365005
rect 504684 364960 504704 364994
rect 504738 364974 504783 364994
rect 504684 364940 504719 364960
rect 504753 364940 504783 364974
rect 505873 364974 505972 365005
rect 504684 364904 504783 364940
rect 504684 364870 504704 364904
rect 504738 364884 504783 364904
rect 504684 364850 504719 364870
rect 504753 364850 504783 364884
rect 504684 364814 504783 364850
rect 504684 364780 504704 364814
rect 504738 364794 504783 364814
rect 504684 364760 504719 364780
rect 504753 364760 504783 364794
rect 504684 364724 504783 364760
rect 504684 364690 504704 364724
rect 504738 364704 504783 364724
rect 504684 364670 504719 364690
rect 504753 364670 504783 364704
rect 504684 364634 504783 364670
rect 504684 364600 504704 364634
rect 504738 364614 504783 364634
rect 504684 364580 504719 364600
rect 504753 364580 504783 364614
rect 504684 364544 504783 364580
rect 504684 364510 504704 364544
rect 504738 364524 504783 364544
rect 504684 364490 504719 364510
rect 504753 364490 504783 364524
rect 504684 364454 504783 364490
rect 504684 364420 504704 364454
rect 504738 364434 504783 364454
rect 504684 364400 504719 364420
rect 504753 364400 504783 364434
rect 504684 364364 504783 364400
rect 504684 364330 504704 364364
rect 504738 364344 504783 364364
rect 504684 364310 504719 364330
rect 504753 364310 504783 364344
rect 504684 364274 504783 364310
rect 504684 364240 504704 364274
rect 504738 364254 504783 364274
rect 504684 364220 504719 364240
rect 504753 364220 504783 364254
rect 504684 364184 504783 364220
rect 504684 364150 504704 364184
rect 504738 364164 504783 364184
rect 504684 364130 504719 364150
rect 504753 364130 504783 364164
rect 504684 364094 504783 364130
rect 504684 364060 504704 364094
rect 504738 364074 504783 364094
rect 504684 364040 504719 364060
rect 504753 364040 504783 364074
rect 504684 364004 504783 364040
rect 504684 363970 504704 364004
rect 504738 363984 504783 364004
rect 504684 363950 504719 363970
rect 504753 363950 504783 363984
rect 504847 364922 505809 364941
rect 504847 364920 504923 364922
rect 504847 364886 504864 364920
rect 504898 364888 504923 364920
rect 504957 364888 505013 364922
rect 505047 364888 505103 364922
rect 505137 364888 505193 364922
rect 505227 364888 505283 364922
rect 505317 364888 505373 364922
rect 505407 364888 505463 364922
rect 505497 364888 505553 364922
rect 505587 364888 505643 364922
rect 505677 364888 505809 364922
rect 504898 364886 505809 364888
rect 504847 364869 505809 364886
rect 504847 364830 504919 364869
rect 504847 364796 504864 364830
rect 504898 364810 504919 364830
rect 504847 364776 504866 364796
rect 504900 364776 504919 364810
rect 505737 364844 505809 364869
rect 505737 364810 505756 364844
rect 505790 364810 505809 364844
rect 504847 364740 504919 364776
rect 504847 364706 504864 364740
rect 504898 364720 504919 364740
rect 504847 364686 504866 364706
rect 504900 364686 504919 364720
rect 504847 364650 504919 364686
rect 504847 364616 504864 364650
rect 504898 364630 504919 364650
rect 504847 364596 504866 364616
rect 504900 364596 504919 364630
rect 504847 364560 504919 364596
rect 504847 364526 504864 364560
rect 504898 364540 504919 364560
rect 504847 364506 504866 364526
rect 504900 364506 504919 364540
rect 504847 364470 504919 364506
rect 504847 364436 504864 364470
rect 504898 364450 504919 364470
rect 504847 364416 504866 364436
rect 504900 364416 504919 364450
rect 504847 364380 504919 364416
rect 504847 364346 504864 364380
rect 504898 364360 504919 364380
rect 504847 364326 504866 364346
rect 504900 364326 504919 364360
rect 504847 364290 504919 364326
rect 504847 364256 504864 364290
rect 504898 364270 504919 364290
rect 504847 364236 504866 364256
rect 504900 364236 504919 364270
rect 504847 364200 504919 364236
rect 504847 364166 504864 364200
rect 504898 364180 504919 364200
rect 504847 364146 504866 364166
rect 504900 364146 504919 364180
rect 504847 364110 504919 364146
rect 504981 364746 505675 364807
rect 504981 364712 505040 364746
rect 505074 364734 505130 364746
rect 505102 364712 505130 364734
rect 505164 364734 505220 364746
rect 505164 364712 505168 364734
rect 504981 364700 505068 364712
rect 505102 364700 505168 364712
rect 505202 364712 505220 364734
rect 505254 364734 505310 364746
rect 505254 364712 505268 364734
rect 505202 364700 505268 364712
rect 505302 364712 505310 364734
rect 505344 364734 505400 364746
rect 505434 364734 505490 364746
rect 505524 364734 505580 364746
rect 505344 364712 505368 364734
rect 505434 364712 505468 364734
rect 505524 364712 505568 364734
rect 505614 364712 505675 364746
rect 505302 364700 505368 364712
rect 505402 364700 505468 364712
rect 505502 364700 505568 364712
rect 505602 364700 505675 364712
rect 504981 364656 505675 364700
rect 504981 364622 505040 364656
rect 505074 364634 505130 364656
rect 505102 364622 505130 364634
rect 505164 364634 505220 364656
rect 505164 364622 505168 364634
rect 504981 364600 505068 364622
rect 505102 364600 505168 364622
rect 505202 364622 505220 364634
rect 505254 364634 505310 364656
rect 505254 364622 505268 364634
rect 505202 364600 505268 364622
rect 505302 364622 505310 364634
rect 505344 364634 505400 364656
rect 505434 364634 505490 364656
rect 505524 364634 505580 364656
rect 505344 364622 505368 364634
rect 505434 364622 505468 364634
rect 505524 364622 505568 364634
rect 505614 364622 505675 364656
rect 505302 364600 505368 364622
rect 505402 364600 505468 364622
rect 505502 364600 505568 364622
rect 505602 364600 505675 364622
rect 504981 364566 505675 364600
rect 504981 364532 505040 364566
rect 505074 364534 505130 364566
rect 505102 364532 505130 364534
rect 505164 364534 505220 364566
rect 505164 364532 505168 364534
rect 504981 364500 505068 364532
rect 505102 364500 505168 364532
rect 505202 364532 505220 364534
rect 505254 364534 505310 364566
rect 505254 364532 505268 364534
rect 505202 364500 505268 364532
rect 505302 364532 505310 364534
rect 505344 364534 505400 364566
rect 505434 364534 505490 364566
rect 505524 364534 505580 364566
rect 505344 364532 505368 364534
rect 505434 364532 505468 364534
rect 505524 364532 505568 364534
rect 505614 364532 505675 364566
rect 505302 364500 505368 364532
rect 505402 364500 505468 364532
rect 505502 364500 505568 364532
rect 505602 364500 505675 364532
rect 504981 364476 505675 364500
rect 504981 364442 505040 364476
rect 505074 364442 505130 364476
rect 505164 364442 505220 364476
rect 505254 364442 505310 364476
rect 505344 364442 505400 364476
rect 505434 364442 505490 364476
rect 505524 364442 505580 364476
rect 505614 364442 505675 364476
rect 504981 364434 505675 364442
rect 504981 364400 505068 364434
rect 505102 364400 505168 364434
rect 505202 364400 505268 364434
rect 505302 364400 505368 364434
rect 505402 364400 505468 364434
rect 505502 364400 505568 364434
rect 505602 364400 505675 364434
rect 504981 364386 505675 364400
rect 504981 364352 505040 364386
rect 505074 364352 505130 364386
rect 505164 364352 505220 364386
rect 505254 364352 505310 364386
rect 505344 364352 505400 364386
rect 505434 364352 505490 364386
rect 505524 364352 505580 364386
rect 505614 364352 505675 364386
rect 504981 364334 505675 364352
rect 504981 364300 505068 364334
rect 505102 364300 505168 364334
rect 505202 364300 505268 364334
rect 505302 364300 505368 364334
rect 505402 364300 505468 364334
rect 505502 364300 505568 364334
rect 505602 364300 505675 364334
rect 504981 364296 505675 364300
rect 504981 364262 505040 364296
rect 505074 364262 505130 364296
rect 505164 364262 505220 364296
rect 505254 364262 505310 364296
rect 505344 364262 505400 364296
rect 505434 364262 505490 364296
rect 505524 364262 505580 364296
rect 505614 364262 505675 364296
rect 504981 364234 505675 364262
rect 504981 364206 505068 364234
rect 505102 364206 505168 364234
rect 504981 364172 505040 364206
rect 505102 364200 505130 364206
rect 505074 364172 505130 364200
rect 505164 364200 505168 364206
rect 505202 364206 505268 364234
rect 505202 364200 505220 364206
rect 505164 364172 505220 364200
rect 505254 364200 505268 364206
rect 505302 364206 505368 364234
rect 505402 364206 505468 364234
rect 505502 364206 505568 364234
rect 505602 364206 505675 364234
rect 505302 364200 505310 364206
rect 505254 364172 505310 364200
rect 505344 364200 505368 364206
rect 505434 364200 505468 364206
rect 505524 364200 505568 364206
rect 505344 364172 505400 364200
rect 505434 364172 505490 364200
rect 505524 364172 505580 364200
rect 505614 364172 505675 364206
rect 504981 364113 505675 364172
rect 505737 364754 505809 364810
rect 505737 364720 505756 364754
rect 505790 364720 505809 364754
rect 505737 364664 505809 364720
rect 505737 364630 505756 364664
rect 505790 364630 505809 364664
rect 505737 364574 505809 364630
rect 505737 364540 505756 364574
rect 505790 364540 505809 364574
rect 505737 364484 505809 364540
rect 505737 364450 505756 364484
rect 505790 364450 505809 364484
rect 505737 364394 505809 364450
rect 505737 364360 505756 364394
rect 505790 364360 505809 364394
rect 505737 364304 505809 364360
rect 505737 364270 505756 364304
rect 505790 364270 505809 364304
rect 505737 364214 505809 364270
rect 505737 364180 505756 364214
rect 505790 364180 505809 364214
rect 505737 364124 505809 364180
rect 504847 364076 504864 364110
rect 504898 364090 504919 364110
rect 504847 364056 504866 364076
rect 504900 364056 504919 364090
rect 504847 364051 504919 364056
rect 505737 364090 505756 364124
rect 505790 364090 505809 364124
rect 505737 364051 505809 364090
rect 504847 364032 505809 364051
rect 504847 364020 504942 364032
rect 504847 363986 504864 364020
rect 504898 363998 504942 364020
rect 504976 363998 505032 364032
rect 505066 363998 505122 364032
rect 505156 363998 505212 364032
rect 505246 363998 505302 364032
rect 505336 363998 505392 364032
rect 505426 363998 505482 364032
rect 505516 363998 505572 364032
rect 505606 363998 505662 364032
rect 505696 363998 505809 364032
rect 504898 363986 505809 363998
rect 504847 363979 505809 363986
rect 505873 364940 505906 364974
rect 505940 364940 505972 364974
rect 505873 364884 505972 364940
rect 505873 364850 505906 364884
rect 505940 364850 505972 364884
rect 505873 364794 505972 364850
rect 505873 364760 505906 364794
rect 505940 364760 505972 364794
rect 505873 364704 505972 364760
rect 505873 364670 505906 364704
rect 505940 364670 505972 364704
rect 505873 364614 505972 364670
rect 505873 364580 505906 364614
rect 505940 364580 505972 364614
rect 505873 364524 505972 364580
rect 505873 364490 505906 364524
rect 505940 364490 505972 364524
rect 505873 364434 505972 364490
rect 505873 364400 505906 364434
rect 505940 364400 505972 364434
rect 505873 364344 505972 364400
rect 505873 364310 505906 364344
rect 505940 364310 505972 364344
rect 505873 364254 505972 364310
rect 505873 364220 505906 364254
rect 505940 364220 505972 364254
rect 505873 364164 505972 364220
rect 505873 364130 505906 364164
rect 505940 364130 505972 364164
rect 505873 364074 505972 364130
rect 505873 364040 505906 364074
rect 505940 364040 505972 364074
rect 505873 363984 505972 364040
rect 504684 363915 504783 363950
rect 505873 363950 505906 363984
rect 505940 363950 505972 363984
rect 505873 363915 505972 363950
rect 504684 363914 505972 363915
rect 504684 363880 504704 363914
rect 504738 363883 505972 363914
rect 504738 363880 504742 363883
rect 504684 363849 504742 363880
rect 504776 363849 504832 363883
rect 504866 363849 504922 363883
rect 504956 363849 505012 363883
rect 505046 363849 505102 363883
rect 505136 363849 505192 363883
rect 505226 363849 505282 363883
rect 505316 363849 505372 363883
rect 505406 363849 505462 363883
rect 505496 363849 505552 363883
rect 505586 363849 505642 363883
rect 505676 363849 505732 363883
rect 505766 363849 505822 363883
rect 505856 363849 505972 363883
rect 504684 363744 505972 363849
rect 504684 363710 504704 363744
rect 504738 363730 505972 363744
rect 504738 363710 504742 363730
rect 504684 363696 504742 363710
rect 504776 363696 504832 363730
rect 504866 363696 504922 363730
rect 504956 363696 505012 363730
rect 505046 363696 505102 363730
rect 505136 363696 505192 363730
rect 505226 363696 505282 363730
rect 505316 363696 505372 363730
rect 505406 363696 505462 363730
rect 505496 363696 505552 363730
rect 505586 363696 505642 363730
rect 505676 363696 505732 363730
rect 505766 363696 505822 363730
rect 505856 363696 505972 363730
rect 504684 363665 505972 363696
rect 504684 363654 504783 363665
rect 504684 363620 504704 363654
rect 504738 363634 504783 363654
rect 504684 363600 504719 363620
rect 504753 363600 504783 363634
rect 505873 363634 505972 363665
rect 504684 363564 504783 363600
rect 504684 363530 504704 363564
rect 504738 363544 504783 363564
rect 504684 363510 504719 363530
rect 504753 363510 504783 363544
rect 504684 363474 504783 363510
rect 504684 363440 504704 363474
rect 504738 363454 504783 363474
rect 504684 363420 504719 363440
rect 504753 363420 504783 363454
rect 504684 363384 504783 363420
rect 504684 363350 504704 363384
rect 504738 363364 504783 363384
rect 504684 363330 504719 363350
rect 504753 363330 504783 363364
rect 504684 363294 504783 363330
rect 504684 363260 504704 363294
rect 504738 363274 504783 363294
rect 504684 363240 504719 363260
rect 504753 363240 504783 363274
rect 504684 363204 504783 363240
rect 504684 363170 504704 363204
rect 504738 363184 504783 363204
rect 504684 363150 504719 363170
rect 504753 363150 504783 363184
rect 504684 363114 504783 363150
rect 504684 363080 504704 363114
rect 504738 363094 504783 363114
rect 504684 363060 504719 363080
rect 504753 363060 504783 363094
rect 504684 363024 504783 363060
rect 504684 362990 504704 363024
rect 504738 363004 504783 363024
rect 504684 362970 504719 362990
rect 504753 362970 504783 363004
rect 504684 362934 504783 362970
rect 504684 362900 504704 362934
rect 504738 362914 504783 362934
rect 504684 362880 504719 362900
rect 504753 362880 504783 362914
rect 504684 362844 504783 362880
rect 504684 362810 504704 362844
rect 504738 362824 504783 362844
rect 504684 362790 504719 362810
rect 504753 362790 504783 362824
rect 504684 362754 504783 362790
rect 504684 362720 504704 362754
rect 504738 362734 504783 362754
rect 504684 362700 504719 362720
rect 504753 362700 504783 362734
rect 504684 362664 504783 362700
rect 504684 362630 504704 362664
rect 504738 362644 504783 362664
rect 504684 362610 504719 362630
rect 504753 362610 504783 362644
rect 504847 363582 505809 363601
rect 504847 363580 504923 363582
rect 504847 363546 504864 363580
rect 504898 363548 504923 363580
rect 504957 363548 505013 363582
rect 505047 363548 505103 363582
rect 505137 363548 505193 363582
rect 505227 363548 505283 363582
rect 505317 363548 505373 363582
rect 505407 363548 505463 363582
rect 505497 363548 505553 363582
rect 505587 363548 505643 363582
rect 505677 363548 505809 363582
rect 504898 363546 505809 363548
rect 504847 363529 505809 363546
rect 504847 363490 504919 363529
rect 504847 363456 504864 363490
rect 504898 363470 504919 363490
rect 504847 363436 504866 363456
rect 504900 363436 504919 363470
rect 505737 363504 505809 363529
rect 505737 363470 505756 363504
rect 505790 363470 505809 363504
rect 504847 363400 504919 363436
rect 504847 363366 504864 363400
rect 504898 363380 504919 363400
rect 504847 363346 504866 363366
rect 504900 363346 504919 363380
rect 504847 363310 504919 363346
rect 504847 363276 504864 363310
rect 504898 363290 504919 363310
rect 504847 363256 504866 363276
rect 504900 363256 504919 363290
rect 504847 363220 504919 363256
rect 504847 363186 504864 363220
rect 504898 363200 504919 363220
rect 504847 363166 504866 363186
rect 504900 363166 504919 363200
rect 504847 363130 504919 363166
rect 504847 363096 504864 363130
rect 504898 363110 504919 363130
rect 504847 363076 504866 363096
rect 504900 363076 504919 363110
rect 504847 363040 504919 363076
rect 504847 363006 504864 363040
rect 504898 363020 504919 363040
rect 504847 362986 504866 363006
rect 504900 362986 504919 363020
rect 504847 362950 504919 362986
rect 504847 362916 504864 362950
rect 504898 362930 504919 362950
rect 504847 362896 504866 362916
rect 504900 362896 504919 362930
rect 504847 362860 504919 362896
rect 504847 362826 504864 362860
rect 504898 362840 504919 362860
rect 504847 362806 504866 362826
rect 504900 362806 504919 362840
rect 504847 362770 504919 362806
rect 504981 363406 505675 363467
rect 504981 363372 505040 363406
rect 505074 363394 505130 363406
rect 505102 363372 505130 363394
rect 505164 363394 505220 363406
rect 505164 363372 505168 363394
rect 504981 363360 505068 363372
rect 505102 363360 505168 363372
rect 505202 363372 505220 363394
rect 505254 363394 505310 363406
rect 505254 363372 505268 363394
rect 505202 363360 505268 363372
rect 505302 363372 505310 363394
rect 505344 363394 505400 363406
rect 505434 363394 505490 363406
rect 505524 363394 505580 363406
rect 505344 363372 505368 363394
rect 505434 363372 505468 363394
rect 505524 363372 505568 363394
rect 505614 363372 505675 363406
rect 505302 363360 505368 363372
rect 505402 363360 505468 363372
rect 505502 363360 505568 363372
rect 505602 363360 505675 363372
rect 504981 363316 505675 363360
rect 504981 363282 505040 363316
rect 505074 363294 505130 363316
rect 505102 363282 505130 363294
rect 505164 363294 505220 363316
rect 505164 363282 505168 363294
rect 504981 363260 505068 363282
rect 505102 363260 505168 363282
rect 505202 363282 505220 363294
rect 505254 363294 505310 363316
rect 505254 363282 505268 363294
rect 505202 363260 505268 363282
rect 505302 363282 505310 363294
rect 505344 363294 505400 363316
rect 505434 363294 505490 363316
rect 505524 363294 505580 363316
rect 505344 363282 505368 363294
rect 505434 363282 505468 363294
rect 505524 363282 505568 363294
rect 505614 363282 505675 363316
rect 505302 363260 505368 363282
rect 505402 363260 505468 363282
rect 505502 363260 505568 363282
rect 505602 363260 505675 363282
rect 504981 363226 505675 363260
rect 504981 363192 505040 363226
rect 505074 363194 505130 363226
rect 505102 363192 505130 363194
rect 505164 363194 505220 363226
rect 505164 363192 505168 363194
rect 504981 363160 505068 363192
rect 505102 363160 505168 363192
rect 505202 363192 505220 363194
rect 505254 363194 505310 363226
rect 505254 363192 505268 363194
rect 505202 363160 505268 363192
rect 505302 363192 505310 363194
rect 505344 363194 505400 363226
rect 505434 363194 505490 363226
rect 505524 363194 505580 363226
rect 505344 363192 505368 363194
rect 505434 363192 505468 363194
rect 505524 363192 505568 363194
rect 505614 363192 505675 363226
rect 505302 363160 505368 363192
rect 505402 363160 505468 363192
rect 505502 363160 505568 363192
rect 505602 363160 505675 363192
rect 504981 363136 505675 363160
rect 504981 363102 505040 363136
rect 505074 363102 505130 363136
rect 505164 363102 505220 363136
rect 505254 363102 505310 363136
rect 505344 363102 505400 363136
rect 505434 363102 505490 363136
rect 505524 363102 505580 363136
rect 505614 363102 505675 363136
rect 504981 363094 505675 363102
rect 504981 363060 505068 363094
rect 505102 363060 505168 363094
rect 505202 363060 505268 363094
rect 505302 363060 505368 363094
rect 505402 363060 505468 363094
rect 505502 363060 505568 363094
rect 505602 363060 505675 363094
rect 504981 363046 505675 363060
rect 504981 363012 505040 363046
rect 505074 363012 505130 363046
rect 505164 363012 505220 363046
rect 505254 363012 505310 363046
rect 505344 363012 505400 363046
rect 505434 363012 505490 363046
rect 505524 363012 505580 363046
rect 505614 363012 505675 363046
rect 504981 362994 505675 363012
rect 504981 362960 505068 362994
rect 505102 362960 505168 362994
rect 505202 362960 505268 362994
rect 505302 362960 505368 362994
rect 505402 362960 505468 362994
rect 505502 362960 505568 362994
rect 505602 362960 505675 362994
rect 504981 362956 505675 362960
rect 504981 362922 505040 362956
rect 505074 362922 505130 362956
rect 505164 362922 505220 362956
rect 505254 362922 505310 362956
rect 505344 362922 505400 362956
rect 505434 362922 505490 362956
rect 505524 362922 505580 362956
rect 505614 362922 505675 362956
rect 504981 362894 505675 362922
rect 504981 362866 505068 362894
rect 505102 362866 505168 362894
rect 504981 362832 505040 362866
rect 505102 362860 505130 362866
rect 505074 362832 505130 362860
rect 505164 362860 505168 362866
rect 505202 362866 505268 362894
rect 505202 362860 505220 362866
rect 505164 362832 505220 362860
rect 505254 362860 505268 362866
rect 505302 362866 505368 362894
rect 505402 362866 505468 362894
rect 505502 362866 505568 362894
rect 505602 362866 505675 362894
rect 505302 362860 505310 362866
rect 505254 362832 505310 362860
rect 505344 362860 505368 362866
rect 505434 362860 505468 362866
rect 505524 362860 505568 362866
rect 505344 362832 505400 362860
rect 505434 362832 505490 362860
rect 505524 362832 505580 362860
rect 505614 362832 505675 362866
rect 504981 362773 505675 362832
rect 505737 363414 505809 363470
rect 505737 363380 505756 363414
rect 505790 363380 505809 363414
rect 505737 363324 505809 363380
rect 505737 363290 505756 363324
rect 505790 363290 505809 363324
rect 505737 363234 505809 363290
rect 505737 363200 505756 363234
rect 505790 363200 505809 363234
rect 505737 363144 505809 363200
rect 505737 363110 505756 363144
rect 505790 363110 505809 363144
rect 505737 363054 505809 363110
rect 505737 363020 505756 363054
rect 505790 363020 505809 363054
rect 505737 362964 505809 363020
rect 505737 362930 505756 362964
rect 505790 362930 505809 362964
rect 505737 362874 505809 362930
rect 505737 362840 505756 362874
rect 505790 362840 505809 362874
rect 505737 362784 505809 362840
rect 504847 362736 504864 362770
rect 504898 362750 504919 362770
rect 504847 362716 504866 362736
rect 504900 362716 504919 362750
rect 504847 362711 504919 362716
rect 505737 362750 505756 362784
rect 505790 362750 505809 362784
rect 505737 362711 505809 362750
rect 504847 362692 505809 362711
rect 504847 362680 504942 362692
rect 504847 362646 504864 362680
rect 504898 362658 504942 362680
rect 504976 362658 505032 362692
rect 505066 362658 505122 362692
rect 505156 362658 505212 362692
rect 505246 362658 505302 362692
rect 505336 362658 505392 362692
rect 505426 362658 505482 362692
rect 505516 362658 505572 362692
rect 505606 362658 505662 362692
rect 505696 362658 505809 362692
rect 504898 362646 505809 362658
rect 504847 362639 505809 362646
rect 505873 363600 505906 363634
rect 505940 363600 505972 363634
rect 505873 363544 505972 363600
rect 505873 363510 505906 363544
rect 505940 363510 505972 363544
rect 505873 363454 505972 363510
rect 505873 363420 505906 363454
rect 505940 363420 505972 363454
rect 505873 363364 505972 363420
rect 505873 363330 505906 363364
rect 505940 363330 505972 363364
rect 505873 363274 505972 363330
rect 505873 363240 505906 363274
rect 505940 363240 505972 363274
rect 505873 363184 505972 363240
rect 505873 363150 505906 363184
rect 505940 363150 505972 363184
rect 505873 363094 505972 363150
rect 505873 363060 505906 363094
rect 505940 363060 505972 363094
rect 505873 363004 505972 363060
rect 505873 362970 505906 363004
rect 505940 362970 505972 363004
rect 505873 362914 505972 362970
rect 505873 362880 505906 362914
rect 505940 362880 505972 362914
rect 505873 362824 505972 362880
rect 505873 362790 505906 362824
rect 505940 362790 505972 362824
rect 505873 362734 505972 362790
rect 505873 362700 505906 362734
rect 505940 362700 505972 362734
rect 505873 362644 505972 362700
rect 504684 362575 504783 362610
rect 505873 362610 505906 362644
rect 505940 362610 505972 362644
rect 505873 362575 505972 362610
rect 504684 362574 505972 362575
rect 504684 362540 504704 362574
rect 504738 362543 505972 362574
rect 504738 362540 504742 362543
rect 504684 362509 504742 362540
rect 504776 362509 504832 362543
rect 504866 362509 504922 362543
rect 504956 362509 505012 362543
rect 505046 362509 505102 362543
rect 505136 362509 505192 362543
rect 505226 362509 505282 362543
rect 505316 362509 505372 362543
rect 505406 362509 505462 362543
rect 505496 362509 505552 362543
rect 505586 362509 505642 362543
rect 505676 362509 505732 362543
rect 505766 362509 505822 362543
rect 505856 362509 505972 362543
rect 504684 362476 505972 362509
rect 506238 372987 506298 373170
rect 506238 372953 506251 372987
rect 506285 372953 506298 372987
rect 506238 372787 506298 372953
rect 506238 372753 506251 372787
rect 506285 372753 506298 372787
rect 506238 372587 506298 372753
rect 506238 372553 506251 372587
rect 506285 372553 506298 372587
rect 506238 372387 506298 372553
rect 506238 372353 506251 372387
rect 506285 372353 506298 372387
rect 506238 372187 506298 372353
rect 506238 372153 506251 372187
rect 506285 372153 506298 372187
rect 506238 371987 506298 372153
rect 506238 371953 506251 371987
rect 506285 371953 506298 371987
rect 506238 371787 506298 371953
rect 506238 371753 506251 371787
rect 506285 371753 506298 371787
rect 506238 371587 506298 371753
rect 506238 371553 506251 371587
rect 506285 371553 506298 371587
rect 506238 371387 506298 371553
rect 506238 371353 506251 371387
rect 506285 371353 506298 371387
rect 506238 371187 506298 371353
rect 506238 371153 506251 371187
rect 506285 371153 506298 371187
rect 506238 370987 506298 371153
rect 506238 370953 506251 370987
rect 506285 370953 506298 370987
rect 506238 370787 506298 370953
rect 506238 370753 506251 370787
rect 506285 370753 506298 370787
rect 506238 370587 506298 370753
rect 506238 370553 506251 370587
rect 506285 370553 506298 370587
rect 506238 370387 506298 370553
rect 506238 370353 506251 370387
rect 506285 370353 506298 370387
rect 506238 370187 506298 370353
rect 506238 370153 506251 370187
rect 506285 370153 506298 370187
rect 506238 369987 506298 370153
rect 506238 369953 506251 369987
rect 506285 369953 506298 369987
rect 506238 369787 506298 369953
rect 506238 369753 506251 369787
rect 506285 369753 506298 369787
rect 506238 369587 506298 369753
rect 506238 369553 506251 369587
rect 506285 369553 506298 369587
rect 506238 369387 506298 369553
rect 506238 369353 506251 369387
rect 506285 369353 506298 369387
rect 506238 369187 506298 369353
rect 506238 369153 506251 369187
rect 506285 369153 506298 369187
rect 506238 368987 506298 369153
rect 506238 368953 506251 368987
rect 506285 368953 506298 368987
rect 506238 368787 506298 368953
rect 506238 368753 506251 368787
rect 506285 368753 506298 368787
rect 506238 368587 506298 368753
rect 506238 368553 506251 368587
rect 506285 368553 506298 368587
rect 506238 368387 506298 368553
rect 506238 368353 506251 368387
rect 506285 368353 506298 368387
rect 506238 368187 506298 368353
rect 506238 368153 506251 368187
rect 506285 368153 506298 368187
rect 506238 367987 506298 368153
rect 506238 367953 506251 367987
rect 506285 367953 506298 367987
rect 506238 367787 506298 367953
rect 506238 367753 506251 367787
rect 506285 367753 506298 367787
rect 506238 367587 506298 367753
rect 506238 367553 506251 367587
rect 506285 367553 506298 367587
rect 506238 367387 506298 367553
rect 506238 367353 506251 367387
rect 506285 367353 506298 367387
rect 506238 367187 506298 367353
rect 506238 367153 506251 367187
rect 506285 367153 506298 367187
rect 506238 366987 506298 367153
rect 506238 366953 506251 366987
rect 506285 366953 506298 366987
rect 506238 366787 506298 366953
rect 506238 366753 506251 366787
rect 506285 366753 506298 366787
rect 506238 366587 506298 366753
rect 506238 366553 506251 366587
rect 506285 366553 506298 366587
rect 506238 366387 506298 366553
rect 506238 366353 506251 366387
rect 506285 366353 506298 366387
rect 506238 366187 506298 366353
rect 506238 366153 506251 366187
rect 506285 366153 506298 366187
rect 506238 365987 506298 366153
rect 506238 365953 506251 365987
rect 506285 365953 506298 365987
rect 506238 365787 506298 365953
rect 506238 365753 506251 365787
rect 506285 365753 506298 365787
rect 506238 365587 506298 365753
rect 506238 365553 506251 365587
rect 506285 365553 506298 365587
rect 506238 365387 506298 365553
rect 506238 365353 506251 365387
rect 506285 365353 506298 365387
rect 506238 365187 506298 365353
rect 506238 365153 506251 365187
rect 506285 365153 506298 365187
rect 506238 364987 506298 365153
rect 506238 364953 506251 364987
rect 506285 364953 506298 364987
rect 506238 364787 506298 364953
rect 506238 364753 506251 364787
rect 506285 364753 506298 364787
rect 506238 364587 506298 364753
rect 506238 364553 506251 364587
rect 506285 364553 506298 364587
rect 506238 364387 506298 364553
rect 506238 364353 506251 364387
rect 506285 364353 506298 364387
rect 506238 364187 506298 364353
rect 506238 364153 506251 364187
rect 506285 364153 506298 364187
rect 506238 363987 506298 364153
rect 506238 363953 506251 363987
rect 506285 363953 506298 363987
rect 506238 363787 506298 363953
rect 506238 363753 506251 363787
rect 506285 363753 506298 363787
rect 506238 363587 506298 363753
rect 506238 363553 506251 363587
rect 506285 363553 506298 363587
rect 506238 363387 506298 363553
rect 506238 363353 506251 363387
rect 506285 363353 506298 363387
rect 506238 363187 506298 363353
rect 506238 363153 506251 363187
rect 506285 363153 506298 363187
rect 506238 362987 506298 363153
rect 506238 362953 506251 362987
rect 506285 362953 506298 362987
rect 506238 362787 506298 362953
rect 506238 362753 506251 362787
rect 506285 362753 506298 362787
rect 506238 362587 506298 362753
rect 506238 362553 506251 362587
rect 506285 362553 506298 362587
rect 506238 362450 506298 362553
rect 508118 372987 508178 373170
rect 508118 372953 508131 372987
rect 508165 372953 508178 372987
rect 508118 372787 508178 372953
rect 508118 372753 508131 372787
rect 508165 372753 508178 372787
rect 508118 372587 508178 372753
rect 508118 372553 508131 372587
rect 508165 372553 508178 372587
rect 508118 372387 508178 372553
rect 508118 372353 508131 372387
rect 508165 372353 508178 372387
rect 508118 372187 508178 372353
rect 508118 372153 508131 372187
rect 508165 372153 508178 372187
rect 508118 371987 508178 372153
rect 508118 371953 508131 371987
rect 508165 371953 508178 371987
rect 508118 371787 508178 371953
rect 508118 371753 508131 371787
rect 508165 371753 508178 371787
rect 508118 371587 508178 371753
rect 508118 371553 508131 371587
rect 508165 371553 508178 371587
rect 508118 371387 508178 371553
rect 508118 371353 508131 371387
rect 508165 371353 508178 371387
rect 508118 371187 508178 371353
rect 508118 371153 508131 371187
rect 508165 371153 508178 371187
rect 508118 370987 508178 371153
rect 508118 370953 508131 370987
rect 508165 370953 508178 370987
rect 508118 370787 508178 370953
rect 508118 370753 508131 370787
rect 508165 370753 508178 370787
rect 508118 370587 508178 370753
rect 508118 370553 508131 370587
rect 508165 370553 508178 370587
rect 508118 370387 508178 370553
rect 508118 370353 508131 370387
rect 508165 370353 508178 370387
rect 508118 370187 508178 370353
rect 508118 370153 508131 370187
rect 508165 370153 508178 370187
rect 508118 369987 508178 370153
rect 508118 369953 508131 369987
rect 508165 369953 508178 369987
rect 508118 369787 508178 369953
rect 508118 369753 508131 369787
rect 508165 369753 508178 369787
rect 508118 369587 508178 369753
rect 508118 369553 508131 369587
rect 508165 369553 508178 369587
rect 508118 369387 508178 369553
rect 508118 369353 508131 369387
rect 508165 369353 508178 369387
rect 508118 369187 508178 369353
rect 508118 369153 508131 369187
rect 508165 369153 508178 369187
rect 508118 368987 508178 369153
rect 508118 368953 508131 368987
rect 508165 368953 508178 368987
rect 508118 368787 508178 368953
rect 508118 368753 508131 368787
rect 508165 368753 508178 368787
rect 508118 368587 508178 368753
rect 508118 368553 508131 368587
rect 508165 368553 508178 368587
rect 508118 368387 508178 368553
rect 508118 368353 508131 368387
rect 508165 368353 508178 368387
rect 508118 368187 508178 368353
rect 508118 368153 508131 368187
rect 508165 368153 508178 368187
rect 508118 367987 508178 368153
rect 508118 367953 508131 367987
rect 508165 367953 508178 367987
rect 508118 367787 508178 367953
rect 508118 367753 508131 367787
rect 508165 367753 508178 367787
rect 508118 367587 508178 367753
rect 508118 367553 508131 367587
rect 508165 367553 508178 367587
rect 508118 367387 508178 367553
rect 508118 367353 508131 367387
rect 508165 367353 508178 367387
rect 508118 367187 508178 367353
rect 508118 367153 508131 367187
rect 508165 367153 508178 367187
rect 508118 366987 508178 367153
rect 508118 366953 508131 366987
rect 508165 366953 508178 366987
rect 508118 366787 508178 366953
rect 508118 366753 508131 366787
rect 508165 366753 508178 366787
rect 508118 366587 508178 366753
rect 508118 366553 508131 366587
rect 508165 366553 508178 366587
rect 508118 366387 508178 366553
rect 508118 366353 508131 366387
rect 508165 366353 508178 366387
rect 508118 366187 508178 366353
rect 508118 366153 508131 366187
rect 508165 366153 508178 366187
rect 508118 365987 508178 366153
rect 508118 365953 508131 365987
rect 508165 365953 508178 365987
rect 508118 365787 508178 365953
rect 508118 365753 508131 365787
rect 508165 365753 508178 365787
rect 508118 365587 508178 365753
rect 508118 365553 508131 365587
rect 508165 365553 508178 365587
rect 508118 365387 508178 365553
rect 508118 365353 508131 365387
rect 508165 365353 508178 365387
rect 508118 365187 508178 365353
rect 508118 365153 508131 365187
rect 508165 365153 508178 365187
rect 508118 364987 508178 365153
rect 508118 364953 508131 364987
rect 508165 364953 508178 364987
rect 508118 364787 508178 364953
rect 508118 364753 508131 364787
rect 508165 364753 508178 364787
rect 508118 364587 508178 364753
rect 508118 364553 508131 364587
rect 508165 364553 508178 364587
rect 508118 364387 508178 364553
rect 508118 364353 508131 364387
rect 508165 364353 508178 364387
rect 508118 364187 508178 364353
rect 508118 364153 508131 364187
rect 508165 364153 508178 364187
rect 508118 363987 508178 364153
rect 508118 363953 508131 363987
rect 508165 363953 508178 363987
rect 508118 363787 508178 363953
rect 508118 363753 508131 363787
rect 508165 363753 508178 363787
rect 508118 363587 508178 363753
rect 508118 363553 508131 363587
rect 508165 363553 508178 363587
rect 508118 363387 508178 363553
rect 508118 363353 508131 363387
rect 508165 363353 508178 363387
rect 508118 363187 508178 363353
rect 508118 363153 508131 363187
rect 508165 363153 508178 363187
rect 508118 362987 508178 363153
rect 508118 362953 508131 362987
rect 508165 362953 508178 362987
rect 508118 362787 508178 362953
rect 508118 362753 508131 362787
rect 508165 362753 508178 362787
rect 508118 362587 508178 362753
rect 508118 362553 508131 362587
rect 508165 362553 508178 362587
rect 508118 362450 508178 362553
rect 508444 373124 509732 373144
rect 508444 373090 508464 373124
rect 508498 373110 509732 373124
rect 508498 373090 508502 373110
rect 508444 373076 508502 373090
rect 508536 373076 508592 373110
rect 508626 373076 508682 373110
rect 508716 373076 508772 373110
rect 508806 373076 508862 373110
rect 508896 373076 508952 373110
rect 508986 373076 509042 373110
rect 509076 373076 509132 373110
rect 509166 373076 509222 373110
rect 509256 373076 509312 373110
rect 509346 373076 509402 373110
rect 509436 373076 509492 373110
rect 509526 373076 509582 373110
rect 509616 373076 509732 373110
rect 508444 373045 509732 373076
rect 508444 373034 508543 373045
rect 508444 373000 508464 373034
rect 508498 373014 508543 373034
rect 508444 372980 508479 373000
rect 508513 372980 508543 373014
rect 509633 373014 509732 373045
rect 508444 372944 508543 372980
rect 508444 372910 508464 372944
rect 508498 372924 508543 372944
rect 508444 372890 508479 372910
rect 508513 372890 508543 372924
rect 508444 372854 508543 372890
rect 508444 372820 508464 372854
rect 508498 372834 508543 372854
rect 508444 372800 508479 372820
rect 508513 372800 508543 372834
rect 508444 372764 508543 372800
rect 508444 372730 508464 372764
rect 508498 372744 508543 372764
rect 508444 372710 508479 372730
rect 508513 372710 508543 372744
rect 508444 372674 508543 372710
rect 508444 372640 508464 372674
rect 508498 372654 508543 372674
rect 508444 372620 508479 372640
rect 508513 372620 508543 372654
rect 508444 372584 508543 372620
rect 508444 372550 508464 372584
rect 508498 372564 508543 372584
rect 508444 372530 508479 372550
rect 508513 372530 508543 372564
rect 508444 372494 508543 372530
rect 508444 372460 508464 372494
rect 508498 372474 508543 372494
rect 508444 372440 508479 372460
rect 508513 372440 508543 372474
rect 508444 372404 508543 372440
rect 508444 372370 508464 372404
rect 508498 372384 508543 372404
rect 508444 372350 508479 372370
rect 508513 372350 508543 372384
rect 508444 372314 508543 372350
rect 508444 372280 508464 372314
rect 508498 372294 508543 372314
rect 508444 372260 508479 372280
rect 508513 372260 508543 372294
rect 508444 372224 508543 372260
rect 508444 372190 508464 372224
rect 508498 372204 508543 372224
rect 508444 372170 508479 372190
rect 508513 372170 508543 372204
rect 508444 372134 508543 372170
rect 508444 372100 508464 372134
rect 508498 372114 508543 372134
rect 508444 372080 508479 372100
rect 508513 372080 508543 372114
rect 508444 372044 508543 372080
rect 508444 372010 508464 372044
rect 508498 372024 508543 372044
rect 508444 371990 508479 372010
rect 508513 371990 508543 372024
rect 508607 372962 509569 372981
rect 508607 372960 508683 372962
rect 508607 372926 508624 372960
rect 508658 372928 508683 372960
rect 508717 372928 508773 372962
rect 508807 372928 508863 372962
rect 508897 372928 508953 372962
rect 508987 372928 509043 372962
rect 509077 372928 509133 372962
rect 509167 372928 509223 372962
rect 509257 372928 509313 372962
rect 509347 372928 509403 372962
rect 509437 372928 509569 372962
rect 508658 372926 509569 372928
rect 508607 372909 509569 372926
rect 508607 372870 508679 372909
rect 508607 372836 508624 372870
rect 508658 372850 508679 372870
rect 508607 372816 508626 372836
rect 508660 372816 508679 372850
rect 509497 372884 509569 372909
rect 509497 372850 509516 372884
rect 509550 372850 509569 372884
rect 508607 372780 508679 372816
rect 508607 372746 508624 372780
rect 508658 372760 508679 372780
rect 508607 372726 508626 372746
rect 508660 372726 508679 372760
rect 508607 372690 508679 372726
rect 508607 372656 508624 372690
rect 508658 372670 508679 372690
rect 508607 372636 508626 372656
rect 508660 372636 508679 372670
rect 508607 372600 508679 372636
rect 508607 372566 508624 372600
rect 508658 372580 508679 372600
rect 508607 372546 508626 372566
rect 508660 372546 508679 372580
rect 508607 372510 508679 372546
rect 508607 372476 508624 372510
rect 508658 372490 508679 372510
rect 508607 372456 508626 372476
rect 508660 372456 508679 372490
rect 508607 372420 508679 372456
rect 508607 372386 508624 372420
rect 508658 372400 508679 372420
rect 508607 372366 508626 372386
rect 508660 372366 508679 372400
rect 508607 372330 508679 372366
rect 508607 372296 508624 372330
rect 508658 372310 508679 372330
rect 508607 372276 508626 372296
rect 508660 372276 508679 372310
rect 508607 372240 508679 372276
rect 508607 372206 508624 372240
rect 508658 372220 508679 372240
rect 508607 372186 508626 372206
rect 508660 372186 508679 372220
rect 508607 372150 508679 372186
rect 508741 372786 509435 372847
rect 508741 372752 508800 372786
rect 508834 372774 508890 372786
rect 508862 372752 508890 372774
rect 508924 372774 508980 372786
rect 508924 372752 508928 372774
rect 508741 372740 508828 372752
rect 508862 372740 508928 372752
rect 508962 372752 508980 372774
rect 509014 372774 509070 372786
rect 509014 372752 509028 372774
rect 508962 372740 509028 372752
rect 509062 372752 509070 372774
rect 509104 372774 509160 372786
rect 509194 372774 509250 372786
rect 509284 372774 509340 372786
rect 509104 372752 509128 372774
rect 509194 372752 509228 372774
rect 509284 372752 509328 372774
rect 509374 372752 509435 372786
rect 509062 372740 509128 372752
rect 509162 372740 509228 372752
rect 509262 372740 509328 372752
rect 509362 372740 509435 372752
rect 508741 372696 509435 372740
rect 508741 372662 508800 372696
rect 508834 372674 508890 372696
rect 508862 372662 508890 372674
rect 508924 372674 508980 372696
rect 508924 372662 508928 372674
rect 508741 372640 508828 372662
rect 508862 372640 508928 372662
rect 508962 372662 508980 372674
rect 509014 372674 509070 372696
rect 509014 372662 509028 372674
rect 508962 372640 509028 372662
rect 509062 372662 509070 372674
rect 509104 372674 509160 372696
rect 509194 372674 509250 372696
rect 509284 372674 509340 372696
rect 509104 372662 509128 372674
rect 509194 372662 509228 372674
rect 509284 372662 509328 372674
rect 509374 372662 509435 372696
rect 509062 372640 509128 372662
rect 509162 372640 509228 372662
rect 509262 372640 509328 372662
rect 509362 372640 509435 372662
rect 508741 372606 509435 372640
rect 508741 372572 508800 372606
rect 508834 372574 508890 372606
rect 508862 372572 508890 372574
rect 508924 372574 508980 372606
rect 508924 372572 508928 372574
rect 508741 372540 508828 372572
rect 508862 372540 508928 372572
rect 508962 372572 508980 372574
rect 509014 372574 509070 372606
rect 509014 372572 509028 372574
rect 508962 372540 509028 372572
rect 509062 372572 509070 372574
rect 509104 372574 509160 372606
rect 509194 372574 509250 372606
rect 509284 372574 509340 372606
rect 509104 372572 509128 372574
rect 509194 372572 509228 372574
rect 509284 372572 509328 372574
rect 509374 372572 509435 372606
rect 509062 372540 509128 372572
rect 509162 372540 509228 372572
rect 509262 372540 509328 372572
rect 509362 372540 509435 372572
rect 508741 372516 509435 372540
rect 508741 372482 508800 372516
rect 508834 372482 508890 372516
rect 508924 372482 508980 372516
rect 509014 372482 509070 372516
rect 509104 372482 509160 372516
rect 509194 372482 509250 372516
rect 509284 372482 509340 372516
rect 509374 372482 509435 372516
rect 508741 372474 509435 372482
rect 508741 372440 508828 372474
rect 508862 372440 508928 372474
rect 508962 372440 509028 372474
rect 509062 372440 509128 372474
rect 509162 372440 509228 372474
rect 509262 372440 509328 372474
rect 509362 372440 509435 372474
rect 508741 372426 509435 372440
rect 508741 372392 508800 372426
rect 508834 372392 508890 372426
rect 508924 372392 508980 372426
rect 509014 372392 509070 372426
rect 509104 372392 509160 372426
rect 509194 372392 509250 372426
rect 509284 372392 509340 372426
rect 509374 372392 509435 372426
rect 508741 372374 509435 372392
rect 508741 372340 508828 372374
rect 508862 372340 508928 372374
rect 508962 372340 509028 372374
rect 509062 372340 509128 372374
rect 509162 372340 509228 372374
rect 509262 372340 509328 372374
rect 509362 372340 509435 372374
rect 508741 372336 509435 372340
rect 508741 372302 508800 372336
rect 508834 372302 508890 372336
rect 508924 372302 508980 372336
rect 509014 372302 509070 372336
rect 509104 372302 509160 372336
rect 509194 372302 509250 372336
rect 509284 372302 509340 372336
rect 509374 372302 509435 372336
rect 508741 372274 509435 372302
rect 508741 372246 508828 372274
rect 508862 372246 508928 372274
rect 508741 372212 508800 372246
rect 508862 372240 508890 372246
rect 508834 372212 508890 372240
rect 508924 372240 508928 372246
rect 508962 372246 509028 372274
rect 508962 372240 508980 372246
rect 508924 372212 508980 372240
rect 509014 372240 509028 372246
rect 509062 372246 509128 372274
rect 509162 372246 509228 372274
rect 509262 372246 509328 372274
rect 509362 372246 509435 372274
rect 509062 372240 509070 372246
rect 509014 372212 509070 372240
rect 509104 372240 509128 372246
rect 509194 372240 509228 372246
rect 509284 372240 509328 372246
rect 509104 372212 509160 372240
rect 509194 372212 509250 372240
rect 509284 372212 509340 372240
rect 509374 372212 509435 372246
rect 508741 372153 509435 372212
rect 509497 372794 509569 372850
rect 509497 372760 509516 372794
rect 509550 372760 509569 372794
rect 509497 372704 509569 372760
rect 509497 372670 509516 372704
rect 509550 372670 509569 372704
rect 509497 372614 509569 372670
rect 509497 372580 509516 372614
rect 509550 372580 509569 372614
rect 509497 372524 509569 372580
rect 509497 372490 509516 372524
rect 509550 372490 509569 372524
rect 509497 372434 509569 372490
rect 509497 372400 509516 372434
rect 509550 372400 509569 372434
rect 509497 372344 509569 372400
rect 509497 372310 509516 372344
rect 509550 372310 509569 372344
rect 509497 372254 509569 372310
rect 509497 372220 509516 372254
rect 509550 372220 509569 372254
rect 509497 372164 509569 372220
rect 508607 372116 508624 372150
rect 508658 372130 508679 372150
rect 508607 372096 508626 372116
rect 508660 372096 508679 372130
rect 508607 372091 508679 372096
rect 509497 372130 509516 372164
rect 509550 372130 509569 372164
rect 509497 372091 509569 372130
rect 508607 372072 509569 372091
rect 508607 372060 508702 372072
rect 508607 372026 508624 372060
rect 508658 372038 508702 372060
rect 508736 372038 508792 372072
rect 508826 372038 508882 372072
rect 508916 372038 508972 372072
rect 509006 372038 509062 372072
rect 509096 372038 509152 372072
rect 509186 372038 509242 372072
rect 509276 372038 509332 372072
rect 509366 372038 509422 372072
rect 509456 372038 509569 372072
rect 508658 372026 509569 372038
rect 508607 372019 509569 372026
rect 509633 372980 509666 373014
rect 509700 372980 509732 373014
rect 509633 372924 509732 372980
rect 509633 372890 509666 372924
rect 509700 372890 509732 372924
rect 509633 372834 509732 372890
rect 509633 372800 509666 372834
rect 509700 372800 509732 372834
rect 509633 372744 509732 372800
rect 509633 372710 509666 372744
rect 509700 372710 509732 372744
rect 509633 372654 509732 372710
rect 509633 372620 509666 372654
rect 509700 372620 509732 372654
rect 509633 372564 509732 372620
rect 509633 372530 509666 372564
rect 509700 372530 509732 372564
rect 509633 372474 509732 372530
rect 509633 372440 509666 372474
rect 509700 372440 509732 372474
rect 509633 372384 509732 372440
rect 509633 372350 509666 372384
rect 509700 372350 509732 372384
rect 509633 372294 509732 372350
rect 509633 372260 509666 372294
rect 509700 372260 509732 372294
rect 509633 372204 509732 372260
rect 509633 372170 509666 372204
rect 509700 372170 509732 372204
rect 509633 372114 509732 372170
rect 509633 372080 509666 372114
rect 509700 372080 509732 372114
rect 509633 372024 509732 372080
rect 508444 371955 508543 371990
rect 509633 371990 509666 372024
rect 509700 371990 509732 372024
rect 509633 371955 509732 371990
rect 508444 371954 509732 371955
rect 508444 371920 508464 371954
rect 508498 371923 509732 371954
rect 508498 371920 508502 371923
rect 508444 371889 508502 371920
rect 508536 371889 508592 371923
rect 508626 371889 508682 371923
rect 508716 371889 508772 371923
rect 508806 371889 508862 371923
rect 508896 371889 508952 371923
rect 508986 371889 509042 371923
rect 509076 371889 509132 371923
rect 509166 371889 509222 371923
rect 509256 371889 509312 371923
rect 509346 371889 509402 371923
rect 509436 371889 509492 371923
rect 509526 371889 509582 371923
rect 509616 371889 509732 371923
rect 508444 371784 509732 371889
rect 508444 371750 508464 371784
rect 508498 371770 509732 371784
rect 508498 371750 508502 371770
rect 508444 371736 508502 371750
rect 508536 371736 508592 371770
rect 508626 371736 508682 371770
rect 508716 371736 508772 371770
rect 508806 371736 508862 371770
rect 508896 371736 508952 371770
rect 508986 371736 509042 371770
rect 509076 371736 509132 371770
rect 509166 371736 509222 371770
rect 509256 371736 509312 371770
rect 509346 371736 509402 371770
rect 509436 371736 509492 371770
rect 509526 371736 509582 371770
rect 509616 371736 509732 371770
rect 508444 371705 509732 371736
rect 508444 371694 508543 371705
rect 508444 371660 508464 371694
rect 508498 371674 508543 371694
rect 508444 371640 508479 371660
rect 508513 371640 508543 371674
rect 509633 371674 509732 371705
rect 508444 371604 508543 371640
rect 508444 371570 508464 371604
rect 508498 371584 508543 371604
rect 508444 371550 508479 371570
rect 508513 371550 508543 371584
rect 508444 371514 508543 371550
rect 508444 371480 508464 371514
rect 508498 371494 508543 371514
rect 508444 371460 508479 371480
rect 508513 371460 508543 371494
rect 508444 371424 508543 371460
rect 508444 371390 508464 371424
rect 508498 371404 508543 371424
rect 508444 371370 508479 371390
rect 508513 371370 508543 371404
rect 508444 371334 508543 371370
rect 508444 371300 508464 371334
rect 508498 371314 508543 371334
rect 508444 371280 508479 371300
rect 508513 371280 508543 371314
rect 508444 371244 508543 371280
rect 508444 371210 508464 371244
rect 508498 371224 508543 371244
rect 508444 371190 508479 371210
rect 508513 371190 508543 371224
rect 508444 371154 508543 371190
rect 508444 371120 508464 371154
rect 508498 371134 508543 371154
rect 508444 371100 508479 371120
rect 508513 371100 508543 371134
rect 508444 371064 508543 371100
rect 508444 371030 508464 371064
rect 508498 371044 508543 371064
rect 508444 371010 508479 371030
rect 508513 371010 508543 371044
rect 508444 370974 508543 371010
rect 508444 370940 508464 370974
rect 508498 370954 508543 370974
rect 508444 370920 508479 370940
rect 508513 370920 508543 370954
rect 508444 370884 508543 370920
rect 508444 370850 508464 370884
rect 508498 370864 508543 370884
rect 508444 370830 508479 370850
rect 508513 370830 508543 370864
rect 508444 370794 508543 370830
rect 508444 370760 508464 370794
rect 508498 370774 508543 370794
rect 508444 370740 508479 370760
rect 508513 370740 508543 370774
rect 508444 370704 508543 370740
rect 508444 370670 508464 370704
rect 508498 370684 508543 370704
rect 508444 370650 508479 370670
rect 508513 370650 508543 370684
rect 508607 371622 509569 371641
rect 508607 371620 508683 371622
rect 508607 371586 508624 371620
rect 508658 371588 508683 371620
rect 508717 371588 508773 371622
rect 508807 371588 508863 371622
rect 508897 371588 508953 371622
rect 508987 371588 509043 371622
rect 509077 371588 509133 371622
rect 509167 371588 509223 371622
rect 509257 371588 509313 371622
rect 509347 371588 509403 371622
rect 509437 371588 509569 371622
rect 508658 371586 509569 371588
rect 508607 371569 509569 371586
rect 508607 371530 508679 371569
rect 508607 371496 508624 371530
rect 508658 371510 508679 371530
rect 508607 371476 508626 371496
rect 508660 371476 508679 371510
rect 509497 371544 509569 371569
rect 509497 371510 509516 371544
rect 509550 371510 509569 371544
rect 508607 371440 508679 371476
rect 508607 371406 508624 371440
rect 508658 371420 508679 371440
rect 508607 371386 508626 371406
rect 508660 371386 508679 371420
rect 508607 371350 508679 371386
rect 508607 371316 508624 371350
rect 508658 371330 508679 371350
rect 508607 371296 508626 371316
rect 508660 371296 508679 371330
rect 508607 371260 508679 371296
rect 508607 371226 508624 371260
rect 508658 371240 508679 371260
rect 508607 371206 508626 371226
rect 508660 371206 508679 371240
rect 508607 371170 508679 371206
rect 508607 371136 508624 371170
rect 508658 371150 508679 371170
rect 508607 371116 508626 371136
rect 508660 371116 508679 371150
rect 508607 371080 508679 371116
rect 508607 371046 508624 371080
rect 508658 371060 508679 371080
rect 508607 371026 508626 371046
rect 508660 371026 508679 371060
rect 508607 370990 508679 371026
rect 508607 370956 508624 370990
rect 508658 370970 508679 370990
rect 508607 370936 508626 370956
rect 508660 370936 508679 370970
rect 508607 370900 508679 370936
rect 508607 370866 508624 370900
rect 508658 370880 508679 370900
rect 508607 370846 508626 370866
rect 508660 370846 508679 370880
rect 508607 370810 508679 370846
rect 508741 371446 509435 371507
rect 508741 371412 508800 371446
rect 508834 371434 508890 371446
rect 508862 371412 508890 371434
rect 508924 371434 508980 371446
rect 508924 371412 508928 371434
rect 508741 371400 508828 371412
rect 508862 371400 508928 371412
rect 508962 371412 508980 371434
rect 509014 371434 509070 371446
rect 509014 371412 509028 371434
rect 508962 371400 509028 371412
rect 509062 371412 509070 371434
rect 509104 371434 509160 371446
rect 509194 371434 509250 371446
rect 509284 371434 509340 371446
rect 509104 371412 509128 371434
rect 509194 371412 509228 371434
rect 509284 371412 509328 371434
rect 509374 371412 509435 371446
rect 509062 371400 509128 371412
rect 509162 371400 509228 371412
rect 509262 371400 509328 371412
rect 509362 371400 509435 371412
rect 508741 371356 509435 371400
rect 508741 371322 508800 371356
rect 508834 371334 508890 371356
rect 508862 371322 508890 371334
rect 508924 371334 508980 371356
rect 508924 371322 508928 371334
rect 508741 371300 508828 371322
rect 508862 371300 508928 371322
rect 508962 371322 508980 371334
rect 509014 371334 509070 371356
rect 509014 371322 509028 371334
rect 508962 371300 509028 371322
rect 509062 371322 509070 371334
rect 509104 371334 509160 371356
rect 509194 371334 509250 371356
rect 509284 371334 509340 371356
rect 509104 371322 509128 371334
rect 509194 371322 509228 371334
rect 509284 371322 509328 371334
rect 509374 371322 509435 371356
rect 509062 371300 509128 371322
rect 509162 371300 509228 371322
rect 509262 371300 509328 371322
rect 509362 371300 509435 371322
rect 508741 371266 509435 371300
rect 508741 371232 508800 371266
rect 508834 371234 508890 371266
rect 508862 371232 508890 371234
rect 508924 371234 508980 371266
rect 508924 371232 508928 371234
rect 508741 371200 508828 371232
rect 508862 371200 508928 371232
rect 508962 371232 508980 371234
rect 509014 371234 509070 371266
rect 509014 371232 509028 371234
rect 508962 371200 509028 371232
rect 509062 371232 509070 371234
rect 509104 371234 509160 371266
rect 509194 371234 509250 371266
rect 509284 371234 509340 371266
rect 509104 371232 509128 371234
rect 509194 371232 509228 371234
rect 509284 371232 509328 371234
rect 509374 371232 509435 371266
rect 509062 371200 509128 371232
rect 509162 371200 509228 371232
rect 509262 371200 509328 371232
rect 509362 371200 509435 371232
rect 508741 371176 509435 371200
rect 508741 371142 508800 371176
rect 508834 371142 508890 371176
rect 508924 371142 508980 371176
rect 509014 371142 509070 371176
rect 509104 371142 509160 371176
rect 509194 371142 509250 371176
rect 509284 371142 509340 371176
rect 509374 371142 509435 371176
rect 508741 371134 509435 371142
rect 508741 371100 508828 371134
rect 508862 371100 508928 371134
rect 508962 371100 509028 371134
rect 509062 371100 509128 371134
rect 509162 371100 509228 371134
rect 509262 371100 509328 371134
rect 509362 371100 509435 371134
rect 508741 371086 509435 371100
rect 508741 371052 508800 371086
rect 508834 371052 508890 371086
rect 508924 371052 508980 371086
rect 509014 371052 509070 371086
rect 509104 371052 509160 371086
rect 509194 371052 509250 371086
rect 509284 371052 509340 371086
rect 509374 371052 509435 371086
rect 508741 371034 509435 371052
rect 508741 371000 508828 371034
rect 508862 371000 508928 371034
rect 508962 371000 509028 371034
rect 509062 371000 509128 371034
rect 509162 371000 509228 371034
rect 509262 371000 509328 371034
rect 509362 371000 509435 371034
rect 508741 370996 509435 371000
rect 508741 370962 508800 370996
rect 508834 370962 508890 370996
rect 508924 370962 508980 370996
rect 509014 370962 509070 370996
rect 509104 370962 509160 370996
rect 509194 370962 509250 370996
rect 509284 370962 509340 370996
rect 509374 370962 509435 370996
rect 508741 370934 509435 370962
rect 508741 370906 508828 370934
rect 508862 370906 508928 370934
rect 508741 370872 508800 370906
rect 508862 370900 508890 370906
rect 508834 370872 508890 370900
rect 508924 370900 508928 370906
rect 508962 370906 509028 370934
rect 508962 370900 508980 370906
rect 508924 370872 508980 370900
rect 509014 370900 509028 370906
rect 509062 370906 509128 370934
rect 509162 370906 509228 370934
rect 509262 370906 509328 370934
rect 509362 370906 509435 370934
rect 509062 370900 509070 370906
rect 509014 370872 509070 370900
rect 509104 370900 509128 370906
rect 509194 370900 509228 370906
rect 509284 370900 509328 370906
rect 509104 370872 509160 370900
rect 509194 370872 509250 370900
rect 509284 370872 509340 370900
rect 509374 370872 509435 370906
rect 508741 370813 509435 370872
rect 509497 371454 509569 371510
rect 509497 371420 509516 371454
rect 509550 371420 509569 371454
rect 509497 371364 509569 371420
rect 509497 371330 509516 371364
rect 509550 371330 509569 371364
rect 509497 371274 509569 371330
rect 509497 371240 509516 371274
rect 509550 371240 509569 371274
rect 509497 371184 509569 371240
rect 509497 371150 509516 371184
rect 509550 371150 509569 371184
rect 509497 371094 509569 371150
rect 509497 371060 509516 371094
rect 509550 371060 509569 371094
rect 509497 371004 509569 371060
rect 509497 370970 509516 371004
rect 509550 370970 509569 371004
rect 509497 370914 509569 370970
rect 509497 370880 509516 370914
rect 509550 370880 509569 370914
rect 509497 370824 509569 370880
rect 508607 370776 508624 370810
rect 508658 370790 508679 370810
rect 508607 370756 508626 370776
rect 508660 370756 508679 370790
rect 508607 370751 508679 370756
rect 509497 370790 509516 370824
rect 509550 370790 509569 370824
rect 509497 370751 509569 370790
rect 508607 370732 509569 370751
rect 508607 370720 508702 370732
rect 508607 370686 508624 370720
rect 508658 370698 508702 370720
rect 508736 370698 508792 370732
rect 508826 370698 508882 370732
rect 508916 370698 508972 370732
rect 509006 370698 509062 370732
rect 509096 370698 509152 370732
rect 509186 370698 509242 370732
rect 509276 370698 509332 370732
rect 509366 370698 509422 370732
rect 509456 370698 509569 370732
rect 508658 370686 509569 370698
rect 508607 370679 509569 370686
rect 509633 371640 509666 371674
rect 509700 371640 509732 371674
rect 509633 371584 509732 371640
rect 509633 371550 509666 371584
rect 509700 371550 509732 371584
rect 509633 371494 509732 371550
rect 509633 371460 509666 371494
rect 509700 371460 509732 371494
rect 509633 371404 509732 371460
rect 509633 371370 509666 371404
rect 509700 371370 509732 371404
rect 509633 371314 509732 371370
rect 509633 371280 509666 371314
rect 509700 371280 509732 371314
rect 509633 371224 509732 371280
rect 509633 371190 509666 371224
rect 509700 371190 509732 371224
rect 509633 371134 509732 371190
rect 509633 371100 509666 371134
rect 509700 371100 509732 371134
rect 509633 371044 509732 371100
rect 509633 371010 509666 371044
rect 509700 371010 509732 371044
rect 509633 370954 509732 371010
rect 509633 370920 509666 370954
rect 509700 370920 509732 370954
rect 509633 370864 509732 370920
rect 509633 370830 509666 370864
rect 509700 370830 509732 370864
rect 509633 370774 509732 370830
rect 509633 370740 509666 370774
rect 509700 370740 509732 370774
rect 509633 370684 509732 370740
rect 508444 370615 508543 370650
rect 509633 370650 509666 370684
rect 509700 370650 509732 370684
rect 509633 370615 509732 370650
rect 508444 370614 509732 370615
rect 508444 370580 508464 370614
rect 508498 370583 509732 370614
rect 508498 370580 508502 370583
rect 508444 370549 508502 370580
rect 508536 370549 508592 370583
rect 508626 370549 508682 370583
rect 508716 370549 508772 370583
rect 508806 370549 508862 370583
rect 508896 370549 508952 370583
rect 508986 370549 509042 370583
rect 509076 370549 509132 370583
rect 509166 370549 509222 370583
rect 509256 370549 509312 370583
rect 509346 370549 509402 370583
rect 509436 370549 509492 370583
rect 509526 370549 509582 370583
rect 509616 370549 509732 370583
rect 508444 370444 509732 370549
rect 508444 370410 508464 370444
rect 508498 370430 509732 370444
rect 508498 370410 508502 370430
rect 508444 370396 508502 370410
rect 508536 370396 508592 370430
rect 508626 370396 508682 370430
rect 508716 370396 508772 370430
rect 508806 370396 508862 370430
rect 508896 370396 508952 370430
rect 508986 370396 509042 370430
rect 509076 370396 509132 370430
rect 509166 370396 509222 370430
rect 509256 370396 509312 370430
rect 509346 370396 509402 370430
rect 509436 370396 509492 370430
rect 509526 370396 509582 370430
rect 509616 370396 509732 370430
rect 508444 370365 509732 370396
rect 508444 370354 508543 370365
rect 508444 370320 508464 370354
rect 508498 370334 508543 370354
rect 508444 370300 508479 370320
rect 508513 370300 508543 370334
rect 509633 370334 509732 370365
rect 508444 370264 508543 370300
rect 508444 370230 508464 370264
rect 508498 370244 508543 370264
rect 508444 370210 508479 370230
rect 508513 370210 508543 370244
rect 508444 370174 508543 370210
rect 508444 370140 508464 370174
rect 508498 370154 508543 370174
rect 508444 370120 508479 370140
rect 508513 370120 508543 370154
rect 508444 370084 508543 370120
rect 508444 370050 508464 370084
rect 508498 370064 508543 370084
rect 508444 370030 508479 370050
rect 508513 370030 508543 370064
rect 508444 369994 508543 370030
rect 508444 369960 508464 369994
rect 508498 369974 508543 369994
rect 508444 369940 508479 369960
rect 508513 369940 508543 369974
rect 508444 369904 508543 369940
rect 508444 369870 508464 369904
rect 508498 369884 508543 369904
rect 508444 369850 508479 369870
rect 508513 369850 508543 369884
rect 508444 369814 508543 369850
rect 508444 369780 508464 369814
rect 508498 369794 508543 369814
rect 508444 369760 508479 369780
rect 508513 369760 508543 369794
rect 508444 369724 508543 369760
rect 508444 369690 508464 369724
rect 508498 369704 508543 369724
rect 508444 369670 508479 369690
rect 508513 369670 508543 369704
rect 508444 369634 508543 369670
rect 508444 369600 508464 369634
rect 508498 369614 508543 369634
rect 508444 369580 508479 369600
rect 508513 369580 508543 369614
rect 508444 369544 508543 369580
rect 508444 369510 508464 369544
rect 508498 369524 508543 369544
rect 508444 369490 508479 369510
rect 508513 369490 508543 369524
rect 508444 369454 508543 369490
rect 508444 369420 508464 369454
rect 508498 369434 508543 369454
rect 508444 369400 508479 369420
rect 508513 369400 508543 369434
rect 508444 369364 508543 369400
rect 508444 369330 508464 369364
rect 508498 369344 508543 369364
rect 508444 369310 508479 369330
rect 508513 369310 508543 369344
rect 508607 370282 509569 370301
rect 508607 370280 508683 370282
rect 508607 370246 508624 370280
rect 508658 370248 508683 370280
rect 508717 370248 508773 370282
rect 508807 370248 508863 370282
rect 508897 370248 508953 370282
rect 508987 370248 509043 370282
rect 509077 370248 509133 370282
rect 509167 370248 509223 370282
rect 509257 370248 509313 370282
rect 509347 370248 509403 370282
rect 509437 370248 509569 370282
rect 508658 370246 509569 370248
rect 508607 370229 509569 370246
rect 508607 370190 508679 370229
rect 508607 370156 508624 370190
rect 508658 370170 508679 370190
rect 508607 370136 508626 370156
rect 508660 370136 508679 370170
rect 509497 370204 509569 370229
rect 509497 370170 509516 370204
rect 509550 370170 509569 370204
rect 508607 370100 508679 370136
rect 508607 370066 508624 370100
rect 508658 370080 508679 370100
rect 508607 370046 508626 370066
rect 508660 370046 508679 370080
rect 508607 370010 508679 370046
rect 508607 369976 508624 370010
rect 508658 369990 508679 370010
rect 508607 369956 508626 369976
rect 508660 369956 508679 369990
rect 508607 369920 508679 369956
rect 508607 369886 508624 369920
rect 508658 369900 508679 369920
rect 508607 369866 508626 369886
rect 508660 369866 508679 369900
rect 508607 369830 508679 369866
rect 508607 369796 508624 369830
rect 508658 369810 508679 369830
rect 508607 369776 508626 369796
rect 508660 369776 508679 369810
rect 508607 369740 508679 369776
rect 508607 369706 508624 369740
rect 508658 369720 508679 369740
rect 508607 369686 508626 369706
rect 508660 369686 508679 369720
rect 508607 369650 508679 369686
rect 508607 369616 508624 369650
rect 508658 369630 508679 369650
rect 508607 369596 508626 369616
rect 508660 369596 508679 369630
rect 508607 369560 508679 369596
rect 508607 369526 508624 369560
rect 508658 369540 508679 369560
rect 508607 369506 508626 369526
rect 508660 369506 508679 369540
rect 508607 369470 508679 369506
rect 508741 370106 509435 370167
rect 508741 370072 508800 370106
rect 508834 370094 508890 370106
rect 508862 370072 508890 370094
rect 508924 370094 508980 370106
rect 508924 370072 508928 370094
rect 508741 370060 508828 370072
rect 508862 370060 508928 370072
rect 508962 370072 508980 370094
rect 509014 370094 509070 370106
rect 509014 370072 509028 370094
rect 508962 370060 509028 370072
rect 509062 370072 509070 370094
rect 509104 370094 509160 370106
rect 509194 370094 509250 370106
rect 509284 370094 509340 370106
rect 509104 370072 509128 370094
rect 509194 370072 509228 370094
rect 509284 370072 509328 370094
rect 509374 370072 509435 370106
rect 509062 370060 509128 370072
rect 509162 370060 509228 370072
rect 509262 370060 509328 370072
rect 509362 370060 509435 370072
rect 508741 370016 509435 370060
rect 508741 369982 508800 370016
rect 508834 369994 508890 370016
rect 508862 369982 508890 369994
rect 508924 369994 508980 370016
rect 508924 369982 508928 369994
rect 508741 369960 508828 369982
rect 508862 369960 508928 369982
rect 508962 369982 508980 369994
rect 509014 369994 509070 370016
rect 509014 369982 509028 369994
rect 508962 369960 509028 369982
rect 509062 369982 509070 369994
rect 509104 369994 509160 370016
rect 509194 369994 509250 370016
rect 509284 369994 509340 370016
rect 509104 369982 509128 369994
rect 509194 369982 509228 369994
rect 509284 369982 509328 369994
rect 509374 369982 509435 370016
rect 509062 369960 509128 369982
rect 509162 369960 509228 369982
rect 509262 369960 509328 369982
rect 509362 369960 509435 369982
rect 508741 369926 509435 369960
rect 508741 369892 508800 369926
rect 508834 369894 508890 369926
rect 508862 369892 508890 369894
rect 508924 369894 508980 369926
rect 508924 369892 508928 369894
rect 508741 369860 508828 369892
rect 508862 369860 508928 369892
rect 508962 369892 508980 369894
rect 509014 369894 509070 369926
rect 509014 369892 509028 369894
rect 508962 369860 509028 369892
rect 509062 369892 509070 369894
rect 509104 369894 509160 369926
rect 509194 369894 509250 369926
rect 509284 369894 509340 369926
rect 509104 369892 509128 369894
rect 509194 369892 509228 369894
rect 509284 369892 509328 369894
rect 509374 369892 509435 369926
rect 509062 369860 509128 369892
rect 509162 369860 509228 369892
rect 509262 369860 509328 369892
rect 509362 369860 509435 369892
rect 508741 369836 509435 369860
rect 508741 369802 508800 369836
rect 508834 369802 508890 369836
rect 508924 369802 508980 369836
rect 509014 369802 509070 369836
rect 509104 369802 509160 369836
rect 509194 369802 509250 369836
rect 509284 369802 509340 369836
rect 509374 369802 509435 369836
rect 508741 369794 509435 369802
rect 508741 369760 508828 369794
rect 508862 369760 508928 369794
rect 508962 369760 509028 369794
rect 509062 369760 509128 369794
rect 509162 369760 509228 369794
rect 509262 369760 509328 369794
rect 509362 369760 509435 369794
rect 508741 369746 509435 369760
rect 508741 369712 508800 369746
rect 508834 369712 508890 369746
rect 508924 369712 508980 369746
rect 509014 369712 509070 369746
rect 509104 369712 509160 369746
rect 509194 369712 509250 369746
rect 509284 369712 509340 369746
rect 509374 369712 509435 369746
rect 508741 369694 509435 369712
rect 508741 369660 508828 369694
rect 508862 369660 508928 369694
rect 508962 369660 509028 369694
rect 509062 369660 509128 369694
rect 509162 369660 509228 369694
rect 509262 369660 509328 369694
rect 509362 369660 509435 369694
rect 508741 369656 509435 369660
rect 508741 369622 508800 369656
rect 508834 369622 508890 369656
rect 508924 369622 508980 369656
rect 509014 369622 509070 369656
rect 509104 369622 509160 369656
rect 509194 369622 509250 369656
rect 509284 369622 509340 369656
rect 509374 369622 509435 369656
rect 508741 369594 509435 369622
rect 508741 369566 508828 369594
rect 508862 369566 508928 369594
rect 508741 369532 508800 369566
rect 508862 369560 508890 369566
rect 508834 369532 508890 369560
rect 508924 369560 508928 369566
rect 508962 369566 509028 369594
rect 508962 369560 508980 369566
rect 508924 369532 508980 369560
rect 509014 369560 509028 369566
rect 509062 369566 509128 369594
rect 509162 369566 509228 369594
rect 509262 369566 509328 369594
rect 509362 369566 509435 369594
rect 509062 369560 509070 369566
rect 509014 369532 509070 369560
rect 509104 369560 509128 369566
rect 509194 369560 509228 369566
rect 509284 369560 509328 369566
rect 509104 369532 509160 369560
rect 509194 369532 509250 369560
rect 509284 369532 509340 369560
rect 509374 369532 509435 369566
rect 508741 369473 509435 369532
rect 509497 370114 509569 370170
rect 509497 370080 509516 370114
rect 509550 370080 509569 370114
rect 509497 370024 509569 370080
rect 509497 369990 509516 370024
rect 509550 369990 509569 370024
rect 509497 369934 509569 369990
rect 509497 369900 509516 369934
rect 509550 369900 509569 369934
rect 509497 369844 509569 369900
rect 509497 369810 509516 369844
rect 509550 369810 509569 369844
rect 509497 369754 509569 369810
rect 509497 369720 509516 369754
rect 509550 369720 509569 369754
rect 509497 369664 509569 369720
rect 509497 369630 509516 369664
rect 509550 369630 509569 369664
rect 509497 369574 509569 369630
rect 509497 369540 509516 369574
rect 509550 369540 509569 369574
rect 509497 369484 509569 369540
rect 508607 369436 508624 369470
rect 508658 369450 508679 369470
rect 508607 369416 508626 369436
rect 508660 369416 508679 369450
rect 508607 369411 508679 369416
rect 509497 369450 509516 369484
rect 509550 369450 509569 369484
rect 509497 369411 509569 369450
rect 508607 369392 509569 369411
rect 508607 369380 508702 369392
rect 508607 369346 508624 369380
rect 508658 369358 508702 369380
rect 508736 369358 508792 369392
rect 508826 369358 508882 369392
rect 508916 369358 508972 369392
rect 509006 369358 509062 369392
rect 509096 369358 509152 369392
rect 509186 369358 509242 369392
rect 509276 369358 509332 369392
rect 509366 369358 509422 369392
rect 509456 369358 509569 369392
rect 508658 369346 509569 369358
rect 508607 369339 509569 369346
rect 509633 370300 509666 370334
rect 509700 370300 509732 370334
rect 509633 370244 509732 370300
rect 509633 370210 509666 370244
rect 509700 370210 509732 370244
rect 509633 370154 509732 370210
rect 509633 370120 509666 370154
rect 509700 370120 509732 370154
rect 509633 370064 509732 370120
rect 509633 370030 509666 370064
rect 509700 370030 509732 370064
rect 509633 369974 509732 370030
rect 509633 369940 509666 369974
rect 509700 369940 509732 369974
rect 509633 369884 509732 369940
rect 509633 369850 509666 369884
rect 509700 369850 509732 369884
rect 509633 369794 509732 369850
rect 509633 369760 509666 369794
rect 509700 369760 509732 369794
rect 509633 369704 509732 369760
rect 509633 369670 509666 369704
rect 509700 369670 509732 369704
rect 509633 369614 509732 369670
rect 509633 369580 509666 369614
rect 509700 369580 509732 369614
rect 509633 369524 509732 369580
rect 509633 369490 509666 369524
rect 509700 369490 509732 369524
rect 509633 369434 509732 369490
rect 509633 369400 509666 369434
rect 509700 369400 509732 369434
rect 509633 369344 509732 369400
rect 508444 369275 508543 369310
rect 509633 369310 509666 369344
rect 509700 369310 509732 369344
rect 509633 369275 509732 369310
rect 508444 369274 509732 369275
rect 508444 369240 508464 369274
rect 508498 369243 509732 369274
rect 508498 369240 508502 369243
rect 508444 369209 508502 369240
rect 508536 369209 508592 369243
rect 508626 369209 508682 369243
rect 508716 369209 508772 369243
rect 508806 369209 508862 369243
rect 508896 369209 508952 369243
rect 508986 369209 509042 369243
rect 509076 369209 509132 369243
rect 509166 369209 509222 369243
rect 509256 369209 509312 369243
rect 509346 369209 509402 369243
rect 509436 369209 509492 369243
rect 509526 369209 509582 369243
rect 509616 369209 509732 369243
rect 508444 369104 509732 369209
rect 508444 369070 508464 369104
rect 508498 369090 509732 369104
rect 508498 369070 508502 369090
rect 508444 369056 508502 369070
rect 508536 369056 508592 369090
rect 508626 369056 508682 369090
rect 508716 369056 508772 369090
rect 508806 369056 508862 369090
rect 508896 369056 508952 369090
rect 508986 369056 509042 369090
rect 509076 369056 509132 369090
rect 509166 369056 509222 369090
rect 509256 369056 509312 369090
rect 509346 369056 509402 369090
rect 509436 369056 509492 369090
rect 509526 369056 509582 369090
rect 509616 369056 509732 369090
rect 508444 369025 509732 369056
rect 508444 369014 508543 369025
rect 508444 368980 508464 369014
rect 508498 368994 508543 369014
rect 508444 368960 508479 368980
rect 508513 368960 508543 368994
rect 509633 368994 509732 369025
rect 508444 368924 508543 368960
rect 508444 368890 508464 368924
rect 508498 368904 508543 368924
rect 508444 368870 508479 368890
rect 508513 368870 508543 368904
rect 508444 368834 508543 368870
rect 508444 368800 508464 368834
rect 508498 368814 508543 368834
rect 508444 368780 508479 368800
rect 508513 368780 508543 368814
rect 508444 368744 508543 368780
rect 508444 368710 508464 368744
rect 508498 368724 508543 368744
rect 508444 368690 508479 368710
rect 508513 368690 508543 368724
rect 508444 368654 508543 368690
rect 508444 368620 508464 368654
rect 508498 368634 508543 368654
rect 508444 368600 508479 368620
rect 508513 368600 508543 368634
rect 508444 368564 508543 368600
rect 508444 368530 508464 368564
rect 508498 368544 508543 368564
rect 508444 368510 508479 368530
rect 508513 368510 508543 368544
rect 508444 368474 508543 368510
rect 508444 368440 508464 368474
rect 508498 368454 508543 368474
rect 508444 368420 508479 368440
rect 508513 368420 508543 368454
rect 508444 368384 508543 368420
rect 508444 368350 508464 368384
rect 508498 368364 508543 368384
rect 508444 368330 508479 368350
rect 508513 368330 508543 368364
rect 508444 368294 508543 368330
rect 508444 368260 508464 368294
rect 508498 368274 508543 368294
rect 508444 368240 508479 368260
rect 508513 368240 508543 368274
rect 508444 368204 508543 368240
rect 508444 368170 508464 368204
rect 508498 368184 508543 368204
rect 508444 368150 508479 368170
rect 508513 368150 508543 368184
rect 508444 368114 508543 368150
rect 508444 368080 508464 368114
rect 508498 368094 508543 368114
rect 508444 368060 508479 368080
rect 508513 368060 508543 368094
rect 508444 368024 508543 368060
rect 508444 367990 508464 368024
rect 508498 368004 508543 368024
rect 508444 367970 508479 367990
rect 508513 367970 508543 368004
rect 508607 368942 509569 368961
rect 508607 368940 508683 368942
rect 508607 368906 508624 368940
rect 508658 368908 508683 368940
rect 508717 368908 508773 368942
rect 508807 368908 508863 368942
rect 508897 368908 508953 368942
rect 508987 368908 509043 368942
rect 509077 368908 509133 368942
rect 509167 368908 509223 368942
rect 509257 368908 509313 368942
rect 509347 368908 509403 368942
rect 509437 368908 509569 368942
rect 508658 368906 509569 368908
rect 508607 368889 509569 368906
rect 508607 368850 508679 368889
rect 508607 368816 508624 368850
rect 508658 368830 508679 368850
rect 508607 368796 508626 368816
rect 508660 368796 508679 368830
rect 509497 368864 509569 368889
rect 509497 368830 509516 368864
rect 509550 368830 509569 368864
rect 508607 368760 508679 368796
rect 508607 368726 508624 368760
rect 508658 368740 508679 368760
rect 508607 368706 508626 368726
rect 508660 368706 508679 368740
rect 508607 368670 508679 368706
rect 508607 368636 508624 368670
rect 508658 368650 508679 368670
rect 508607 368616 508626 368636
rect 508660 368616 508679 368650
rect 508607 368580 508679 368616
rect 508607 368546 508624 368580
rect 508658 368560 508679 368580
rect 508607 368526 508626 368546
rect 508660 368526 508679 368560
rect 508607 368490 508679 368526
rect 508607 368456 508624 368490
rect 508658 368470 508679 368490
rect 508607 368436 508626 368456
rect 508660 368436 508679 368470
rect 508607 368400 508679 368436
rect 508607 368366 508624 368400
rect 508658 368380 508679 368400
rect 508607 368346 508626 368366
rect 508660 368346 508679 368380
rect 508607 368310 508679 368346
rect 508607 368276 508624 368310
rect 508658 368290 508679 368310
rect 508607 368256 508626 368276
rect 508660 368256 508679 368290
rect 508607 368220 508679 368256
rect 508607 368186 508624 368220
rect 508658 368200 508679 368220
rect 508607 368166 508626 368186
rect 508660 368166 508679 368200
rect 508607 368130 508679 368166
rect 508741 368766 509435 368827
rect 508741 368732 508800 368766
rect 508834 368754 508890 368766
rect 508862 368732 508890 368754
rect 508924 368754 508980 368766
rect 508924 368732 508928 368754
rect 508741 368720 508828 368732
rect 508862 368720 508928 368732
rect 508962 368732 508980 368754
rect 509014 368754 509070 368766
rect 509014 368732 509028 368754
rect 508962 368720 509028 368732
rect 509062 368732 509070 368754
rect 509104 368754 509160 368766
rect 509194 368754 509250 368766
rect 509284 368754 509340 368766
rect 509104 368732 509128 368754
rect 509194 368732 509228 368754
rect 509284 368732 509328 368754
rect 509374 368732 509435 368766
rect 509062 368720 509128 368732
rect 509162 368720 509228 368732
rect 509262 368720 509328 368732
rect 509362 368720 509435 368732
rect 508741 368676 509435 368720
rect 508741 368642 508800 368676
rect 508834 368654 508890 368676
rect 508862 368642 508890 368654
rect 508924 368654 508980 368676
rect 508924 368642 508928 368654
rect 508741 368620 508828 368642
rect 508862 368620 508928 368642
rect 508962 368642 508980 368654
rect 509014 368654 509070 368676
rect 509014 368642 509028 368654
rect 508962 368620 509028 368642
rect 509062 368642 509070 368654
rect 509104 368654 509160 368676
rect 509194 368654 509250 368676
rect 509284 368654 509340 368676
rect 509104 368642 509128 368654
rect 509194 368642 509228 368654
rect 509284 368642 509328 368654
rect 509374 368642 509435 368676
rect 509062 368620 509128 368642
rect 509162 368620 509228 368642
rect 509262 368620 509328 368642
rect 509362 368620 509435 368642
rect 508741 368586 509435 368620
rect 508741 368552 508800 368586
rect 508834 368554 508890 368586
rect 508862 368552 508890 368554
rect 508924 368554 508980 368586
rect 508924 368552 508928 368554
rect 508741 368520 508828 368552
rect 508862 368520 508928 368552
rect 508962 368552 508980 368554
rect 509014 368554 509070 368586
rect 509014 368552 509028 368554
rect 508962 368520 509028 368552
rect 509062 368552 509070 368554
rect 509104 368554 509160 368586
rect 509194 368554 509250 368586
rect 509284 368554 509340 368586
rect 509104 368552 509128 368554
rect 509194 368552 509228 368554
rect 509284 368552 509328 368554
rect 509374 368552 509435 368586
rect 509062 368520 509128 368552
rect 509162 368520 509228 368552
rect 509262 368520 509328 368552
rect 509362 368520 509435 368552
rect 508741 368496 509435 368520
rect 508741 368462 508800 368496
rect 508834 368462 508890 368496
rect 508924 368462 508980 368496
rect 509014 368462 509070 368496
rect 509104 368462 509160 368496
rect 509194 368462 509250 368496
rect 509284 368462 509340 368496
rect 509374 368462 509435 368496
rect 508741 368454 509435 368462
rect 508741 368420 508828 368454
rect 508862 368420 508928 368454
rect 508962 368420 509028 368454
rect 509062 368420 509128 368454
rect 509162 368420 509228 368454
rect 509262 368420 509328 368454
rect 509362 368420 509435 368454
rect 508741 368406 509435 368420
rect 508741 368372 508800 368406
rect 508834 368372 508890 368406
rect 508924 368372 508980 368406
rect 509014 368372 509070 368406
rect 509104 368372 509160 368406
rect 509194 368372 509250 368406
rect 509284 368372 509340 368406
rect 509374 368372 509435 368406
rect 508741 368354 509435 368372
rect 508741 368320 508828 368354
rect 508862 368320 508928 368354
rect 508962 368320 509028 368354
rect 509062 368320 509128 368354
rect 509162 368320 509228 368354
rect 509262 368320 509328 368354
rect 509362 368320 509435 368354
rect 508741 368316 509435 368320
rect 508741 368282 508800 368316
rect 508834 368282 508890 368316
rect 508924 368282 508980 368316
rect 509014 368282 509070 368316
rect 509104 368282 509160 368316
rect 509194 368282 509250 368316
rect 509284 368282 509340 368316
rect 509374 368282 509435 368316
rect 508741 368254 509435 368282
rect 508741 368226 508828 368254
rect 508862 368226 508928 368254
rect 508741 368192 508800 368226
rect 508862 368220 508890 368226
rect 508834 368192 508890 368220
rect 508924 368220 508928 368226
rect 508962 368226 509028 368254
rect 508962 368220 508980 368226
rect 508924 368192 508980 368220
rect 509014 368220 509028 368226
rect 509062 368226 509128 368254
rect 509162 368226 509228 368254
rect 509262 368226 509328 368254
rect 509362 368226 509435 368254
rect 509062 368220 509070 368226
rect 509014 368192 509070 368220
rect 509104 368220 509128 368226
rect 509194 368220 509228 368226
rect 509284 368220 509328 368226
rect 509104 368192 509160 368220
rect 509194 368192 509250 368220
rect 509284 368192 509340 368220
rect 509374 368192 509435 368226
rect 508741 368133 509435 368192
rect 509497 368774 509569 368830
rect 509497 368740 509516 368774
rect 509550 368740 509569 368774
rect 509497 368684 509569 368740
rect 509497 368650 509516 368684
rect 509550 368650 509569 368684
rect 509497 368594 509569 368650
rect 509497 368560 509516 368594
rect 509550 368560 509569 368594
rect 509497 368504 509569 368560
rect 509497 368470 509516 368504
rect 509550 368470 509569 368504
rect 509497 368414 509569 368470
rect 509497 368380 509516 368414
rect 509550 368380 509569 368414
rect 509497 368324 509569 368380
rect 509497 368290 509516 368324
rect 509550 368290 509569 368324
rect 509497 368234 509569 368290
rect 509497 368200 509516 368234
rect 509550 368200 509569 368234
rect 509497 368144 509569 368200
rect 508607 368096 508624 368130
rect 508658 368110 508679 368130
rect 508607 368076 508626 368096
rect 508660 368076 508679 368110
rect 508607 368071 508679 368076
rect 509497 368110 509516 368144
rect 509550 368110 509569 368144
rect 509497 368071 509569 368110
rect 508607 368052 509569 368071
rect 508607 368040 508702 368052
rect 508607 368006 508624 368040
rect 508658 368018 508702 368040
rect 508736 368018 508792 368052
rect 508826 368018 508882 368052
rect 508916 368018 508972 368052
rect 509006 368018 509062 368052
rect 509096 368018 509152 368052
rect 509186 368018 509242 368052
rect 509276 368018 509332 368052
rect 509366 368018 509422 368052
rect 509456 368018 509569 368052
rect 508658 368006 509569 368018
rect 508607 367999 509569 368006
rect 509633 368960 509666 368994
rect 509700 368960 509732 368994
rect 509633 368904 509732 368960
rect 509633 368870 509666 368904
rect 509700 368870 509732 368904
rect 509633 368814 509732 368870
rect 509633 368780 509666 368814
rect 509700 368780 509732 368814
rect 509633 368724 509732 368780
rect 509633 368690 509666 368724
rect 509700 368690 509732 368724
rect 509633 368634 509732 368690
rect 509633 368600 509666 368634
rect 509700 368600 509732 368634
rect 509633 368544 509732 368600
rect 509633 368510 509666 368544
rect 509700 368510 509732 368544
rect 509633 368454 509732 368510
rect 509633 368420 509666 368454
rect 509700 368420 509732 368454
rect 509633 368364 509732 368420
rect 509633 368330 509666 368364
rect 509700 368330 509732 368364
rect 509633 368274 509732 368330
rect 509633 368240 509666 368274
rect 509700 368240 509732 368274
rect 509633 368184 509732 368240
rect 509633 368150 509666 368184
rect 509700 368150 509732 368184
rect 509633 368094 509732 368150
rect 509633 368060 509666 368094
rect 509700 368060 509732 368094
rect 509633 368004 509732 368060
rect 508444 367935 508543 367970
rect 509633 367970 509666 368004
rect 509700 367970 509732 368004
rect 509633 367935 509732 367970
rect 508444 367934 509732 367935
rect 508444 367900 508464 367934
rect 508498 367903 509732 367934
rect 508498 367900 508502 367903
rect 508444 367869 508502 367900
rect 508536 367869 508592 367903
rect 508626 367869 508682 367903
rect 508716 367869 508772 367903
rect 508806 367869 508862 367903
rect 508896 367869 508952 367903
rect 508986 367869 509042 367903
rect 509076 367869 509132 367903
rect 509166 367869 509222 367903
rect 509256 367869 509312 367903
rect 509346 367869 509402 367903
rect 509436 367869 509492 367903
rect 509526 367869 509582 367903
rect 509616 367869 509732 367903
rect 508444 367764 509732 367869
rect 508444 367730 508464 367764
rect 508498 367750 509732 367764
rect 508498 367730 508502 367750
rect 508444 367716 508502 367730
rect 508536 367716 508592 367750
rect 508626 367716 508682 367750
rect 508716 367716 508772 367750
rect 508806 367716 508862 367750
rect 508896 367716 508952 367750
rect 508986 367716 509042 367750
rect 509076 367716 509132 367750
rect 509166 367716 509222 367750
rect 509256 367716 509312 367750
rect 509346 367716 509402 367750
rect 509436 367716 509492 367750
rect 509526 367716 509582 367750
rect 509616 367716 509732 367750
rect 508444 367685 509732 367716
rect 508444 367674 508543 367685
rect 508444 367640 508464 367674
rect 508498 367654 508543 367674
rect 508444 367620 508479 367640
rect 508513 367620 508543 367654
rect 509633 367654 509732 367685
rect 508444 367584 508543 367620
rect 508444 367550 508464 367584
rect 508498 367564 508543 367584
rect 508444 367530 508479 367550
rect 508513 367530 508543 367564
rect 508444 367494 508543 367530
rect 508444 367460 508464 367494
rect 508498 367474 508543 367494
rect 508444 367440 508479 367460
rect 508513 367440 508543 367474
rect 508444 367404 508543 367440
rect 508444 367370 508464 367404
rect 508498 367384 508543 367404
rect 508444 367350 508479 367370
rect 508513 367350 508543 367384
rect 508444 367314 508543 367350
rect 508444 367280 508464 367314
rect 508498 367294 508543 367314
rect 508444 367260 508479 367280
rect 508513 367260 508543 367294
rect 508444 367224 508543 367260
rect 508444 367190 508464 367224
rect 508498 367204 508543 367224
rect 508444 367170 508479 367190
rect 508513 367170 508543 367204
rect 508444 367134 508543 367170
rect 508444 367100 508464 367134
rect 508498 367114 508543 367134
rect 508444 367080 508479 367100
rect 508513 367080 508543 367114
rect 508444 367044 508543 367080
rect 508444 367010 508464 367044
rect 508498 367024 508543 367044
rect 508444 366990 508479 367010
rect 508513 366990 508543 367024
rect 508444 366954 508543 366990
rect 508444 366920 508464 366954
rect 508498 366934 508543 366954
rect 508444 366900 508479 366920
rect 508513 366900 508543 366934
rect 508444 366864 508543 366900
rect 508444 366830 508464 366864
rect 508498 366844 508543 366864
rect 508444 366810 508479 366830
rect 508513 366810 508543 366844
rect 508444 366774 508543 366810
rect 508444 366740 508464 366774
rect 508498 366754 508543 366774
rect 508444 366720 508479 366740
rect 508513 366720 508543 366754
rect 508444 366684 508543 366720
rect 508444 366650 508464 366684
rect 508498 366664 508543 366684
rect 508444 366630 508479 366650
rect 508513 366630 508543 366664
rect 508607 367602 509569 367621
rect 508607 367600 508683 367602
rect 508607 367566 508624 367600
rect 508658 367568 508683 367600
rect 508717 367568 508773 367602
rect 508807 367568 508863 367602
rect 508897 367568 508953 367602
rect 508987 367568 509043 367602
rect 509077 367568 509133 367602
rect 509167 367568 509223 367602
rect 509257 367568 509313 367602
rect 509347 367568 509403 367602
rect 509437 367568 509569 367602
rect 508658 367566 509569 367568
rect 508607 367549 509569 367566
rect 508607 367510 508679 367549
rect 508607 367476 508624 367510
rect 508658 367490 508679 367510
rect 508607 367456 508626 367476
rect 508660 367456 508679 367490
rect 509497 367524 509569 367549
rect 509497 367490 509516 367524
rect 509550 367490 509569 367524
rect 508607 367420 508679 367456
rect 508607 367386 508624 367420
rect 508658 367400 508679 367420
rect 508607 367366 508626 367386
rect 508660 367366 508679 367400
rect 508607 367330 508679 367366
rect 508607 367296 508624 367330
rect 508658 367310 508679 367330
rect 508607 367276 508626 367296
rect 508660 367276 508679 367310
rect 508607 367240 508679 367276
rect 508607 367206 508624 367240
rect 508658 367220 508679 367240
rect 508607 367186 508626 367206
rect 508660 367186 508679 367220
rect 508607 367150 508679 367186
rect 508607 367116 508624 367150
rect 508658 367130 508679 367150
rect 508607 367096 508626 367116
rect 508660 367096 508679 367130
rect 508607 367060 508679 367096
rect 508607 367026 508624 367060
rect 508658 367040 508679 367060
rect 508607 367006 508626 367026
rect 508660 367006 508679 367040
rect 508607 366970 508679 367006
rect 508607 366936 508624 366970
rect 508658 366950 508679 366970
rect 508607 366916 508626 366936
rect 508660 366916 508679 366950
rect 508607 366880 508679 366916
rect 508607 366846 508624 366880
rect 508658 366860 508679 366880
rect 508607 366826 508626 366846
rect 508660 366826 508679 366860
rect 508607 366790 508679 366826
rect 508741 367426 509435 367487
rect 508741 367392 508800 367426
rect 508834 367414 508890 367426
rect 508862 367392 508890 367414
rect 508924 367414 508980 367426
rect 508924 367392 508928 367414
rect 508741 367380 508828 367392
rect 508862 367380 508928 367392
rect 508962 367392 508980 367414
rect 509014 367414 509070 367426
rect 509014 367392 509028 367414
rect 508962 367380 509028 367392
rect 509062 367392 509070 367414
rect 509104 367414 509160 367426
rect 509194 367414 509250 367426
rect 509284 367414 509340 367426
rect 509104 367392 509128 367414
rect 509194 367392 509228 367414
rect 509284 367392 509328 367414
rect 509374 367392 509435 367426
rect 509062 367380 509128 367392
rect 509162 367380 509228 367392
rect 509262 367380 509328 367392
rect 509362 367380 509435 367392
rect 508741 367336 509435 367380
rect 508741 367302 508800 367336
rect 508834 367314 508890 367336
rect 508862 367302 508890 367314
rect 508924 367314 508980 367336
rect 508924 367302 508928 367314
rect 508741 367280 508828 367302
rect 508862 367280 508928 367302
rect 508962 367302 508980 367314
rect 509014 367314 509070 367336
rect 509014 367302 509028 367314
rect 508962 367280 509028 367302
rect 509062 367302 509070 367314
rect 509104 367314 509160 367336
rect 509194 367314 509250 367336
rect 509284 367314 509340 367336
rect 509104 367302 509128 367314
rect 509194 367302 509228 367314
rect 509284 367302 509328 367314
rect 509374 367302 509435 367336
rect 509062 367280 509128 367302
rect 509162 367280 509228 367302
rect 509262 367280 509328 367302
rect 509362 367280 509435 367302
rect 508741 367246 509435 367280
rect 508741 367212 508800 367246
rect 508834 367214 508890 367246
rect 508862 367212 508890 367214
rect 508924 367214 508980 367246
rect 508924 367212 508928 367214
rect 508741 367180 508828 367212
rect 508862 367180 508928 367212
rect 508962 367212 508980 367214
rect 509014 367214 509070 367246
rect 509014 367212 509028 367214
rect 508962 367180 509028 367212
rect 509062 367212 509070 367214
rect 509104 367214 509160 367246
rect 509194 367214 509250 367246
rect 509284 367214 509340 367246
rect 509104 367212 509128 367214
rect 509194 367212 509228 367214
rect 509284 367212 509328 367214
rect 509374 367212 509435 367246
rect 509062 367180 509128 367212
rect 509162 367180 509228 367212
rect 509262 367180 509328 367212
rect 509362 367180 509435 367212
rect 508741 367156 509435 367180
rect 508741 367122 508800 367156
rect 508834 367122 508890 367156
rect 508924 367122 508980 367156
rect 509014 367122 509070 367156
rect 509104 367122 509160 367156
rect 509194 367122 509250 367156
rect 509284 367122 509340 367156
rect 509374 367122 509435 367156
rect 508741 367114 509435 367122
rect 508741 367080 508828 367114
rect 508862 367080 508928 367114
rect 508962 367080 509028 367114
rect 509062 367080 509128 367114
rect 509162 367080 509228 367114
rect 509262 367080 509328 367114
rect 509362 367080 509435 367114
rect 508741 367066 509435 367080
rect 508741 367032 508800 367066
rect 508834 367032 508890 367066
rect 508924 367032 508980 367066
rect 509014 367032 509070 367066
rect 509104 367032 509160 367066
rect 509194 367032 509250 367066
rect 509284 367032 509340 367066
rect 509374 367032 509435 367066
rect 508741 367014 509435 367032
rect 508741 366980 508828 367014
rect 508862 366980 508928 367014
rect 508962 366980 509028 367014
rect 509062 366980 509128 367014
rect 509162 366980 509228 367014
rect 509262 366980 509328 367014
rect 509362 366980 509435 367014
rect 508741 366976 509435 366980
rect 508741 366942 508800 366976
rect 508834 366942 508890 366976
rect 508924 366942 508980 366976
rect 509014 366942 509070 366976
rect 509104 366942 509160 366976
rect 509194 366942 509250 366976
rect 509284 366942 509340 366976
rect 509374 366942 509435 366976
rect 508741 366914 509435 366942
rect 508741 366886 508828 366914
rect 508862 366886 508928 366914
rect 508741 366852 508800 366886
rect 508862 366880 508890 366886
rect 508834 366852 508890 366880
rect 508924 366880 508928 366886
rect 508962 366886 509028 366914
rect 508962 366880 508980 366886
rect 508924 366852 508980 366880
rect 509014 366880 509028 366886
rect 509062 366886 509128 366914
rect 509162 366886 509228 366914
rect 509262 366886 509328 366914
rect 509362 366886 509435 366914
rect 509062 366880 509070 366886
rect 509014 366852 509070 366880
rect 509104 366880 509128 366886
rect 509194 366880 509228 366886
rect 509284 366880 509328 366886
rect 509104 366852 509160 366880
rect 509194 366852 509250 366880
rect 509284 366852 509340 366880
rect 509374 366852 509435 366886
rect 508741 366793 509435 366852
rect 509497 367434 509569 367490
rect 509497 367400 509516 367434
rect 509550 367400 509569 367434
rect 509497 367344 509569 367400
rect 509497 367310 509516 367344
rect 509550 367310 509569 367344
rect 509497 367254 509569 367310
rect 509497 367220 509516 367254
rect 509550 367220 509569 367254
rect 509497 367164 509569 367220
rect 509497 367130 509516 367164
rect 509550 367130 509569 367164
rect 509497 367074 509569 367130
rect 509497 367040 509516 367074
rect 509550 367040 509569 367074
rect 509497 366984 509569 367040
rect 509497 366950 509516 366984
rect 509550 366950 509569 366984
rect 509497 366894 509569 366950
rect 509497 366860 509516 366894
rect 509550 366860 509569 366894
rect 509497 366804 509569 366860
rect 508607 366756 508624 366790
rect 508658 366770 508679 366790
rect 508607 366736 508626 366756
rect 508660 366736 508679 366770
rect 508607 366731 508679 366736
rect 509497 366770 509516 366804
rect 509550 366770 509569 366804
rect 509497 366731 509569 366770
rect 508607 366712 509569 366731
rect 508607 366700 508702 366712
rect 508607 366666 508624 366700
rect 508658 366678 508702 366700
rect 508736 366678 508792 366712
rect 508826 366678 508882 366712
rect 508916 366678 508972 366712
rect 509006 366678 509062 366712
rect 509096 366678 509152 366712
rect 509186 366678 509242 366712
rect 509276 366678 509332 366712
rect 509366 366678 509422 366712
rect 509456 366678 509569 366712
rect 508658 366666 509569 366678
rect 508607 366659 509569 366666
rect 509633 367620 509666 367654
rect 509700 367620 509732 367654
rect 509633 367564 509732 367620
rect 509633 367530 509666 367564
rect 509700 367530 509732 367564
rect 509633 367474 509732 367530
rect 509633 367440 509666 367474
rect 509700 367440 509732 367474
rect 509633 367384 509732 367440
rect 509633 367350 509666 367384
rect 509700 367350 509732 367384
rect 509633 367294 509732 367350
rect 509633 367260 509666 367294
rect 509700 367260 509732 367294
rect 509633 367204 509732 367260
rect 509633 367170 509666 367204
rect 509700 367170 509732 367204
rect 509633 367114 509732 367170
rect 509633 367080 509666 367114
rect 509700 367080 509732 367114
rect 509633 367024 509732 367080
rect 509633 366990 509666 367024
rect 509700 366990 509732 367024
rect 509633 366934 509732 366990
rect 509633 366900 509666 366934
rect 509700 366900 509732 366934
rect 509633 366844 509732 366900
rect 509633 366810 509666 366844
rect 509700 366810 509732 366844
rect 509633 366754 509732 366810
rect 509633 366720 509666 366754
rect 509700 366720 509732 366754
rect 509633 366664 509732 366720
rect 508444 366595 508543 366630
rect 509633 366630 509666 366664
rect 509700 366630 509732 366664
rect 509633 366595 509732 366630
rect 508444 366594 509732 366595
rect 508444 366560 508464 366594
rect 508498 366563 509732 366594
rect 508498 366560 508502 366563
rect 508444 366529 508502 366560
rect 508536 366529 508592 366563
rect 508626 366529 508682 366563
rect 508716 366529 508772 366563
rect 508806 366529 508862 366563
rect 508896 366529 508952 366563
rect 508986 366529 509042 366563
rect 509076 366529 509132 366563
rect 509166 366529 509222 366563
rect 509256 366529 509312 366563
rect 509346 366529 509402 366563
rect 509436 366529 509492 366563
rect 509526 366529 509582 366563
rect 509616 366529 509732 366563
rect 508444 366424 509732 366529
rect 508444 366390 508464 366424
rect 508498 366410 509732 366424
rect 508498 366390 508502 366410
rect 508444 366376 508502 366390
rect 508536 366376 508592 366410
rect 508626 366376 508682 366410
rect 508716 366376 508772 366410
rect 508806 366376 508862 366410
rect 508896 366376 508952 366410
rect 508986 366376 509042 366410
rect 509076 366376 509132 366410
rect 509166 366376 509222 366410
rect 509256 366376 509312 366410
rect 509346 366376 509402 366410
rect 509436 366376 509492 366410
rect 509526 366376 509582 366410
rect 509616 366376 509732 366410
rect 508444 366345 509732 366376
rect 508444 366334 508543 366345
rect 508444 366300 508464 366334
rect 508498 366314 508543 366334
rect 508444 366280 508479 366300
rect 508513 366280 508543 366314
rect 509633 366314 509732 366345
rect 508444 366244 508543 366280
rect 508444 366210 508464 366244
rect 508498 366224 508543 366244
rect 508444 366190 508479 366210
rect 508513 366190 508543 366224
rect 508444 366154 508543 366190
rect 508444 366120 508464 366154
rect 508498 366134 508543 366154
rect 508444 366100 508479 366120
rect 508513 366100 508543 366134
rect 508444 366064 508543 366100
rect 508444 366030 508464 366064
rect 508498 366044 508543 366064
rect 508444 366010 508479 366030
rect 508513 366010 508543 366044
rect 508444 365974 508543 366010
rect 508444 365940 508464 365974
rect 508498 365954 508543 365974
rect 508444 365920 508479 365940
rect 508513 365920 508543 365954
rect 508444 365884 508543 365920
rect 508444 365850 508464 365884
rect 508498 365864 508543 365884
rect 508444 365830 508479 365850
rect 508513 365830 508543 365864
rect 508444 365794 508543 365830
rect 508444 365760 508464 365794
rect 508498 365774 508543 365794
rect 508444 365740 508479 365760
rect 508513 365740 508543 365774
rect 508444 365704 508543 365740
rect 508444 365670 508464 365704
rect 508498 365684 508543 365704
rect 508444 365650 508479 365670
rect 508513 365650 508543 365684
rect 508444 365614 508543 365650
rect 508444 365580 508464 365614
rect 508498 365594 508543 365614
rect 508444 365560 508479 365580
rect 508513 365560 508543 365594
rect 508444 365524 508543 365560
rect 508444 365490 508464 365524
rect 508498 365504 508543 365524
rect 508444 365470 508479 365490
rect 508513 365470 508543 365504
rect 508444 365434 508543 365470
rect 508444 365400 508464 365434
rect 508498 365414 508543 365434
rect 508444 365380 508479 365400
rect 508513 365380 508543 365414
rect 508444 365344 508543 365380
rect 508444 365310 508464 365344
rect 508498 365324 508543 365344
rect 508444 365290 508479 365310
rect 508513 365290 508543 365324
rect 508607 366262 509569 366281
rect 508607 366260 508683 366262
rect 508607 366226 508624 366260
rect 508658 366228 508683 366260
rect 508717 366228 508773 366262
rect 508807 366228 508863 366262
rect 508897 366228 508953 366262
rect 508987 366228 509043 366262
rect 509077 366228 509133 366262
rect 509167 366228 509223 366262
rect 509257 366228 509313 366262
rect 509347 366228 509403 366262
rect 509437 366228 509569 366262
rect 508658 366226 509569 366228
rect 508607 366209 509569 366226
rect 508607 366170 508679 366209
rect 508607 366136 508624 366170
rect 508658 366150 508679 366170
rect 508607 366116 508626 366136
rect 508660 366116 508679 366150
rect 509497 366184 509569 366209
rect 509497 366150 509516 366184
rect 509550 366150 509569 366184
rect 508607 366080 508679 366116
rect 508607 366046 508624 366080
rect 508658 366060 508679 366080
rect 508607 366026 508626 366046
rect 508660 366026 508679 366060
rect 508607 365990 508679 366026
rect 508607 365956 508624 365990
rect 508658 365970 508679 365990
rect 508607 365936 508626 365956
rect 508660 365936 508679 365970
rect 508607 365900 508679 365936
rect 508607 365866 508624 365900
rect 508658 365880 508679 365900
rect 508607 365846 508626 365866
rect 508660 365846 508679 365880
rect 508607 365810 508679 365846
rect 508607 365776 508624 365810
rect 508658 365790 508679 365810
rect 508607 365756 508626 365776
rect 508660 365756 508679 365790
rect 508607 365720 508679 365756
rect 508607 365686 508624 365720
rect 508658 365700 508679 365720
rect 508607 365666 508626 365686
rect 508660 365666 508679 365700
rect 508607 365630 508679 365666
rect 508607 365596 508624 365630
rect 508658 365610 508679 365630
rect 508607 365576 508626 365596
rect 508660 365576 508679 365610
rect 508607 365540 508679 365576
rect 508607 365506 508624 365540
rect 508658 365520 508679 365540
rect 508607 365486 508626 365506
rect 508660 365486 508679 365520
rect 508607 365450 508679 365486
rect 508741 366086 509435 366147
rect 508741 366052 508800 366086
rect 508834 366074 508890 366086
rect 508862 366052 508890 366074
rect 508924 366074 508980 366086
rect 508924 366052 508928 366074
rect 508741 366040 508828 366052
rect 508862 366040 508928 366052
rect 508962 366052 508980 366074
rect 509014 366074 509070 366086
rect 509014 366052 509028 366074
rect 508962 366040 509028 366052
rect 509062 366052 509070 366074
rect 509104 366074 509160 366086
rect 509194 366074 509250 366086
rect 509284 366074 509340 366086
rect 509104 366052 509128 366074
rect 509194 366052 509228 366074
rect 509284 366052 509328 366074
rect 509374 366052 509435 366086
rect 509062 366040 509128 366052
rect 509162 366040 509228 366052
rect 509262 366040 509328 366052
rect 509362 366040 509435 366052
rect 508741 365996 509435 366040
rect 508741 365962 508800 365996
rect 508834 365974 508890 365996
rect 508862 365962 508890 365974
rect 508924 365974 508980 365996
rect 508924 365962 508928 365974
rect 508741 365940 508828 365962
rect 508862 365940 508928 365962
rect 508962 365962 508980 365974
rect 509014 365974 509070 365996
rect 509014 365962 509028 365974
rect 508962 365940 509028 365962
rect 509062 365962 509070 365974
rect 509104 365974 509160 365996
rect 509194 365974 509250 365996
rect 509284 365974 509340 365996
rect 509104 365962 509128 365974
rect 509194 365962 509228 365974
rect 509284 365962 509328 365974
rect 509374 365962 509435 365996
rect 509062 365940 509128 365962
rect 509162 365940 509228 365962
rect 509262 365940 509328 365962
rect 509362 365940 509435 365962
rect 508741 365906 509435 365940
rect 508741 365872 508800 365906
rect 508834 365874 508890 365906
rect 508862 365872 508890 365874
rect 508924 365874 508980 365906
rect 508924 365872 508928 365874
rect 508741 365840 508828 365872
rect 508862 365840 508928 365872
rect 508962 365872 508980 365874
rect 509014 365874 509070 365906
rect 509014 365872 509028 365874
rect 508962 365840 509028 365872
rect 509062 365872 509070 365874
rect 509104 365874 509160 365906
rect 509194 365874 509250 365906
rect 509284 365874 509340 365906
rect 509104 365872 509128 365874
rect 509194 365872 509228 365874
rect 509284 365872 509328 365874
rect 509374 365872 509435 365906
rect 509062 365840 509128 365872
rect 509162 365840 509228 365872
rect 509262 365840 509328 365872
rect 509362 365840 509435 365872
rect 508741 365816 509435 365840
rect 508741 365782 508800 365816
rect 508834 365782 508890 365816
rect 508924 365782 508980 365816
rect 509014 365782 509070 365816
rect 509104 365782 509160 365816
rect 509194 365782 509250 365816
rect 509284 365782 509340 365816
rect 509374 365782 509435 365816
rect 508741 365774 509435 365782
rect 508741 365740 508828 365774
rect 508862 365740 508928 365774
rect 508962 365740 509028 365774
rect 509062 365740 509128 365774
rect 509162 365740 509228 365774
rect 509262 365740 509328 365774
rect 509362 365740 509435 365774
rect 508741 365726 509435 365740
rect 508741 365692 508800 365726
rect 508834 365692 508890 365726
rect 508924 365692 508980 365726
rect 509014 365692 509070 365726
rect 509104 365692 509160 365726
rect 509194 365692 509250 365726
rect 509284 365692 509340 365726
rect 509374 365692 509435 365726
rect 508741 365674 509435 365692
rect 508741 365640 508828 365674
rect 508862 365640 508928 365674
rect 508962 365640 509028 365674
rect 509062 365640 509128 365674
rect 509162 365640 509228 365674
rect 509262 365640 509328 365674
rect 509362 365640 509435 365674
rect 508741 365636 509435 365640
rect 508741 365602 508800 365636
rect 508834 365602 508890 365636
rect 508924 365602 508980 365636
rect 509014 365602 509070 365636
rect 509104 365602 509160 365636
rect 509194 365602 509250 365636
rect 509284 365602 509340 365636
rect 509374 365602 509435 365636
rect 508741 365574 509435 365602
rect 508741 365546 508828 365574
rect 508862 365546 508928 365574
rect 508741 365512 508800 365546
rect 508862 365540 508890 365546
rect 508834 365512 508890 365540
rect 508924 365540 508928 365546
rect 508962 365546 509028 365574
rect 508962 365540 508980 365546
rect 508924 365512 508980 365540
rect 509014 365540 509028 365546
rect 509062 365546 509128 365574
rect 509162 365546 509228 365574
rect 509262 365546 509328 365574
rect 509362 365546 509435 365574
rect 509062 365540 509070 365546
rect 509014 365512 509070 365540
rect 509104 365540 509128 365546
rect 509194 365540 509228 365546
rect 509284 365540 509328 365546
rect 509104 365512 509160 365540
rect 509194 365512 509250 365540
rect 509284 365512 509340 365540
rect 509374 365512 509435 365546
rect 508741 365453 509435 365512
rect 509497 366094 509569 366150
rect 509497 366060 509516 366094
rect 509550 366060 509569 366094
rect 509497 366004 509569 366060
rect 509497 365970 509516 366004
rect 509550 365970 509569 366004
rect 509497 365914 509569 365970
rect 509497 365880 509516 365914
rect 509550 365880 509569 365914
rect 509497 365824 509569 365880
rect 509497 365790 509516 365824
rect 509550 365790 509569 365824
rect 509497 365734 509569 365790
rect 509497 365700 509516 365734
rect 509550 365700 509569 365734
rect 509497 365644 509569 365700
rect 509497 365610 509516 365644
rect 509550 365610 509569 365644
rect 509497 365554 509569 365610
rect 509497 365520 509516 365554
rect 509550 365520 509569 365554
rect 509497 365464 509569 365520
rect 508607 365416 508624 365450
rect 508658 365430 508679 365450
rect 508607 365396 508626 365416
rect 508660 365396 508679 365430
rect 508607 365391 508679 365396
rect 509497 365430 509516 365464
rect 509550 365430 509569 365464
rect 509497 365391 509569 365430
rect 508607 365372 509569 365391
rect 508607 365360 508702 365372
rect 508607 365326 508624 365360
rect 508658 365338 508702 365360
rect 508736 365338 508792 365372
rect 508826 365338 508882 365372
rect 508916 365338 508972 365372
rect 509006 365338 509062 365372
rect 509096 365338 509152 365372
rect 509186 365338 509242 365372
rect 509276 365338 509332 365372
rect 509366 365338 509422 365372
rect 509456 365338 509569 365372
rect 508658 365326 509569 365338
rect 508607 365319 509569 365326
rect 509633 366280 509666 366314
rect 509700 366280 509732 366314
rect 509633 366224 509732 366280
rect 509633 366190 509666 366224
rect 509700 366190 509732 366224
rect 509633 366134 509732 366190
rect 509633 366100 509666 366134
rect 509700 366100 509732 366134
rect 509633 366044 509732 366100
rect 509633 366010 509666 366044
rect 509700 366010 509732 366044
rect 509633 365954 509732 366010
rect 509633 365920 509666 365954
rect 509700 365920 509732 365954
rect 509633 365864 509732 365920
rect 509633 365830 509666 365864
rect 509700 365830 509732 365864
rect 509633 365774 509732 365830
rect 509633 365740 509666 365774
rect 509700 365740 509732 365774
rect 509633 365684 509732 365740
rect 509633 365650 509666 365684
rect 509700 365650 509732 365684
rect 509633 365594 509732 365650
rect 509633 365560 509666 365594
rect 509700 365560 509732 365594
rect 509633 365504 509732 365560
rect 509633 365470 509666 365504
rect 509700 365470 509732 365504
rect 509633 365414 509732 365470
rect 509633 365380 509666 365414
rect 509700 365380 509732 365414
rect 509633 365324 509732 365380
rect 508444 365255 508543 365290
rect 509633 365290 509666 365324
rect 509700 365290 509732 365324
rect 509633 365255 509732 365290
rect 508444 365254 509732 365255
rect 508444 365220 508464 365254
rect 508498 365223 509732 365254
rect 508498 365220 508502 365223
rect 508444 365189 508502 365220
rect 508536 365189 508592 365223
rect 508626 365189 508682 365223
rect 508716 365189 508772 365223
rect 508806 365189 508862 365223
rect 508896 365189 508952 365223
rect 508986 365189 509042 365223
rect 509076 365189 509132 365223
rect 509166 365189 509222 365223
rect 509256 365189 509312 365223
rect 509346 365189 509402 365223
rect 509436 365189 509492 365223
rect 509526 365189 509582 365223
rect 509616 365189 509732 365223
rect 508444 365084 509732 365189
rect 508444 365050 508464 365084
rect 508498 365070 509732 365084
rect 508498 365050 508502 365070
rect 508444 365036 508502 365050
rect 508536 365036 508592 365070
rect 508626 365036 508682 365070
rect 508716 365036 508772 365070
rect 508806 365036 508862 365070
rect 508896 365036 508952 365070
rect 508986 365036 509042 365070
rect 509076 365036 509132 365070
rect 509166 365036 509222 365070
rect 509256 365036 509312 365070
rect 509346 365036 509402 365070
rect 509436 365036 509492 365070
rect 509526 365036 509582 365070
rect 509616 365036 509732 365070
rect 508444 365005 509732 365036
rect 508444 364994 508543 365005
rect 508444 364960 508464 364994
rect 508498 364974 508543 364994
rect 508444 364940 508479 364960
rect 508513 364940 508543 364974
rect 509633 364974 509732 365005
rect 508444 364904 508543 364940
rect 508444 364870 508464 364904
rect 508498 364884 508543 364904
rect 508444 364850 508479 364870
rect 508513 364850 508543 364884
rect 508444 364814 508543 364850
rect 508444 364780 508464 364814
rect 508498 364794 508543 364814
rect 508444 364760 508479 364780
rect 508513 364760 508543 364794
rect 508444 364724 508543 364760
rect 508444 364690 508464 364724
rect 508498 364704 508543 364724
rect 508444 364670 508479 364690
rect 508513 364670 508543 364704
rect 508444 364634 508543 364670
rect 508444 364600 508464 364634
rect 508498 364614 508543 364634
rect 508444 364580 508479 364600
rect 508513 364580 508543 364614
rect 508444 364544 508543 364580
rect 508444 364510 508464 364544
rect 508498 364524 508543 364544
rect 508444 364490 508479 364510
rect 508513 364490 508543 364524
rect 508444 364454 508543 364490
rect 508444 364420 508464 364454
rect 508498 364434 508543 364454
rect 508444 364400 508479 364420
rect 508513 364400 508543 364434
rect 508444 364364 508543 364400
rect 508444 364330 508464 364364
rect 508498 364344 508543 364364
rect 508444 364310 508479 364330
rect 508513 364310 508543 364344
rect 508444 364274 508543 364310
rect 508444 364240 508464 364274
rect 508498 364254 508543 364274
rect 508444 364220 508479 364240
rect 508513 364220 508543 364254
rect 508444 364184 508543 364220
rect 508444 364150 508464 364184
rect 508498 364164 508543 364184
rect 508444 364130 508479 364150
rect 508513 364130 508543 364164
rect 508444 364094 508543 364130
rect 508444 364060 508464 364094
rect 508498 364074 508543 364094
rect 508444 364040 508479 364060
rect 508513 364040 508543 364074
rect 508444 364004 508543 364040
rect 508444 363970 508464 364004
rect 508498 363984 508543 364004
rect 508444 363950 508479 363970
rect 508513 363950 508543 363984
rect 508607 364922 509569 364941
rect 508607 364920 508683 364922
rect 508607 364886 508624 364920
rect 508658 364888 508683 364920
rect 508717 364888 508773 364922
rect 508807 364888 508863 364922
rect 508897 364888 508953 364922
rect 508987 364888 509043 364922
rect 509077 364888 509133 364922
rect 509167 364888 509223 364922
rect 509257 364888 509313 364922
rect 509347 364888 509403 364922
rect 509437 364888 509569 364922
rect 508658 364886 509569 364888
rect 508607 364869 509569 364886
rect 508607 364830 508679 364869
rect 508607 364796 508624 364830
rect 508658 364810 508679 364830
rect 508607 364776 508626 364796
rect 508660 364776 508679 364810
rect 509497 364844 509569 364869
rect 509497 364810 509516 364844
rect 509550 364810 509569 364844
rect 508607 364740 508679 364776
rect 508607 364706 508624 364740
rect 508658 364720 508679 364740
rect 508607 364686 508626 364706
rect 508660 364686 508679 364720
rect 508607 364650 508679 364686
rect 508607 364616 508624 364650
rect 508658 364630 508679 364650
rect 508607 364596 508626 364616
rect 508660 364596 508679 364630
rect 508607 364560 508679 364596
rect 508607 364526 508624 364560
rect 508658 364540 508679 364560
rect 508607 364506 508626 364526
rect 508660 364506 508679 364540
rect 508607 364470 508679 364506
rect 508607 364436 508624 364470
rect 508658 364450 508679 364470
rect 508607 364416 508626 364436
rect 508660 364416 508679 364450
rect 508607 364380 508679 364416
rect 508607 364346 508624 364380
rect 508658 364360 508679 364380
rect 508607 364326 508626 364346
rect 508660 364326 508679 364360
rect 508607 364290 508679 364326
rect 508607 364256 508624 364290
rect 508658 364270 508679 364290
rect 508607 364236 508626 364256
rect 508660 364236 508679 364270
rect 508607 364200 508679 364236
rect 508607 364166 508624 364200
rect 508658 364180 508679 364200
rect 508607 364146 508626 364166
rect 508660 364146 508679 364180
rect 508607 364110 508679 364146
rect 508741 364746 509435 364807
rect 508741 364712 508800 364746
rect 508834 364734 508890 364746
rect 508862 364712 508890 364734
rect 508924 364734 508980 364746
rect 508924 364712 508928 364734
rect 508741 364700 508828 364712
rect 508862 364700 508928 364712
rect 508962 364712 508980 364734
rect 509014 364734 509070 364746
rect 509014 364712 509028 364734
rect 508962 364700 509028 364712
rect 509062 364712 509070 364734
rect 509104 364734 509160 364746
rect 509194 364734 509250 364746
rect 509284 364734 509340 364746
rect 509104 364712 509128 364734
rect 509194 364712 509228 364734
rect 509284 364712 509328 364734
rect 509374 364712 509435 364746
rect 509062 364700 509128 364712
rect 509162 364700 509228 364712
rect 509262 364700 509328 364712
rect 509362 364700 509435 364712
rect 508741 364656 509435 364700
rect 508741 364622 508800 364656
rect 508834 364634 508890 364656
rect 508862 364622 508890 364634
rect 508924 364634 508980 364656
rect 508924 364622 508928 364634
rect 508741 364600 508828 364622
rect 508862 364600 508928 364622
rect 508962 364622 508980 364634
rect 509014 364634 509070 364656
rect 509014 364622 509028 364634
rect 508962 364600 509028 364622
rect 509062 364622 509070 364634
rect 509104 364634 509160 364656
rect 509194 364634 509250 364656
rect 509284 364634 509340 364656
rect 509104 364622 509128 364634
rect 509194 364622 509228 364634
rect 509284 364622 509328 364634
rect 509374 364622 509435 364656
rect 509062 364600 509128 364622
rect 509162 364600 509228 364622
rect 509262 364600 509328 364622
rect 509362 364600 509435 364622
rect 508741 364566 509435 364600
rect 508741 364532 508800 364566
rect 508834 364534 508890 364566
rect 508862 364532 508890 364534
rect 508924 364534 508980 364566
rect 508924 364532 508928 364534
rect 508741 364500 508828 364532
rect 508862 364500 508928 364532
rect 508962 364532 508980 364534
rect 509014 364534 509070 364566
rect 509014 364532 509028 364534
rect 508962 364500 509028 364532
rect 509062 364532 509070 364534
rect 509104 364534 509160 364566
rect 509194 364534 509250 364566
rect 509284 364534 509340 364566
rect 509104 364532 509128 364534
rect 509194 364532 509228 364534
rect 509284 364532 509328 364534
rect 509374 364532 509435 364566
rect 509062 364500 509128 364532
rect 509162 364500 509228 364532
rect 509262 364500 509328 364532
rect 509362 364500 509435 364532
rect 508741 364476 509435 364500
rect 508741 364442 508800 364476
rect 508834 364442 508890 364476
rect 508924 364442 508980 364476
rect 509014 364442 509070 364476
rect 509104 364442 509160 364476
rect 509194 364442 509250 364476
rect 509284 364442 509340 364476
rect 509374 364442 509435 364476
rect 508741 364434 509435 364442
rect 508741 364400 508828 364434
rect 508862 364400 508928 364434
rect 508962 364400 509028 364434
rect 509062 364400 509128 364434
rect 509162 364400 509228 364434
rect 509262 364400 509328 364434
rect 509362 364400 509435 364434
rect 508741 364386 509435 364400
rect 508741 364352 508800 364386
rect 508834 364352 508890 364386
rect 508924 364352 508980 364386
rect 509014 364352 509070 364386
rect 509104 364352 509160 364386
rect 509194 364352 509250 364386
rect 509284 364352 509340 364386
rect 509374 364352 509435 364386
rect 508741 364334 509435 364352
rect 508741 364300 508828 364334
rect 508862 364300 508928 364334
rect 508962 364300 509028 364334
rect 509062 364300 509128 364334
rect 509162 364300 509228 364334
rect 509262 364300 509328 364334
rect 509362 364300 509435 364334
rect 508741 364296 509435 364300
rect 508741 364262 508800 364296
rect 508834 364262 508890 364296
rect 508924 364262 508980 364296
rect 509014 364262 509070 364296
rect 509104 364262 509160 364296
rect 509194 364262 509250 364296
rect 509284 364262 509340 364296
rect 509374 364262 509435 364296
rect 508741 364234 509435 364262
rect 508741 364206 508828 364234
rect 508862 364206 508928 364234
rect 508741 364172 508800 364206
rect 508862 364200 508890 364206
rect 508834 364172 508890 364200
rect 508924 364200 508928 364206
rect 508962 364206 509028 364234
rect 508962 364200 508980 364206
rect 508924 364172 508980 364200
rect 509014 364200 509028 364206
rect 509062 364206 509128 364234
rect 509162 364206 509228 364234
rect 509262 364206 509328 364234
rect 509362 364206 509435 364234
rect 509062 364200 509070 364206
rect 509014 364172 509070 364200
rect 509104 364200 509128 364206
rect 509194 364200 509228 364206
rect 509284 364200 509328 364206
rect 509104 364172 509160 364200
rect 509194 364172 509250 364200
rect 509284 364172 509340 364200
rect 509374 364172 509435 364206
rect 508741 364113 509435 364172
rect 509497 364754 509569 364810
rect 509497 364720 509516 364754
rect 509550 364720 509569 364754
rect 509497 364664 509569 364720
rect 509497 364630 509516 364664
rect 509550 364630 509569 364664
rect 509497 364574 509569 364630
rect 509497 364540 509516 364574
rect 509550 364540 509569 364574
rect 509497 364484 509569 364540
rect 509497 364450 509516 364484
rect 509550 364450 509569 364484
rect 509497 364394 509569 364450
rect 509497 364360 509516 364394
rect 509550 364360 509569 364394
rect 509497 364304 509569 364360
rect 509497 364270 509516 364304
rect 509550 364270 509569 364304
rect 509497 364214 509569 364270
rect 509497 364180 509516 364214
rect 509550 364180 509569 364214
rect 509497 364124 509569 364180
rect 508607 364076 508624 364110
rect 508658 364090 508679 364110
rect 508607 364056 508626 364076
rect 508660 364056 508679 364090
rect 508607 364051 508679 364056
rect 509497 364090 509516 364124
rect 509550 364090 509569 364124
rect 509497 364051 509569 364090
rect 508607 364032 509569 364051
rect 508607 364020 508702 364032
rect 508607 363986 508624 364020
rect 508658 363998 508702 364020
rect 508736 363998 508792 364032
rect 508826 363998 508882 364032
rect 508916 363998 508972 364032
rect 509006 363998 509062 364032
rect 509096 363998 509152 364032
rect 509186 363998 509242 364032
rect 509276 363998 509332 364032
rect 509366 363998 509422 364032
rect 509456 363998 509569 364032
rect 508658 363986 509569 363998
rect 508607 363979 509569 363986
rect 509633 364940 509666 364974
rect 509700 364940 509732 364974
rect 509633 364884 509732 364940
rect 509633 364850 509666 364884
rect 509700 364850 509732 364884
rect 509633 364794 509732 364850
rect 509633 364760 509666 364794
rect 509700 364760 509732 364794
rect 509633 364704 509732 364760
rect 509633 364670 509666 364704
rect 509700 364670 509732 364704
rect 509633 364614 509732 364670
rect 509633 364580 509666 364614
rect 509700 364580 509732 364614
rect 509633 364524 509732 364580
rect 509633 364490 509666 364524
rect 509700 364490 509732 364524
rect 509633 364434 509732 364490
rect 509633 364400 509666 364434
rect 509700 364400 509732 364434
rect 509633 364344 509732 364400
rect 509633 364310 509666 364344
rect 509700 364310 509732 364344
rect 509633 364254 509732 364310
rect 509633 364220 509666 364254
rect 509700 364220 509732 364254
rect 509633 364164 509732 364220
rect 509633 364130 509666 364164
rect 509700 364130 509732 364164
rect 509633 364074 509732 364130
rect 509633 364040 509666 364074
rect 509700 364040 509732 364074
rect 509633 363984 509732 364040
rect 508444 363915 508543 363950
rect 509633 363950 509666 363984
rect 509700 363950 509732 363984
rect 509633 363915 509732 363950
rect 508444 363914 509732 363915
rect 508444 363880 508464 363914
rect 508498 363883 509732 363914
rect 508498 363880 508502 363883
rect 508444 363849 508502 363880
rect 508536 363849 508592 363883
rect 508626 363849 508682 363883
rect 508716 363849 508772 363883
rect 508806 363849 508862 363883
rect 508896 363849 508952 363883
rect 508986 363849 509042 363883
rect 509076 363849 509132 363883
rect 509166 363849 509222 363883
rect 509256 363849 509312 363883
rect 509346 363849 509402 363883
rect 509436 363849 509492 363883
rect 509526 363849 509582 363883
rect 509616 363849 509732 363883
rect 508444 363744 509732 363849
rect 508444 363710 508464 363744
rect 508498 363730 509732 363744
rect 508498 363710 508502 363730
rect 508444 363696 508502 363710
rect 508536 363696 508592 363730
rect 508626 363696 508682 363730
rect 508716 363696 508772 363730
rect 508806 363696 508862 363730
rect 508896 363696 508952 363730
rect 508986 363696 509042 363730
rect 509076 363696 509132 363730
rect 509166 363696 509222 363730
rect 509256 363696 509312 363730
rect 509346 363696 509402 363730
rect 509436 363696 509492 363730
rect 509526 363696 509582 363730
rect 509616 363696 509732 363730
rect 508444 363665 509732 363696
rect 508444 363654 508543 363665
rect 508444 363620 508464 363654
rect 508498 363634 508543 363654
rect 508444 363600 508479 363620
rect 508513 363600 508543 363634
rect 509633 363634 509732 363665
rect 508444 363564 508543 363600
rect 508444 363530 508464 363564
rect 508498 363544 508543 363564
rect 508444 363510 508479 363530
rect 508513 363510 508543 363544
rect 508444 363474 508543 363510
rect 508444 363440 508464 363474
rect 508498 363454 508543 363474
rect 508444 363420 508479 363440
rect 508513 363420 508543 363454
rect 508444 363384 508543 363420
rect 508444 363350 508464 363384
rect 508498 363364 508543 363384
rect 508444 363330 508479 363350
rect 508513 363330 508543 363364
rect 508444 363294 508543 363330
rect 508444 363260 508464 363294
rect 508498 363274 508543 363294
rect 508444 363240 508479 363260
rect 508513 363240 508543 363274
rect 508444 363204 508543 363240
rect 508444 363170 508464 363204
rect 508498 363184 508543 363204
rect 508444 363150 508479 363170
rect 508513 363150 508543 363184
rect 508444 363114 508543 363150
rect 508444 363080 508464 363114
rect 508498 363094 508543 363114
rect 508444 363060 508479 363080
rect 508513 363060 508543 363094
rect 508444 363024 508543 363060
rect 508444 362990 508464 363024
rect 508498 363004 508543 363024
rect 508444 362970 508479 362990
rect 508513 362970 508543 363004
rect 508444 362934 508543 362970
rect 508444 362900 508464 362934
rect 508498 362914 508543 362934
rect 508444 362880 508479 362900
rect 508513 362880 508543 362914
rect 508444 362844 508543 362880
rect 508444 362810 508464 362844
rect 508498 362824 508543 362844
rect 508444 362790 508479 362810
rect 508513 362790 508543 362824
rect 508444 362754 508543 362790
rect 508444 362720 508464 362754
rect 508498 362734 508543 362754
rect 508444 362700 508479 362720
rect 508513 362700 508543 362734
rect 508444 362664 508543 362700
rect 508444 362630 508464 362664
rect 508498 362644 508543 362664
rect 508444 362610 508479 362630
rect 508513 362610 508543 362644
rect 508607 363582 509569 363601
rect 508607 363580 508683 363582
rect 508607 363546 508624 363580
rect 508658 363548 508683 363580
rect 508717 363548 508773 363582
rect 508807 363548 508863 363582
rect 508897 363548 508953 363582
rect 508987 363548 509043 363582
rect 509077 363548 509133 363582
rect 509167 363548 509223 363582
rect 509257 363548 509313 363582
rect 509347 363548 509403 363582
rect 509437 363548 509569 363582
rect 508658 363546 509569 363548
rect 508607 363529 509569 363546
rect 508607 363490 508679 363529
rect 508607 363456 508624 363490
rect 508658 363470 508679 363490
rect 508607 363436 508626 363456
rect 508660 363436 508679 363470
rect 509497 363504 509569 363529
rect 509497 363470 509516 363504
rect 509550 363470 509569 363504
rect 508607 363400 508679 363436
rect 508607 363366 508624 363400
rect 508658 363380 508679 363400
rect 508607 363346 508626 363366
rect 508660 363346 508679 363380
rect 508607 363310 508679 363346
rect 508607 363276 508624 363310
rect 508658 363290 508679 363310
rect 508607 363256 508626 363276
rect 508660 363256 508679 363290
rect 508607 363220 508679 363256
rect 508607 363186 508624 363220
rect 508658 363200 508679 363220
rect 508607 363166 508626 363186
rect 508660 363166 508679 363200
rect 508607 363130 508679 363166
rect 508607 363096 508624 363130
rect 508658 363110 508679 363130
rect 508607 363076 508626 363096
rect 508660 363076 508679 363110
rect 508607 363040 508679 363076
rect 508607 363006 508624 363040
rect 508658 363020 508679 363040
rect 508607 362986 508626 363006
rect 508660 362986 508679 363020
rect 508607 362950 508679 362986
rect 508607 362916 508624 362950
rect 508658 362930 508679 362950
rect 508607 362896 508626 362916
rect 508660 362896 508679 362930
rect 508607 362860 508679 362896
rect 508607 362826 508624 362860
rect 508658 362840 508679 362860
rect 508607 362806 508626 362826
rect 508660 362806 508679 362840
rect 508607 362770 508679 362806
rect 508741 363406 509435 363467
rect 508741 363372 508800 363406
rect 508834 363394 508890 363406
rect 508862 363372 508890 363394
rect 508924 363394 508980 363406
rect 508924 363372 508928 363394
rect 508741 363360 508828 363372
rect 508862 363360 508928 363372
rect 508962 363372 508980 363394
rect 509014 363394 509070 363406
rect 509014 363372 509028 363394
rect 508962 363360 509028 363372
rect 509062 363372 509070 363394
rect 509104 363394 509160 363406
rect 509194 363394 509250 363406
rect 509284 363394 509340 363406
rect 509104 363372 509128 363394
rect 509194 363372 509228 363394
rect 509284 363372 509328 363394
rect 509374 363372 509435 363406
rect 509062 363360 509128 363372
rect 509162 363360 509228 363372
rect 509262 363360 509328 363372
rect 509362 363360 509435 363372
rect 508741 363316 509435 363360
rect 508741 363282 508800 363316
rect 508834 363294 508890 363316
rect 508862 363282 508890 363294
rect 508924 363294 508980 363316
rect 508924 363282 508928 363294
rect 508741 363260 508828 363282
rect 508862 363260 508928 363282
rect 508962 363282 508980 363294
rect 509014 363294 509070 363316
rect 509014 363282 509028 363294
rect 508962 363260 509028 363282
rect 509062 363282 509070 363294
rect 509104 363294 509160 363316
rect 509194 363294 509250 363316
rect 509284 363294 509340 363316
rect 509104 363282 509128 363294
rect 509194 363282 509228 363294
rect 509284 363282 509328 363294
rect 509374 363282 509435 363316
rect 509062 363260 509128 363282
rect 509162 363260 509228 363282
rect 509262 363260 509328 363282
rect 509362 363260 509435 363282
rect 508741 363226 509435 363260
rect 508741 363192 508800 363226
rect 508834 363194 508890 363226
rect 508862 363192 508890 363194
rect 508924 363194 508980 363226
rect 508924 363192 508928 363194
rect 508741 363160 508828 363192
rect 508862 363160 508928 363192
rect 508962 363192 508980 363194
rect 509014 363194 509070 363226
rect 509014 363192 509028 363194
rect 508962 363160 509028 363192
rect 509062 363192 509070 363194
rect 509104 363194 509160 363226
rect 509194 363194 509250 363226
rect 509284 363194 509340 363226
rect 509104 363192 509128 363194
rect 509194 363192 509228 363194
rect 509284 363192 509328 363194
rect 509374 363192 509435 363226
rect 509062 363160 509128 363192
rect 509162 363160 509228 363192
rect 509262 363160 509328 363192
rect 509362 363160 509435 363192
rect 508741 363136 509435 363160
rect 508741 363102 508800 363136
rect 508834 363102 508890 363136
rect 508924 363102 508980 363136
rect 509014 363102 509070 363136
rect 509104 363102 509160 363136
rect 509194 363102 509250 363136
rect 509284 363102 509340 363136
rect 509374 363102 509435 363136
rect 508741 363094 509435 363102
rect 508741 363060 508828 363094
rect 508862 363060 508928 363094
rect 508962 363060 509028 363094
rect 509062 363060 509128 363094
rect 509162 363060 509228 363094
rect 509262 363060 509328 363094
rect 509362 363060 509435 363094
rect 508741 363046 509435 363060
rect 508741 363012 508800 363046
rect 508834 363012 508890 363046
rect 508924 363012 508980 363046
rect 509014 363012 509070 363046
rect 509104 363012 509160 363046
rect 509194 363012 509250 363046
rect 509284 363012 509340 363046
rect 509374 363012 509435 363046
rect 508741 362994 509435 363012
rect 508741 362960 508828 362994
rect 508862 362960 508928 362994
rect 508962 362960 509028 362994
rect 509062 362960 509128 362994
rect 509162 362960 509228 362994
rect 509262 362960 509328 362994
rect 509362 362960 509435 362994
rect 508741 362956 509435 362960
rect 508741 362922 508800 362956
rect 508834 362922 508890 362956
rect 508924 362922 508980 362956
rect 509014 362922 509070 362956
rect 509104 362922 509160 362956
rect 509194 362922 509250 362956
rect 509284 362922 509340 362956
rect 509374 362922 509435 362956
rect 508741 362894 509435 362922
rect 508741 362866 508828 362894
rect 508862 362866 508928 362894
rect 508741 362832 508800 362866
rect 508862 362860 508890 362866
rect 508834 362832 508890 362860
rect 508924 362860 508928 362866
rect 508962 362866 509028 362894
rect 508962 362860 508980 362866
rect 508924 362832 508980 362860
rect 509014 362860 509028 362866
rect 509062 362866 509128 362894
rect 509162 362866 509228 362894
rect 509262 362866 509328 362894
rect 509362 362866 509435 362894
rect 509062 362860 509070 362866
rect 509014 362832 509070 362860
rect 509104 362860 509128 362866
rect 509194 362860 509228 362866
rect 509284 362860 509328 362866
rect 509104 362832 509160 362860
rect 509194 362832 509250 362860
rect 509284 362832 509340 362860
rect 509374 362832 509435 362866
rect 508741 362773 509435 362832
rect 509497 363414 509569 363470
rect 509497 363380 509516 363414
rect 509550 363380 509569 363414
rect 509497 363324 509569 363380
rect 509497 363290 509516 363324
rect 509550 363290 509569 363324
rect 509497 363234 509569 363290
rect 509497 363200 509516 363234
rect 509550 363200 509569 363234
rect 509497 363144 509569 363200
rect 509497 363110 509516 363144
rect 509550 363110 509569 363144
rect 509497 363054 509569 363110
rect 509497 363020 509516 363054
rect 509550 363020 509569 363054
rect 509497 362964 509569 363020
rect 509497 362930 509516 362964
rect 509550 362930 509569 362964
rect 509497 362874 509569 362930
rect 509497 362840 509516 362874
rect 509550 362840 509569 362874
rect 509497 362784 509569 362840
rect 508607 362736 508624 362770
rect 508658 362750 508679 362770
rect 508607 362716 508626 362736
rect 508660 362716 508679 362750
rect 508607 362711 508679 362716
rect 509497 362750 509516 362784
rect 509550 362750 509569 362784
rect 509497 362711 509569 362750
rect 508607 362692 509569 362711
rect 508607 362680 508702 362692
rect 508607 362646 508624 362680
rect 508658 362658 508702 362680
rect 508736 362658 508792 362692
rect 508826 362658 508882 362692
rect 508916 362658 508972 362692
rect 509006 362658 509062 362692
rect 509096 362658 509152 362692
rect 509186 362658 509242 362692
rect 509276 362658 509332 362692
rect 509366 362658 509422 362692
rect 509456 362658 509569 362692
rect 508658 362646 509569 362658
rect 508607 362639 509569 362646
rect 509633 363600 509666 363634
rect 509700 363600 509732 363634
rect 509633 363544 509732 363600
rect 509633 363510 509666 363544
rect 509700 363510 509732 363544
rect 509633 363454 509732 363510
rect 509633 363420 509666 363454
rect 509700 363420 509732 363454
rect 509633 363364 509732 363420
rect 509633 363330 509666 363364
rect 509700 363330 509732 363364
rect 509633 363274 509732 363330
rect 509633 363240 509666 363274
rect 509700 363240 509732 363274
rect 509633 363184 509732 363240
rect 509633 363150 509666 363184
rect 509700 363150 509732 363184
rect 509633 363094 509732 363150
rect 509633 363060 509666 363094
rect 509700 363060 509732 363094
rect 509633 363004 509732 363060
rect 509633 362970 509666 363004
rect 509700 362970 509732 363004
rect 509633 362914 509732 362970
rect 509633 362880 509666 362914
rect 509700 362880 509732 362914
rect 509633 362824 509732 362880
rect 509633 362790 509666 362824
rect 509700 362790 509732 362824
rect 509633 362734 509732 362790
rect 509633 362700 509666 362734
rect 509700 362700 509732 362734
rect 509633 362644 509732 362700
rect 508444 362575 508543 362610
rect 509633 362610 509666 362644
rect 509700 362610 509732 362644
rect 509633 362575 509732 362610
rect 508444 362574 509732 362575
rect 508444 362540 508464 362574
rect 508498 362543 509732 362574
rect 508498 362540 508502 362543
rect 508444 362509 508502 362540
rect 508536 362509 508592 362543
rect 508626 362509 508682 362543
rect 508716 362509 508772 362543
rect 508806 362509 508862 362543
rect 508896 362509 508952 362543
rect 508986 362509 509042 362543
rect 509076 362509 509132 362543
rect 509166 362509 509222 362543
rect 509256 362509 509312 362543
rect 509346 362509 509402 362543
rect 509436 362509 509492 362543
rect 509526 362509 509582 362543
rect 509616 362509 509732 362543
rect 508444 362476 509732 362509
rect 509998 372987 510058 373170
rect 509998 372953 510011 372987
rect 510045 372953 510058 372987
rect 509998 372787 510058 372953
rect 509998 372753 510011 372787
rect 510045 372753 510058 372787
rect 509998 372587 510058 372753
rect 509998 372553 510011 372587
rect 510045 372553 510058 372587
rect 509998 372387 510058 372553
rect 509998 372353 510011 372387
rect 510045 372353 510058 372387
rect 509998 372187 510058 372353
rect 509998 372153 510011 372187
rect 510045 372153 510058 372187
rect 509998 371987 510058 372153
rect 509998 371953 510011 371987
rect 510045 371953 510058 371987
rect 509998 371787 510058 371953
rect 509998 371753 510011 371787
rect 510045 371753 510058 371787
rect 509998 371587 510058 371753
rect 509998 371553 510011 371587
rect 510045 371553 510058 371587
rect 509998 371387 510058 371553
rect 509998 371353 510011 371387
rect 510045 371353 510058 371387
rect 509998 371187 510058 371353
rect 509998 371153 510011 371187
rect 510045 371153 510058 371187
rect 509998 370987 510058 371153
rect 509998 370953 510011 370987
rect 510045 370953 510058 370987
rect 509998 370787 510058 370953
rect 509998 370753 510011 370787
rect 510045 370753 510058 370787
rect 509998 370587 510058 370753
rect 509998 370553 510011 370587
rect 510045 370553 510058 370587
rect 509998 370387 510058 370553
rect 509998 370353 510011 370387
rect 510045 370353 510058 370387
rect 509998 370187 510058 370353
rect 509998 370153 510011 370187
rect 510045 370153 510058 370187
rect 509998 369987 510058 370153
rect 509998 369953 510011 369987
rect 510045 369953 510058 369987
rect 509998 369787 510058 369953
rect 509998 369753 510011 369787
rect 510045 369753 510058 369787
rect 509998 369587 510058 369753
rect 509998 369553 510011 369587
rect 510045 369553 510058 369587
rect 509998 369387 510058 369553
rect 509998 369353 510011 369387
rect 510045 369353 510058 369387
rect 509998 369187 510058 369353
rect 509998 369153 510011 369187
rect 510045 369153 510058 369187
rect 509998 368987 510058 369153
rect 509998 368953 510011 368987
rect 510045 368953 510058 368987
rect 509998 368787 510058 368953
rect 509998 368753 510011 368787
rect 510045 368753 510058 368787
rect 509998 368587 510058 368753
rect 509998 368553 510011 368587
rect 510045 368553 510058 368587
rect 509998 368387 510058 368553
rect 509998 368353 510011 368387
rect 510045 368353 510058 368387
rect 509998 368187 510058 368353
rect 509998 368153 510011 368187
rect 510045 368153 510058 368187
rect 509998 367987 510058 368153
rect 509998 367953 510011 367987
rect 510045 367953 510058 367987
rect 509998 367787 510058 367953
rect 509998 367753 510011 367787
rect 510045 367753 510058 367787
rect 509998 367587 510058 367753
rect 509998 367553 510011 367587
rect 510045 367553 510058 367587
rect 509998 367387 510058 367553
rect 509998 367353 510011 367387
rect 510045 367353 510058 367387
rect 509998 367187 510058 367353
rect 509998 367153 510011 367187
rect 510045 367153 510058 367187
rect 509998 366987 510058 367153
rect 509998 366953 510011 366987
rect 510045 366953 510058 366987
rect 509998 366787 510058 366953
rect 509998 366753 510011 366787
rect 510045 366753 510058 366787
rect 509998 366587 510058 366753
rect 509998 366553 510011 366587
rect 510045 366553 510058 366587
rect 509998 366387 510058 366553
rect 509998 366353 510011 366387
rect 510045 366353 510058 366387
rect 509998 366187 510058 366353
rect 509998 366153 510011 366187
rect 510045 366153 510058 366187
rect 509998 365987 510058 366153
rect 509998 365953 510011 365987
rect 510045 365953 510058 365987
rect 509998 365787 510058 365953
rect 509998 365753 510011 365787
rect 510045 365753 510058 365787
rect 509998 365587 510058 365753
rect 509998 365553 510011 365587
rect 510045 365553 510058 365587
rect 509998 365387 510058 365553
rect 509998 365353 510011 365387
rect 510045 365353 510058 365387
rect 509998 365187 510058 365353
rect 509998 365153 510011 365187
rect 510045 365153 510058 365187
rect 509998 364987 510058 365153
rect 509998 364953 510011 364987
rect 510045 364953 510058 364987
rect 509998 364787 510058 364953
rect 509998 364753 510011 364787
rect 510045 364753 510058 364787
rect 509998 364587 510058 364753
rect 509998 364553 510011 364587
rect 510045 364553 510058 364587
rect 509998 364387 510058 364553
rect 509998 364353 510011 364387
rect 510045 364353 510058 364387
rect 509998 364187 510058 364353
rect 509998 364153 510011 364187
rect 510045 364153 510058 364187
rect 509998 363987 510058 364153
rect 509998 363953 510011 363987
rect 510045 363953 510058 363987
rect 509998 363787 510058 363953
rect 509998 363753 510011 363787
rect 510045 363753 510058 363787
rect 509998 363587 510058 363753
rect 509998 363553 510011 363587
rect 510045 363553 510058 363587
rect 509998 363387 510058 363553
rect 509998 363353 510011 363387
rect 510045 363353 510058 363387
rect 509998 363187 510058 363353
rect 509998 363153 510011 363187
rect 510045 363153 510058 363187
rect 509998 362987 510058 363153
rect 509998 362953 510011 362987
rect 510045 362953 510058 362987
rect 509998 362787 510058 362953
rect 509998 362753 510011 362787
rect 510045 362753 510058 362787
rect 509998 362587 510058 362753
rect 509998 362553 510011 362587
rect 510045 362553 510058 362587
rect 509998 362450 510058 362553
rect 511878 372987 511938 373170
rect 511878 372953 511891 372987
rect 511925 372953 511938 372987
rect 511878 372787 511938 372953
rect 511878 372753 511891 372787
rect 511925 372753 511938 372787
rect 511878 372587 511938 372753
rect 511878 372553 511891 372587
rect 511925 372553 511938 372587
rect 511878 372387 511938 372553
rect 511878 372353 511891 372387
rect 511925 372353 511938 372387
rect 511878 372187 511938 372353
rect 511878 372153 511891 372187
rect 511925 372153 511938 372187
rect 511878 371987 511938 372153
rect 511878 371953 511891 371987
rect 511925 371953 511938 371987
rect 511878 371787 511938 371953
rect 511878 371753 511891 371787
rect 511925 371753 511938 371787
rect 511878 371587 511938 371753
rect 511878 371553 511891 371587
rect 511925 371553 511938 371587
rect 511878 371387 511938 371553
rect 511878 371353 511891 371387
rect 511925 371353 511938 371387
rect 511878 371187 511938 371353
rect 511878 371153 511891 371187
rect 511925 371153 511938 371187
rect 511878 370987 511938 371153
rect 511878 370953 511891 370987
rect 511925 370953 511938 370987
rect 511878 370787 511938 370953
rect 511878 370753 511891 370787
rect 511925 370753 511938 370787
rect 511878 370587 511938 370753
rect 511878 370553 511891 370587
rect 511925 370553 511938 370587
rect 511878 370387 511938 370553
rect 511878 370353 511891 370387
rect 511925 370353 511938 370387
rect 511878 370187 511938 370353
rect 511878 370153 511891 370187
rect 511925 370153 511938 370187
rect 511878 369987 511938 370153
rect 511878 369953 511891 369987
rect 511925 369953 511938 369987
rect 511878 369787 511938 369953
rect 511878 369753 511891 369787
rect 511925 369753 511938 369787
rect 511878 369587 511938 369753
rect 511878 369553 511891 369587
rect 511925 369553 511938 369587
rect 511878 369387 511938 369553
rect 511878 369353 511891 369387
rect 511925 369353 511938 369387
rect 511878 369187 511938 369353
rect 511878 369153 511891 369187
rect 511925 369153 511938 369187
rect 511878 368987 511938 369153
rect 511878 368953 511891 368987
rect 511925 368953 511938 368987
rect 511878 368787 511938 368953
rect 511878 368753 511891 368787
rect 511925 368753 511938 368787
rect 511878 368587 511938 368753
rect 511878 368553 511891 368587
rect 511925 368553 511938 368587
rect 511878 368387 511938 368553
rect 511878 368353 511891 368387
rect 511925 368353 511938 368387
rect 511878 368187 511938 368353
rect 511878 368153 511891 368187
rect 511925 368153 511938 368187
rect 511878 367987 511938 368153
rect 511878 367953 511891 367987
rect 511925 367953 511938 367987
rect 511878 367787 511938 367953
rect 511878 367753 511891 367787
rect 511925 367753 511938 367787
rect 511878 367587 511938 367753
rect 511878 367553 511891 367587
rect 511925 367553 511938 367587
rect 511878 367387 511938 367553
rect 511878 367353 511891 367387
rect 511925 367353 511938 367387
rect 511878 367187 511938 367353
rect 511878 367153 511891 367187
rect 511925 367153 511938 367187
rect 511878 366987 511938 367153
rect 511878 366953 511891 366987
rect 511925 366953 511938 366987
rect 511878 366787 511938 366953
rect 511878 366753 511891 366787
rect 511925 366753 511938 366787
rect 511878 366587 511938 366753
rect 511878 366553 511891 366587
rect 511925 366553 511938 366587
rect 511878 366387 511938 366553
rect 511878 366353 511891 366387
rect 511925 366353 511938 366387
rect 511878 366187 511938 366353
rect 511878 366153 511891 366187
rect 511925 366153 511938 366187
rect 511878 365987 511938 366153
rect 511878 365953 511891 365987
rect 511925 365953 511938 365987
rect 511878 365787 511938 365953
rect 511878 365753 511891 365787
rect 511925 365753 511938 365787
rect 511878 365587 511938 365753
rect 511878 365553 511891 365587
rect 511925 365553 511938 365587
rect 511878 365387 511938 365553
rect 511878 365353 511891 365387
rect 511925 365353 511938 365387
rect 511878 365187 511938 365353
rect 511878 365153 511891 365187
rect 511925 365153 511938 365187
rect 511878 364987 511938 365153
rect 511878 364953 511891 364987
rect 511925 364953 511938 364987
rect 511878 364787 511938 364953
rect 511878 364753 511891 364787
rect 511925 364753 511938 364787
rect 511878 364587 511938 364753
rect 511878 364553 511891 364587
rect 511925 364553 511938 364587
rect 511878 364387 511938 364553
rect 511878 364353 511891 364387
rect 511925 364353 511938 364387
rect 511878 364187 511938 364353
rect 511878 364153 511891 364187
rect 511925 364153 511938 364187
rect 511878 363987 511938 364153
rect 511878 363953 511891 363987
rect 511925 363953 511938 363987
rect 511878 363787 511938 363953
rect 511878 363753 511891 363787
rect 511925 363753 511938 363787
rect 511878 363587 511938 363753
rect 511878 363553 511891 363587
rect 511925 363553 511938 363587
rect 511878 363387 511938 363553
rect 511878 363353 511891 363387
rect 511925 363353 511938 363387
rect 511878 363187 511938 363353
rect 511878 363153 511891 363187
rect 511925 363153 511938 363187
rect 511878 362987 511938 363153
rect 511878 362953 511891 362987
rect 511925 362953 511938 362987
rect 511878 362787 511938 362953
rect 511878 362753 511891 362787
rect 511925 362753 511938 362787
rect 511878 362587 511938 362753
rect 511878 362553 511891 362587
rect 511925 362553 511938 362587
rect 511878 362450 511938 362553
rect 512204 373124 513492 373144
rect 512204 373090 512224 373124
rect 512258 373110 513492 373124
rect 512258 373090 512262 373110
rect 512204 373076 512262 373090
rect 512296 373076 512352 373110
rect 512386 373076 512442 373110
rect 512476 373076 512532 373110
rect 512566 373076 512622 373110
rect 512656 373076 512712 373110
rect 512746 373076 512802 373110
rect 512836 373076 512892 373110
rect 512926 373076 512982 373110
rect 513016 373076 513072 373110
rect 513106 373076 513162 373110
rect 513196 373076 513252 373110
rect 513286 373076 513342 373110
rect 513376 373076 513492 373110
rect 512204 373045 513492 373076
rect 512204 373034 512303 373045
rect 512204 373000 512224 373034
rect 512258 373014 512303 373034
rect 512204 372980 512239 373000
rect 512273 372980 512303 373014
rect 513393 373014 513492 373045
rect 512204 372944 512303 372980
rect 512204 372910 512224 372944
rect 512258 372924 512303 372944
rect 512204 372890 512239 372910
rect 512273 372890 512303 372924
rect 512204 372854 512303 372890
rect 512204 372820 512224 372854
rect 512258 372834 512303 372854
rect 512204 372800 512239 372820
rect 512273 372800 512303 372834
rect 512204 372764 512303 372800
rect 512204 372730 512224 372764
rect 512258 372744 512303 372764
rect 512204 372710 512239 372730
rect 512273 372710 512303 372744
rect 512204 372674 512303 372710
rect 512204 372640 512224 372674
rect 512258 372654 512303 372674
rect 512204 372620 512239 372640
rect 512273 372620 512303 372654
rect 512204 372584 512303 372620
rect 512204 372550 512224 372584
rect 512258 372564 512303 372584
rect 512204 372530 512239 372550
rect 512273 372530 512303 372564
rect 512204 372494 512303 372530
rect 512204 372460 512224 372494
rect 512258 372474 512303 372494
rect 512204 372440 512239 372460
rect 512273 372440 512303 372474
rect 512204 372404 512303 372440
rect 512204 372370 512224 372404
rect 512258 372384 512303 372404
rect 512204 372350 512239 372370
rect 512273 372350 512303 372384
rect 512204 372314 512303 372350
rect 512204 372280 512224 372314
rect 512258 372294 512303 372314
rect 512204 372260 512239 372280
rect 512273 372260 512303 372294
rect 512204 372224 512303 372260
rect 512204 372190 512224 372224
rect 512258 372204 512303 372224
rect 512204 372170 512239 372190
rect 512273 372170 512303 372204
rect 512204 372134 512303 372170
rect 512204 372100 512224 372134
rect 512258 372114 512303 372134
rect 512204 372080 512239 372100
rect 512273 372080 512303 372114
rect 512204 372044 512303 372080
rect 512204 372010 512224 372044
rect 512258 372024 512303 372044
rect 512204 371990 512239 372010
rect 512273 371990 512303 372024
rect 512367 372962 513329 372981
rect 512367 372960 512443 372962
rect 512367 372926 512384 372960
rect 512418 372928 512443 372960
rect 512477 372928 512533 372962
rect 512567 372928 512623 372962
rect 512657 372928 512713 372962
rect 512747 372928 512803 372962
rect 512837 372928 512893 372962
rect 512927 372928 512983 372962
rect 513017 372928 513073 372962
rect 513107 372928 513163 372962
rect 513197 372928 513329 372962
rect 512418 372926 513329 372928
rect 512367 372909 513329 372926
rect 512367 372870 512439 372909
rect 512367 372836 512384 372870
rect 512418 372850 512439 372870
rect 512367 372816 512386 372836
rect 512420 372816 512439 372850
rect 513257 372884 513329 372909
rect 513257 372850 513276 372884
rect 513310 372850 513329 372884
rect 512367 372780 512439 372816
rect 512367 372746 512384 372780
rect 512418 372760 512439 372780
rect 512367 372726 512386 372746
rect 512420 372726 512439 372760
rect 512367 372690 512439 372726
rect 512367 372656 512384 372690
rect 512418 372670 512439 372690
rect 512367 372636 512386 372656
rect 512420 372636 512439 372670
rect 512367 372600 512439 372636
rect 512367 372566 512384 372600
rect 512418 372580 512439 372600
rect 512367 372546 512386 372566
rect 512420 372546 512439 372580
rect 512367 372510 512439 372546
rect 512367 372476 512384 372510
rect 512418 372490 512439 372510
rect 512367 372456 512386 372476
rect 512420 372456 512439 372490
rect 512367 372420 512439 372456
rect 512367 372386 512384 372420
rect 512418 372400 512439 372420
rect 512367 372366 512386 372386
rect 512420 372366 512439 372400
rect 512367 372330 512439 372366
rect 512367 372296 512384 372330
rect 512418 372310 512439 372330
rect 512367 372276 512386 372296
rect 512420 372276 512439 372310
rect 512367 372240 512439 372276
rect 512367 372206 512384 372240
rect 512418 372220 512439 372240
rect 512367 372186 512386 372206
rect 512420 372186 512439 372220
rect 512367 372150 512439 372186
rect 512501 372786 513195 372847
rect 512501 372752 512560 372786
rect 512594 372774 512650 372786
rect 512622 372752 512650 372774
rect 512684 372774 512740 372786
rect 512684 372752 512688 372774
rect 512501 372740 512588 372752
rect 512622 372740 512688 372752
rect 512722 372752 512740 372774
rect 512774 372774 512830 372786
rect 512774 372752 512788 372774
rect 512722 372740 512788 372752
rect 512822 372752 512830 372774
rect 512864 372774 512920 372786
rect 512954 372774 513010 372786
rect 513044 372774 513100 372786
rect 512864 372752 512888 372774
rect 512954 372752 512988 372774
rect 513044 372752 513088 372774
rect 513134 372752 513195 372786
rect 512822 372740 512888 372752
rect 512922 372740 512988 372752
rect 513022 372740 513088 372752
rect 513122 372740 513195 372752
rect 512501 372696 513195 372740
rect 512501 372662 512560 372696
rect 512594 372674 512650 372696
rect 512622 372662 512650 372674
rect 512684 372674 512740 372696
rect 512684 372662 512688 372674
rect 512501 372640 512588 372662
rect 512622 372640 512688 372662
rect 512722 372662 512740 372674
rect 512774 372674 512830 372696
rect 512774 372662 512788 372674
rect 512722 372640 512788 372662
rect 512822 372662 512830 372674
rect 512864 372674 512920 372696
rect 512954 372674 513010 372696
rect 513044 372674 513100 372696
rect 512864 372662 512888 372674
rect 512954 372662 512988 372674
rect 513044 372662 513088 372674
rect 513134 372662 513195 372696
rect 512822 372640 512888 372662
rect 512922 372640 512988 372662
rect 513022 372640 513088 372662
rect 513122 372640 513195 372662
rect 512501 372606 513195 372640
rect 512501 372572 512560 372606
rect 512594 372574 512650 372606
rect 512622 372572 512650 372574
rect 512684 372574 512740 372606
rect 512684 372572 512688 372574
rect 512501 372540 512588 372572
rect 512622 372540 512688 372572
rect 512722 372572 512740 372574
rect 512774 372574 512830 372606
rect 512774 372572 512788 372574
rect 512722 372540 512788 372572
rect 512822 372572 512830 372574
rect 512864 372574 512920 372606
rect 512954 372574 513010 372606
rect 513044 372574 513100 372606
rect 512864 372572 512888 372574
rect 512954 372572 512988 372574
rect 513044 372572 513088 372574
rect 513134 372572 513195 372606
rect 512822 372540 512888 372572
rect 512922 372540 512988 372572
rect 513022 372540 513088 372572
rect 513122 372540 513195 372572
rect 512501 372516 513195 372540
rect 512501 372482 512560 372516
rect 512594 372482 512650 372516
rect 512684 372482 512740 372516
rect 512774 372482 512830 372516
rect 512864 372482 512920 372516
rect 512954 372482 513010 372516
rect 513044 372482 513100 372516
rect 513134 372482 513195 372516
rect 512501 372474 513195 372482
rect 512501 372440 512588 372474
rect 512622 372440 512688 372474
rect 512722 372440 512788 372474
rect 512822 372440 512888 372474
rect 512922 372440 512988 372474
rect 513022 372440 513088 372474
rect 513122 372440 513195 372474
rect 512501 372426 513195 372440
rect 512501 372392 512560 372426
rect 512594 372392 512650 372426
rect 512684 372392 512740 372426
rect 512774 372392 512830 372426
rect 512864 372392 512920 372426
rect 512954 372392 513010 372426
rect 513044 372392 513100 372426
rect 513134 372392 513195 372426
rect 512501 372374 513195 372392
rect 512501 372340 512588 372374
rect 512622 372340 512688 372374
rect 512722 372340 512788 372374
rect 512822 372340 512888 372374
rect 512922 372340 512988 372374
rect 513022 372340 513088 372374
rect 513122 372340 513195 372374
rect 512501 372336 513195 372340
rect 512501 372302 512560 372336
rect 512594 372302 512650 372336
rect 512684 372302 512740 372336
rect 512774 372302 512830 372336
rect 512864 372302 512920 372336
rect 512954 372302 513010 372336
rect 513044 372302 513100 372336
rect 513134 372302 513195 372336
rect 512501 372274 513195 372302
rect 512501 372246 512588 372274
rect 512622 372246 512688 372274
rect 512501 372212 512560 372246
rect 512622 372240 512650 372246
rect 512594 372212 512650 372240
rect 512684 372240 512688 372246
rect 512722 372246 512788 372274
rect 512722 372240 512740 372246
rect 512684 372212 512740 372240
rect 512774 372240 512788 372246
rect 512822 372246 512888 372274
rect 512922 372246 512988 372274
rect 513022 372246 513088 372274
rect 513122 372246 513195 372274
rect 512822 372240 512830 372246
rect 512774 372212 512830 372240
rect 512864 372240 512888 372246
rect 512954 372240 512988 372246
rect 513044 372240 513088 372246
rect 512864 372212 512920 372240
rect 512954 372212 513010 372240
rect 513044 372212 513100 372240
rect 513134 372212 513195 372246
rect 512501 372153 513195 372212
rect 513257 372794 513329 372850
rect 513257 372760 513276 372794
rect 513310 372760 513329 372794
rect 513257 372704 513329 372760
rect 513257 372670 513276 372704
rect 513310 372670 513329 372704
rect 513257 372614 513329 372670
rect 513257 372580 513276 372614
rect 513310 372580 513329 372614
rect 513257 372524 513329 372580
rect 513257 372490 513276 372524
rect 513310 372490 513329 372524
rect 513257 372434 513329 372490
rect 513257 372400 513276 372434
rect 513310 372400 513329 372434
rect 513257 372344 513329 372400
rect 513257 372310 513276 372344
rect 513310 372310 513329 372344
rect 513257 372254 513329 372310
rect 513257 372220 513276 372254
rect 513310 372220 513329 372254
rect 513257 372164 513329 372220
rect 512367 372116 512384 372150
rect 512418 372130 512439 372150
rect 512367 372096 512386 372116
rect 512420 372096 512439 372130
rect 512367 372091 512439 372096
rect 513257 372130 513276 372164
rect 513310 372130 513329 372164
rect 513257 372091 513329 372130
rect 512367 372072 513329 372091
rect 512367 372060 512462 372072
rect 512367 372026 512384 372060
rect 512418 372038 512462 372060
rect 512496 372038 512552 372072
rect 512586 372038 512642 372072
rect 512676 372038 512732 372072
rect 512766 372038 512822 372072
rect 512856 372038 512912 372072
rect 512946 372038 513002 372072
rect 513036 372038 513092 372072
rect 513126 372038 513182 372072
rect 513216 372038 513329 372072
rect 512418 372026 513329 372038
rect 512367 372019 513329 372026
rect 513393 372980 513426 373014
rect 513460 372980 513492 373014
rect 513393 372924 513492 372980
rect 513393 372890 513426 372924
rect 513460 372890 513492 372924
rect 513393 372834 513492 372890
rect 513393 372800 513426 372834
rect 513460 372800 513492 372834
rect 513393 372744 513492 372800
rect 513393 372710 513426 372744
rect 513460 372710 513492 372744
rect 513393 372654 513492 372710
rect 513393 372620 513426 372654
rect 513460 372620 513492 372654
rect 513393 372564 513492 372620
rect 513393 372530 513426 372564
rect 513460 372530 513492 372564
rect 513393 372474 513492 372530
rect 513393 372440 513426 372474
rect 513460 372440 513492 372474
rect 513393 372384 513492 372440
rect 513393 372350 513426 372384
rect 513460 372350 513492 372384
rect 513393 372294 513492 372350
rect 513393 372260 513426 372294
rect 513460 372260 513492 372294
rect 513393 372204 513492 372260
rect 513393 372170 513426 372204
rect 513460 372170 513492 372204
rect 513393 372114 513492 372170
rect 513393 372080 513426 372114
rect 513460 372080 513492 372114
rect 513393 372024 513492 372080
rect 512204 371955 512303 371990
rect 513393 371990 513426 372024
rect 513460 371990 513492 372024
rect 513393 371955 513492 371990
rect 512204 371954 513492 371955
rect 512204 371920 512224 371954
rect 512258 371923 513492 371954
rect 512258 371920 512262 371923
rect 512204 371889 512262 371920
rect 512296 371889 512352 371923
rect 512386 371889 512442 371923
rect 512476 371889 512532 371923
rect 512566 371889 512622 371923
rect 512656 371889 512712 371923
rect 512746 371889 512802 371923
rect 512836 371889 512892 371923
rect 512926 371889 512982 371923
rect 513016 371889 513072 371923
rect 513106 371889 513162 371923
rect 513196 371889 513252 371923
rect 513286 371889 513342 371923
rect 513376 371889 513492 371923
rect 512204 371784 513492 371889
rect 512204 371750 512224 371784
rect 512258 371770 513492 371784
rect 512258 371750 512262 371770
rect 512204 371736 512262 371750
rect 512296 371736 512352 371770
rect 512386 371736 512442 371770
rect 512476 371736 512532 371770
rect 512566 371736 512622 371770
rect 512656 371736 512712 371770
rect 512746 371736 512802 371770
rect 512836 371736 512892 371770
rect 512926 371736 512982 371770
rect 513016 371736 513072 371770
rect 513106 371736 513162 371770
rect 513196 371736 513252 371770
rect 513286 371736 513342 371770
rect 513376 371736 513492 371770
rect 512204 371705 513492 371736
rect 512204 371694 512303 371705
rect 512204 371660 512224 371694
rect 512258 371674 512303 371694
rect 512204 371640 512239 371660
rect 512273 371640 512303 371674
rect 513393 371674 513492 371705
rect 512204 371604 512303 371640
rect 512204 371570 512224 371604
rect 512258 371584 512303 371604
rect 512204 371550 512239 371570
rect 512273 371550 512303 371584
rect 512204 371514 512303 371550
rect 512204 371480 512224 371514
rect 512258 371494 512303 371514
rect 512204 371460 512239 371480
rect 512273 371460 512303 371494
rect 512204 371424 512303 371460
rect 512204 371390 512224 371424
rect 512258 371404 512303 371424
rect 512204 371370 512239 371390
rect 512273 371370 512303 371404
rect 512204 371334 512303 371370
rect 512204 371300 512224 371334
rect 512258 371314 512303 371334
rect 512204 371280 512239 371300
rect 512273 371280 512303 371314
rect 512204 371244 512303 371280
rect 512204 371210 512224 371244
rect 512258 371224 512303 371244
rect 512204 371190 512239 371210
rect 512273 371190 512303 371224
rect 512204 371154 512303 371190
rect 512204 371120 512224 371154
rect 512258 371134 512303 371154
rect 512204 371100 512239 371120
rect 512273 371100 512303 371134
rect 512204 371064 512303 371100
rect 512204 371030 512224 371064
rect 512258 371044 512303 371064
rect 512204 371010 512239 371030
rect 512273 371010 512303 371044
rect 512204 370974 512303 371010
rect 512204 370940 512224 370974
rect 512258 370954 512303 370974
rect 512204 370920 512239 370940
rect 512273 370920 512303 370954
rect 512204 370884 512303 370920
rect 512204 370850 512224 370884
rect 512258 370864 512303 370884
rect 512204 370830 512239 370850
rect 512273 370830 512303 370864
rect 512204 370794 512303 370830
rect 512204 370760 512224 370794
rect 512258 370774 512303 370794
rect 512204 370740 512239 370760
rect 512273 370740 512303 370774
rect 512204 370704 512303 370740
rect 512204 370670 512224 370704
rect 512258 370684 512303 370704
rect 512204 370650 512239 370670
rect 512273 370650 512303 370684
rect 512367 371622 513329 371641
rect 512367 371620 512443 371622
rect 512367 371586 512384 371620
rect 512418 371588 512443 371620
rect 512477 371588 512533 371622
rect 512567 371588 512623 371622
rect 512657 371588 512713 371622
rect 512747 371588 512803 371622
rect 512837 371588 512893 371622
rect 512927 371588 512983 371622
rect 513017 371588 513073 371622
rect 513107 371588 513163 371622
rect 513197 371588 513329 371622
rect 512418 371586 513329 371588
rect 512367 371569 513329 371586
rect 512367 371530 512439 371569
rect 512367 371496 512384 371530
rect 512418 371510 512439 371530
rect 512367 371476 512386 371496
rect 512420 371476 512439 371510
rect 513257 371544 513329 371569
rect 513257 371510 513276 371544
rect 513310 371510 513329 371544
rect 512367 371440 512439 371476
rect 512367 371406 512384 371440
rect 512418 371420 512439 371440
rect 512367 371386 512386 371406
rect 512420 371386 512439 371420
rect 512367 371350 512439 371386
rect 512367 371316 512384 371350
rect 512418 371330 512439 371350
rect 512367 371296 512386 371316
rect 512420 371296 512439 371330
rect 512367 371260 512439 371296
rect 512367 371226 512384 371260
rect 512418 371240 512439 371260
rect 512367 371206 512386 371226
rect 512420 371206 512439 371240
rect 512367 371170 512439 371206
rect 512367 371136 512384 371170
rect 512418 371150 512439 371170
rect 512367 371116 512386 371136
rect 512420 371116 512439 371150
rect 512367 371080 512439 371116
rect 512367 371046 512384 371080
rect 512418 371060 512439 371080
rect 512367 371026 512386 371046
rect 512420 371026 512439 371060
rect 512367 370990 512439 371026
rect 512367 370956 512384 370990
rect 512418 370970 512439 370990
rect 512367 370936 512386 370956
rect 512420 370936 512439 370970
rect 512367 370900 512439 370936
rect 512367 370866 512384 370900
rect 512418 370880 512439 370900
rect 512367 370846 512386 370866
rect 512420 370846 512439 370880
rect 512367 370810 512439 370846
rect 512501 371446 513195 371507
rect 512501 371412 512560 371446
rect 512594 371434 512650 371446
rect 512622 371412 512650 371434
rect 512684 371434 512740 371446
rect 512684 371412 512688 371434
rect 512501 371400 512588 371412
rect 512622 371400 512688 371412
rect 512722 371412 512740 371434
rect 512774 371434 512830 371446
rect 512774 371412 512788 371434
rect 512722 371400 512788 371412
rect 512822 371412 512830 371434
rect 512864 371434 512920 371446
rect 512954 371434 513010 371446
rect 513044 371434 513100 371446
rect 512864 371412 512888 371434
rect 512954 371412 512988 371434
rect 513044 371412 513088 371434
rect 513134 371412 513195 371446
rect 512822 371400 512888 371412
rect 512922 371400 512988 371412
rect 513022 371400 513088 371412
rect 513122 371400 513195 371412
rect 512501 371356 513195 371400
rect 512501 371322 512560 371356
rect 512594 371334 512650 371356
rect 512622 371322 512650 371334
rect 512684 371334 512740 371356
rect 512684 371322 512688 371334
rect 512501 371300 512588 371322
rect 512622 371300 512688 371322
rect 512722 371322 512740 371334
rect 512774 371334 512830 371356
rect 512774 371322 512788 371334
rect 512722 371300 512788 371322
rect 512822 371322 512830 371334
rect 512864 371334 512920 371356
rect 512954 371334 513010 371356
rect 513044 371334 513100 371356
rect 512864 371322 512888 371334
rect 512954 371322 512988 371334
rect 513044 371322 513088 371334
rect 513134 371322 513195 371356
rect 512822 371300 512888 371322
rect 512922 371300 512988 371322
rect 513022 371300 513088 371322
rect 513122 371300 513195 371322
rect 512501 371266 513195 371300
rect 512501 371232 512560 371266
rect 512594 371234 512650 371266
rect 512622 371232 512650 371234
rect 512684 371234 512740 371266
rect 512684 371232 512688 371234
rect 512501 371200 512588 371232
rect 512622 371200 512688 371232
rect 512722 371232 512740 371234
rect 512774 371234 512830 371266
rect 512774 371232 512788 371234
rect 512722 371200 512788 371232
rect 512822 371232 512830 371234
rect 512864 371234 512920 371266
rect 512954 371234 513010 371266
rect 513044 371234 513100 371266
rect 512864 371232 512888 371234
rect 512954 371232 512988 371234
rect 513044 371232 513088 371234
rect 513134 371232 513195 371266
rect 512822 371200 512888 371232
rect 512922 371200 512988 371232
rect 513022 371200 513088 371232
rect 513122 371200 513195 371232
rect 512501 371176 513195 371200
rect 512501 371142 512560 371176
rect 512594 371142 512650 371176
rect 512684 371142 512740 371176
rect 512774 371142 512830 371176
rect 512864 371142 512920 371176
rect 512954 371142 513010 371176
rect 513044 371142 513100 371176
rect 513134 371142 513195 371176
rect 512501 371134 513195 371142
rect 512501 371100 512588 371134
rect 512622 371100 512688 371134
rect 512722 371100 512788 371134
rect 512822 371100 512888 371134
rect 512922 371100 512988 371134
rect 513022 371100 513088 371134
rect 513122 371100 513195 371134
rect 512501 371086 513195 371100
rect 512501 371052 512560 371086
rect 512594 371052 512650 371086
rect 512684 371052 512740 371086
rect 512774 371052 512830 371086
rect 512864 371052 512920 371086
rect 512954 371052 513010 371086
rect 513044 371052 513100 371086
rect 513134 371052 513195 371086
rect 512501 371034 513195 371052
rect 512501 371000 512588 371034
rect 512622 371000 512688 371034
rect 512722 371000 512788 371034
rect 512822 371000 512888 371034
rect 512922 371000 512988 371034
rect 513022 371000 513088 371034
rect 513122 371000 513195 371034
rect 512501 370996 513195 371000
rect 512501 370962 512560 370996
rect 512594 370962 512650 370996
rect 512684 370962 512740 370996
rect 512774 370962 512830 370996
rect 512864 370962 512920 370996
rect 512954 370962 513010 370996
rect 513044 370962 513100 370996
rect 513134 370962 513195 370996
rect 512501 370934 513195 370962
rect 512501 370906 512588 370934
rect 512622 370906 512688 370934
rect 512501 370872 512560 370906
rect 512622 370900 512650 370906
rect 512594 370872 512650 370900
rect 512684 370900 512688 370906
rect 512722 370906 512788 370934
rect 512722 370900 512740 370906
rect 512684 370872 512740 370900
rect 512774 370900 512788 370906
rect 512822 370906 512888 370934
rect 512922 370906 512988 370934
rect 513022 370906 513088 370934
rect 513122 370906 513195 370934
rect 512822 370900 512830 370906
rect 512774 370872 512830 370900
rect 512864 370900 512888 370906
rect 512954 370900 512988 370906
rect 513044 370900 513088 370906
rect 512864 370872 512920 370900
rect 512954 370872 513010 370900
rect 513044 370872 513100 370900
rect 513134 370872 513195 370906
rect 512501 370813 513195 370872
rect 513257 371454 513329 371510
rect 513257 371420 513276 371454
rect 513310 371420 513329 371454
rect 513257 371364 513329 371420
rect 513257 371330 513276 371364
rect 513310 371330 513329 371364
rect 513257 371274 513329 371330
rect 513257 371240 513276 371274
rect 513310 371240 513329 371274
rect 513257 371184 513329 371240
rect 513257 371150 513276 371184
rect 513310 371150 513329 371184
rect 513257 371094 513329 371150
rect 513257 371060 513276 371094
rect 513310 371060 513329 371094
rect 513257 371004 513329 371060
rect 513257 370970 513276 371004
rect 513310 370970 513329 371004
rect 513257 370914 513329 370970
rect 513257 370880 513276 370914
rect 513310 370880 513329 370914
rect 513257 370824 513329 370880
rect 512367 370776 512384 370810
rect 512418 370790 512439 370810
rect 512367 370756 512386 370776
rect 512420 370756 512439 370790
rect 512367 370751 512439 370756
rect 513257 370790 513276 370824
rect 513310 370790 513329 370824
rect 513257 370751 513329 370790
rect 512367 370732 513329 370751
rect 512367 370720 512462 370732
rect 512367 370686 512384 370720
rect 512418 370698 512462 370720
rect 512496 370698 512552 370732
rect 512586 370698 512642 370732
rect 512676 370698 512732 370732
rect 512766 370698 512822 370732
rect 512856 370698 512912 370732
rect 512946 370698 513002 370732
rect 513036 370698 513092 370732
rect 513126 370698 513182 370732
rect 513216 370698 513329 370732
rect 512418 370686 513329 370698
rect 512367 370679 513329 370686
rect 513393 371640 513426 371674
rect 513460 371640 513492 371674
rect 513393 371584 513492 371640
rect 513393 371550 513426 371584
rect 513460 371550 513492 371584
rect 513393 371494 513492 371550
rect 513393 371460 513426 371494
rect 513460 371460 513492 371494
rect 513393 371404 513492 371460
rect 513393 371370 513426 371404
rect 513460 371370 513492 371404
rect 513393 371314 513492 371370
rect 513393 371280 513426 371314
rect 513460 371280 513492 371314
rect 513393 371224 513492 371280
rect 513393 371190 513426 371224
rect 513460 371190 513492 371224
rect 513393 371134 513492 371190
rect 513393 371100 513426 371134
rect 513460 371100 513492 371134
rect 513393 371044 513492 371100
rect 513393 371010 513426 371044
rect 513460 371010 513492 371044
rect 513393 370954 513492 371010
rect 513393 370920 513426 370954
rect 513460 370920 513492 370954
rect 513393 370864 513492 370920
rect 513393 370830 513426 370864
rect 513460 370830 513492 370864
rect 513393 370774 513492 370830
rect 513393 370740 513426 370774
rect 513460 370740 513492 370774
rect 513393 370684 513492 370740
rect 512204 370615 512303 370650
rect 513393 370650 513426 370684
rect 513460 370650 513492 370684
rect 513393 370615 513492 370650
rect 512204 370614 513492 370615
rect 512204 370580 512224 370614
rect 512258 370583 513492 370614
rect 512258 370580 512262 370583
rect 512204 370549 512262 370580
rect 512296 370549 512352 370583
rect 512386 370549 512442 370583
rect 512476 370549 512532 370583
rect 512566 370549 512622 370583
rect 512656 370549 512712 370583
rect 512746 370549 512802 370583
rect 512836 370549 512892 370583
rect 512926 370549 512982 370583
rect 513016 370549 513072 370583
rect 513106 370549 513162 370583
rect 513196 370549 513252 370583
rect 513286 370549 513342 370583
rect 513376 370549 513492 370583
rect 512204 370444 513492 370549
rect 512204 370410 512224 370444
rect 512258 370430 513492 370444
rect 512258 370410 512262 370430
rect 512204 370396 512262 370410
rect 512296 370396 512352 370430
rect 512386 370396 512442 370430
rect 512476 370396 512532 370430
rect 512566 370396 512622 370430
rect 512656 370396 512712 370430
rect 512746 370396 512802 370430
rect 512836 370396 512892 370430
rect 512926 370396 512982 370430
rect 513016 370396 513072 370430
rect 513106 370396 513162 370430
rect 513196 370396 513252 370430
rect 513286 370396 513342 370430
rect 513376 370396 513492 370430
rect 512204 370365 513492 370396
rect 512204 370354 512303 370365
rect 512204 370320 512224 370354
rect 512258 370334 512303 370354
rect 512204 370300 512239 370320
rect 512273 370300 512303 370334
rect 513393 370334 513492 370365
rect 512204 370264 512303 370300
rect 512204 370230 512224 370264
rect 512258 370244 512303 370264
rect 512204 370210 512239 370230
rect 512273 370210 512303 370244
rect 512204 370174 512303 370210
rect 512204 370140 512224 370174
rect 512258 370154 512303 370174
rect 512204 370120 512239 370140
rect 512273 370120 512303 370154
rect 512204 370084 512303 370120
rect 512204 370050 512224 370084
rect 512258 370064 512303 370084
rect 512204 370030 512239 370050
rect 512273 370030 512303 370064
rect 512204 369994 512303 370030
rect 512204 369960 512224 369994
rect 512258 369974 512303 369994
rect 512204 369940 512239 369960
rect 512273 369940 512303 369974
rect 512204 369904 512303 369940
rect 512204 369870 512224 369904
rect 512258 369884 512303 369904
rect 512204 369850 512239 369870
rect 512273 369850 512303 369884
rect 512204 369814 512303 369850
rect 512204 369780 512224 369814
rect 512258 369794 512303 369814
rect 512204 369760 512239 369780
rect 512273 369760 512303 369794
rect 512204 369724 512303 369760
rect 512204 369690 512224 369724
rect 512258 369704 512303 369724
rect 512204 369670 512239 369690
rect 512273 369670 512303 369704
rect 512204 369634 512303 369670
rect 512204 369600 512224 369634
rect 512258 369614 512303 369634
rect 512204 369580 512239 369600
rect 512273 369580 512303 369614
rect 512204 369544 512303 369580
rect 512204 369510 512224 369544
rect 512258 369524 512303 369544
rect 512204 369490 512239 369510
rect 512273 369490 512303 369524
rect 512204 369454 512303 369490
rect 512204 369420 512224 369454
rect 512258 369434 512303 369454
rect 512204 369400 512239 369420
rect 512273 369400 512303 369434
rect 512204 369364 512303 369400
rect 512204 369330 512224 369364
rect 512258 369344 512303 369364
rect 512204 369310 512239 369330
rect 512273 369310 512303 369344
rect 512367 370282 513329 370301
rect 512367 370280 512443 370282
rect 512367 370246 512384 370280
rect 512418 370248 512443 370280
rect 512477 370248 512533 370282
rect 512567 370248 512623 370282
rect 512657 370248 512713 370282
rect 512747 370248 512803 370282
rect 512837 370248 512893 370282
rect 512927 370248 512983 370282
rect 513017 370248 513073 370282
rect 513107 370248 513163 370282
rect 513197 370248 513329 370282
rect 512418 370246 513329 370248
rect 512367 370229 513329 370246
rect 512367 370190 512439 370229
rect 512367 370156 512384 370190
rect 512418 370170 512439 370190
rect 512367 370136 512386 370156
rect 512420 370136 512439 370170
rect 513257 370204 513329 370229
rect 513257 370170 513276 370204
rect 513310 370170 513329 370204
rect 512367 370100 512439 370136
rect 512367 370066 512384 370100
rect 512418 370080 512439 370100
rect 512367 370046 512386 370066
rect 512420 370046 512439 370080
rect 512367 370010 512439 370046
rect 512367 369976 512384 370010
rect 512418 369990 512439 370010
rect 512367 369956 512386 369976
rect 512420 369956 512439 369990
rect 512367 369920 512439 369956
rect 512367 369886 512384 369920
rect 512418 369900 512439 369920
rect 512367 369866 512386 369886
rect 512420 369866 512439 369900
rect 512367 369830 512439 369866
rect 512367 369796 512384 369830
rect 512418 369810 512439 369830
rect 512367 369776 512386 369796
rect 512420 369776 512439 369810
rect 512367 369740 512439 369776
rect 512367 369706 512384 369740
rect 512418 369720 512439 369740
rect 512367 369686 512386 369706
rect 512420 369686 512439 369720
rect 512367 369650 512439 369686
rect 512367 369616 512384 369650
rect 512418 369630 512439 369650
rect 512367 369596 512386 369616
rect 512420 369596 512439 369630
rect 512367 369560 512439 369596
rect 512367 369526 512384 369560
rect 512418 369540 512439 369560
rect 512367 369506 512386 369526
rect 512420 369506 512439 369540
rect 512367 369470 512439 369506
rect 512501 370106 513195 370167
rect 512501 370072 512560 370106
rect 512594 370094 512650 370106
rect 512622 370072 512650 370094
rect 512684 370094 512740 370106
rect 512684 370072 512688 370094
rect 512501 370060 512588 370072
rect 512622 370060 512688 370072
rect 512722 370072 512740 370094
rect 512774 370094 512830 370106
rect 512774 370072 512788 370094
rect 512722 370060 512788 370072
rect 512822 370072 512830 370094
rect 512864 370094 512920 370106
rect 512954 370094 513010 370106
rect 513044 370094 513100 370106
rect 512864 370072 512888 370094
rect 512954 370072 512988 370094
rect 513044 370072 513088 370094
rect 513134 370072 513195 370106
rect 512822 370060 512888 370072
rect 512922 370060 512988 370072
rect 513022 370060 513088 370072
rect 513122 370060 513195 370072
rect 512501 370016 513195 370060
rect 512501 369982 512560 370016
rect 512594 369994 512650 370016
rect 512622 369982 512650 369994
rect 512684 369994 512740 370016
rect 512684 369982 512688 369994
rect 512501 369960 512588 369982
rect 512622 369960 512688 369982
rect 512722 369982 512740 369994
rect 512774 369994 512830 370016
rect 512774 369982 512788 369994
rect 512722 369960 512788 369982
rect 512822 369982 512830 369994
rect 512864 369994 512920 370016
rect 512954 369994 513010 370016
rect 513044 369994 513100 370016
rect 512864 369982 512888 369994
rect 512954 369982 512988 369994
rect 513044 369982 513088 369994
rect 513134 369982 513195 370016
rect 512822 369960 512888 369982
rect 512922 369960 512988 369982
rect 513022 369960 513088 369982
rect 513122 369960 513195 369982
rect 512501 369926 513195 369960
rect 512501 369892 512560 369926
rect 512594 369894 512650 369926
rect 512622 369892 512650 369894
rect 512684 369894 512740 369926
rect 512684 369892 512688 369894
rect 512501 369860 512588 369892
rect 512622 369860 512688 369892
rect 512722 369892 512740 369894
rect 512774 369894 512830 369926
rect 512774 369892 512788 369894
rect 512722 369860 512788 369892
rect 512822 369892 512830 369894
rect 512864 369894 512920 369926
rect 512954 369894 513010 369926
rect 513044 369894 513100 369926
rect 512864 369892 512888 369894
rect 512954 369892 512988 369894
rect 513044 369892 513088 369894
rect 513134 369892 513195 369926
rect 512822 369860 512888 369892
rect 512922 369860 512988 369892
rect 513022 369860 513088 369892
rect 513122 369860 513195 369892
rect 512501 369836 513195 369860
rect 512501 369802 512560 369836
rect 512594 369802 512650 369836
rect 512684 369802 512740 369836
rect 512774 369802 512830 369836
rect 512864 369802 512920 369836
rect 512954 369802 513010 369836
rect 513044 369802 513100 369836
rect 513134 369802 513195 369836
rect 512501 369794 513195 369802
rect 512501 369760 512588 369794
rect 512622 369760 512688 369794
rect 512722 369760 512788 369794
rect 512822 369760 512888 369794
rect 512922 369760 512988 369794
rect 513022 369760 513088 369794
rect 513122 369760 513195 369794
rect 512501 369746 513195 369760
rect 512501 369712 512560 369746
rect 512594 369712 512650 369746
rect 512684 369712 512740 369746
rect 512774 369712 512830 369746
rect 512864 369712 512920 369746
rect 512954 369712 513010 369746
rect 513044 369712 513100 369746
rect 513134 369712 513195 369746
rect 512501 369694 513195 369712
rect 512501 369660 512588 369694
rect 512622 369660 512688 369694
rect 512722 369660 512788 369694
rect 512822 369660 512888 369694
rect 512922 369660 512988 369694
rect 513022 369660 513088 369694
rect 513122 369660 513195 369694
rect 512501 369656 513195 369660
rect 512501 369622 512560 369656
rect 512594 369622 512650 369656
rect 512684 369622 512740 369656
rect 512774 369622 512830 369656
rect 512864 369622 512920 369656
rect 512954 369622 513010 369656
rect 513044 369622 513100 369656
rect 513134 369622 513195 369656
rect 512501 369594 513195 369622
rect 512501 369566 512588 369594
rect 512622 369566 512688 369594
rect 512501 369532 512560 369566
rect 512622 369560 512650 369566
rect 512594 369532 512650 369560
rect 512684 369560 512688 369566
rect 512722 369566 512788 369594
rect 512722 369560 512740 369566
rect 512684 369532 512740 369560
rect 512774 369560 512788 369566
rect 512822 369566 512888 369594
rect 512922 369566 512988 369594
rect 513022 369566 513088 369594
rect 513122 369566 513195 369594
rect 512822 369560 512830 369566
rect 512774 369532 512830 369560
rect 512864 369560 512888 369566
rect 512954 369560 512988 369566
rect 513044 369560 513088 369566
rect 512864 369532 512920 369560
rect 512954 369532 513010 369560
rect 513044 369532 513100 369560
rect 513134 369532 513195 369566
rect 512501 369473 513195 369532
rect 513257 370114 513329 370170
rect 513257 370080 513276 370114
rect 513310 370080 513329 370114
rect 513257 370024 513329 370080
rect 513257 369990 513276 370024
rect 513310 369990 513329 370024
rect 513257 369934 513329 369990
rect 513257 369900 513276 369934
rect 513310 369900 513329 369934
rect 513257 369844 513329 369900
rect 513257 369810 513276 369844
rect 513310 369810 513329 369844
rect 513257 369754 513329 369810
rect 513257 369720 513276 369754
rect 513310 369720 513329 369754
rect 513257 369664 513329 369720
rect 513257 369630 513276 369664
rect 513310 369630 513329 369664
rect 513257 369574 513329 369630
rect 513257 369540 513276 369574
rect 513310 369540 513329 369574
rect 513257 369484 513329 369540
rect 512367 369436 512384 369470
rect 512418 369450 512439 369470
rect 512367 369416 512386 369436
rect 512420 369416 512439 369450
rect 512367 369411 512439 369416
rect 513257 369450 513276 369484
rect 513310 369450 513329 369484
rect 513257 369411 513329 369450
rect 512367 369392 513329 369411
rect 512367 369380 512462 369392
rect 512367 369346 512384 369380
rect 512418 369358 512462 369380
rect 512496 369358 512552 369392
rect 512586 369358 512642 369392
rect 512676 369358 512732 369392
rect 512766 369358 512822 369392
rect 512856 369358 512912 369392
rect 512946 369358 513002 369392
rect 513036 369358 513092 369392
rect 513126 369358 513182 369392
rect 513216 369358 513329 369392
rect 512418 369346 513329 369358
rect 512367 369339 513329 369346
rect 513393 370300 513426 370334
rect 513460 370300 513492 370334
rect 513393 370244 513492 370300
rect 513393 370210 513426 370244
rect 513460 370210 513492 370244
rect 513393 370154 513492 370210
rect 513393 370120 513426 370154
rect 513460 370120 513492 370154
rect 513393 370064 513492 370120
rect 513393 370030 513426 370064
rect 513460 370030 513492 370064
rect 513393 369974 513492 370030
rect 513393 369940 513426 369974
rect 513460 369940 513492 369974
rect 513393 369884 513492 369940
rect 513393 369850 513426 369884
rect 513460 369850 513492 369884
rect 513393 369794 513492 369850
rect 513393 369760 513426 369794
rect 513460 369760 513492 369794
rect 513393 369704 513492 369760
rect 513393 369670 513426 369704
rect 513460 369670 513492 369704
rect 513393 369614 513492 369670
rect 513393 369580 513426 369614
rect 513460 369580 513492 369614
rect 513393 369524 513492 369580
rect 513393 369490 513426 369524
rect 513460 369490 513492 369524
rect 513393 369434 513492 369490
rect 513393 369400 513426 369434
rect 513460 369400 513492 369434
rect 513393 369344 513492 369400
rect 512204 369275 512303 369310
rect 513393 369310 513426 369344
rect 513460 369310 513492 369344
rect 513393 369275 513492 369310
rect 512204 369274 513492 369275
rect 512204 369240 512224 369274
rect 512258 369243 513492 369274
rect 512258 369240 512262 369243
rect 512204 369209 512262 369240
rect 512296 369209 512352 369243
rect 512386 369209 512442 369243
rect 512476 369209 512532 369243
rect 512566 369209 512622 369243
rect 512656 369209 512712 369243
rect 512746 369209 512802 369243
rect 512836 369209 512892 369243
rect 512926 369209 512982 369243
rect 513016 369209 513072 369243
rect 513106 369209 513162 369243
rect 513196 369209 513252 369243
rect 513286 369209 513342 369243
rect 513376 369209 513492 369243
rect 512204 369104 513492 369209
rect 512204 369070 512224 369104
rect 512258 369090 513492 369104
rect 512258 369070 512262 369090
rect 512204 369056 512262 369070
rect 512296 369056 512352 369090
rect 512386 369056 512442 369090
rect 512476 369056 512532 369090
rect 512566 369056 512622 369090
rect 512656 369056 512712 369090
rect 512746 369056 512802 369090
rect 512836 369056 512892 369090
rect 512926 369056 512982 369090
rect 513016 369056 513072 369090
rect 513106 369056 513162 369090
rect 513196 369056 513252 369090
rect 513286 369056 513342 369090
rect 513376 369056 513492 369090
rect 512204 369025 513492 369056
rect 512204 369014 512303 369025
rect 512204 368980 512224 369014
rect 512258 368994 512303 369014
rect 512204 368960 512239 368980
rect 512273 368960 512303 368994
rect 513393 368994 513492 369025
rect 512204 368924 512303 368960
rect 512204 368890 512224 368924
rect 512258 368904 512303 368924
rect 512204 368870 512239 368890
rect 512273 368870 512303 368904
rect 512204 368834 512303 368870
rect 512204 368800 512224 368834
rect 512258 368814 512303 368834
rect 512204 368780 512239 368800
rect 512273 368780 512303 368814
rect 512204 368744 512303 368780
rect 512204 368710 512224 368744
rect 512258 368724 512303 368744
rect 512204 368690 512239 368710
rect 512273 368690 512303 368724
rect 512204 368654 512303 368690
rect 512204 368620 512224 368654
rect 512258 368634 512303 368654
rect 512204 368600 512239 368620
rect 512273 368600 512303 368634
rect 512204 368564 512303 368600
rect 512204 368530 512224 368564
rect 512258 368544 512303 368564
rect 512204 368510 512239 368530
rect 512273 368510 512303 368544
rect 512204 368474 512303 368510
rect 512204 368440 512224 368474
rect 512258 368454 512303 368474
rect 512204 368420 512239 368440
rect 512273 368420 512303 368454
rect 512204 368384 512303 368420
rect 512204 368350 512224 368384
rect 512258 368364 512303 368384
rect 512204 368330 512239 368350
rect 512273 368330 512303 368364
rect 512204 368294 512303 368330
rect 512204 368260 512224 368294
rect 512258 368274 512303 368294
rect 512204 368240 512239 368260
rect 512273 368240 512303 368274
rect 512204 368204 512303 368240
rect 512204 368170 512224 368204
rect 512258 368184 512303 368204
rect 512204 368150 512239 368170
rect 512273 368150 512303 368184
rect 512204 368114 512303 368150
rect 512204 368080 512224 368114
rect 512258 368094 512303 368114
rect 512204 368060 512239 368080
rect 512273 368060 512303 368094
rect 512204 368024 512303 368060
rect 512204 367990 512224 368024
rect 512258 368004 512303 368024
rect 512204 367970 512239 367990
rect 512273 367970 512303 368004
rect 512367 368942 513329 368961
rect 512367 368940 512443 368942
rect 512367 368906 512384 368940
rect 512418 368908 512443 368940
rect 512477 368908 512533 368942
rect 512567 368908 512623 368942
rect 512657 368908 512713 368942
rect 512747 368908 512803 368942
rect 512837 368908 512893 368942
rect 512927 368908 512983 368942
rect 513017 368908 513073 368942
rect 513107 368908 513163 368942
rect 513197 368908 513329 368942
rect 512418 368906 513329 368908
rect 512367 368889 513329 368906
rect 512367 368850 512439 368889
rect 512367 368816 512384 368850
rect 512418 368830 512439 368850
rect 512367 368796 512386 368816
rect 512420 368796 512439 368830
rect 513257 368864 513329 368889
rect 513257 368830 513276 368864
rect 513310 368830 513329 368864
rect 512367 368760 512439 368796
rect 512367 368726 512384 368760
rect 512418 368740 512439 368760
rect 512367 368706 512386 368726
rect 512420 368706 512439 368740
rect 512367 368670 512439 368706
rect 512367 368636 512384 368670
rect 512418 368650 512439 368670
rect 512367 368616 512386 368636
rect 512420 368616 512439 368650
rect 512367 368580 512439 368616
rect 512367 368546 512384 368580
rect 512418 368560 512439 368580
rect 512367 368526 512386 368546
rect 512420 368526 512439 368560
rect 512367 368490 512439 368526
rect 512367 368456 512384 368490
rect 512418 368470 512439 368490
rect 512367 368436 512386 368456
rect 512420 368436 512439 368470
rect 512367 368400 512439 368436
rect 512367 368366 512384 368400
rect 512418 368380 512439 368400
rect 512367 368346 512386 368366
rect 512420 368346 512439 368380
rect 512367 368310 512439 368346
rect 512367 368276 512384 368310
rect 512418 368290 512439 368310
rect 512367 368256 512386 368276
rect 512420 368256 512439 368290
rect 512367 368220 512439 368256
rect 512367 368186 512384 368220
rect 512418 368200 512439 368220
rect 512367 368166 512386 368186
rect 512420 368166 512439 368200
rect 512367 368130 512439 368166
rect 512501 368766 513195 368827
rect 512501 368732 512560 368766
rect 512594 368754 512650 368766
rect 512622 368732 512650 368754
rect 512684 368754 512740 368766
rect 512684 368732 512688 368754
rect 512501 368720 512588 368732
rect 512622 368720 512688 368732
rect 512722 368732 512740 368754
rect 512774 368754 512830 368766
rect 512774 368732 512788 368754
rect 512722 368720 512788 368732
rect 512822 368732 512830 368754
rect 512864 368754 512920 368766
rect 512954 368754 513010 368766
rect 513044 368754 513100 368766
rect 512864 368732 512888 368754
rect 512954 368732 512988 368754
rect 513044 368732 513088 368754
rect 513134 368732 513195 368766
rect 512822 368720 512888 368732
rect 512922 368720 512988 368732
rect 513022 368720 513088 368732
rect 513122 368720 513195 368732
rect 512501 368676 513195 368720
rect 512501 368642 512560 368676
rect 512594 368654 512650 368676
rect 512622 368642 512650 368654
rect 512684 368654 512740 368676
rect 512684 368642 512688 368654
rect 512501 368620 512588 368642
rect 512622 368620 512688 368642
rect 512722 368642 512740 368654
rect 512774 368654 512830 368676
rect 512774 368642 512788 368654
rect 512722 368620 512788 368642
rect 512822 368642 512830 368654
rect 512864 368654 512920 368676
rect 512954 368654 513010 368676
rect 513044 368654 513100 368676
rect 512864 368642 512888 368654
rect 512954 368642 512988 368654
rect 513044 368642 513088 368654
rect 513134 368642 513195 368676
rect 512822 368620 512888 368642
rect 512922 368620 512988 368642
rect 513022 368620 513088 368642
rect 513122 368620 513195 368642
rect 512501 368586 513195 368620
rect 512501 368552 512560 368586
rect 512594 368554 512650 368586
rect 512622 368552 512650 368554
rect 512684 368554 512740 368586
rect 512684 368552 512688 368554
rect 512501 368520 512588 368552
rect 512622 368520 512688 368552
rect 512722 368552 512740 368554
rect 512774 368554 512830 368586
rect 512774 368552 512788 368554
rect 512722 368520 512788 368552
rect 512822 368552 512830 368554
rect 512864 368554 512920 368586
rect 512954 368554 513010 368586
rect 513044 368554 513100 368586
rect 512864 368552 512888 368554
rect 512954 368552 512988 368554
rect 513044 368552 513088 368554
rect 513134 368552 513195 368586
rect 512822 368520 512888 368552
rect 512922 368520 512988 368552
rect 513022 368520 513088 368552
rect 513122 368520 513195 368552
rect 512501 368496 513195 368520
rect 512501 368462 512560 368496
rect 512594 368462 512650 368496
rect 512684 368462 512740 368496
rect 512774 368462 512830 368496
rect 512864 368462 512920 368496
rect 512954 368462 513010 368496
rect 513044 368462 513100 368496
rect 513134 368462 513195 368496
rect 512501 368454 513195 368462
rect 512501 368420 512588 368454
rect 512622 368420 512688 368454
rect 512722 368420 512788 368454
rect 512822 368420 512888 368454
rect 512922 368420 512988 368454
rect 513022 368420 513088 368454
rect 513122 368420 513195 368454
rect 512501 368406 513195 368420
rect 512501 368372 512560 368406
rect 512594 368372 512650 368406
rect 512684 368372 512740 368406
rect 512774 368372 512830 368406
rect 512864 368372 512920 368406
rect 512954 368372 513010 368406
rect 513044 368372 513100 368406
rect 513134 368372 513195 368406
rect 512501 368354 513195 368372
rect 512501 368320 512588 368354
rect 512622 368320 512688 368354
rect 512722 368320 512788 368354
rect 512822 368320 512888 368354
rect 512922 368320 512988 368354
rect 513022 368320 513088 368354
rect 513122 368320 513195 368354
rect 512501 368316 513195 368320
rect 512501 368282 512560 368316
rect 512594 368282 512650 368316
rect 512684 368282 512740 368316
rect 512774 368282 512830 368316
rect 512864 368282 512920 368316
rect 512954 368282 513010 368316
rect 513044 368282 513100 368316
rect 513134 368282 513195 368316
rect 512501 368254 513195 368282
rect 512501 368226 512588 368254
rect 512622 368226 512688 368254
rect 512501 368192 512560 368226
rect 512622 368220 512650 368226
rect 512594 368192 512650 368220
rect 512684 368220 512688 368226
rect 512722 368226 512788 368254
rect 512722 368220 512740 368226
rect 512684 368192 512740 368220
rect 512774 368220 512788 368226
rect 512822 368226 512888 368254
rect 512922 368226 512988 368254
rect 513022 368226 513088 368254
rect 513122 368226 513195 368254
rect 512822 368220 512830 368226
rect 512774 368192 512830 368220
rect 512864 368220 512888 368226
rect 512954 368220 512988 368226
rect 513044 368220 513088 368226
rect 512864 368192 512920 368220
rect 512954 368192 513010 368220
rect 513044 368192 513100 368220
rect 513134 368192 513195 368226
rect 512501 368133 513195 368192
rect 513257 368774 513329 368830
rect 513257 368740 513276 368774
rect 513310 368740 513329 368774
rect 513257 368684 513329 368740
rect 513257 368650 513276 368684
rect 513310 368650 513329 368684
rect 513257 368594 513329 368650
rect 513257 368560 513276 368594
rect 513310 368560 513329 368594
rect 513257 368504 513329 368560
rect 513257 368470 513276 368504
rect 513310 368470 513329 368504
rect 513257 368414 513329 368470
rect 513257 368380 513276 368414
rect 513310 368380 513329 368414
rect 513257 368324 513329 368380
rect 513257 368290 513276 368324
rect 513310 368290 513329 368324
rect 513257 368234 513329 368290
rect 513257 368200 513276 368234
rect 513310 368200 513329 368234
rect 513257 368144 513329 368200
rect 512367 368096 512384 368130
rect 512418 368110 512439 368130
rect 512367 368076 512386 368096
rect 512420 368076 512439 368110
rect 512367 368071 512439 368076
rect 513257 368110 513276 368144
rect 513310 368110 513329 368144
rect 513257 368071 513329 368110
rect 512367 368052 513329 368071
rect 512367 368040 512462 368052
rect 512367 368006 512384 368040
rect 512418 368018 512462 368040
rect 512496 368018 512552 368052
rect 512586 368018 512642 368052
rect 512676 368018 512732 368052
rect 512766 368018 512822 368052
rect 512856 368018 512912 368052
rect 512946 368018 513002 368052
rect 513036 368018 513092 368052
rect 513126 368018 513182 368052
rect 513216 368018 513329 368052
rect 512418 368006 513329 368018
rect 512367 367999 513329 368006
rect 513393 368960 513426 368994
rect 513460 368960 513492 368994
rect 513393 368904 513492 368960
rect 513393 368870 513426 368904
rect 513460 368870 513492 368904
rect 513393 368814 513492 368870
rect 513393 368780 513426 368814
rect 513460 368780 513492 368814
rect 513393 368724 513492 368780
rect 513393 368690 513426 368724
rect 513460 368690 513492 368724
rect 513393 368634 513492 368690
rect 513393 368600 513426 368634
rect 513460 368600 513492 368634
rect 513393 368544 513492 368600
rect 513393 368510 513426 368544
rect 513460 368510 513492 368544
rect 513393 368454 513492 368510
rect 513393 368420 513426 368454
rect 513460 368420 513492 368454
rect 513393 368364 513492 368420
rect 513393 368330 513426 368364
rect 513460 368330 513492 368364
rect 513393 368274 513492 368330
rect 513393 368240 513426 368274
rect 513460 368240 513492 368274
rect 513393 368184 513492 368240
rect 513393 368150 513426 368184
rect 513460 368150 513492 368184
rect 513393 368094 513492 368150
rect 513393 368060 513426 368094
rect 513460 368060 513492 368094
rect 513393 368004 513492 368060
rect 512204 367935 512303 367970
rect 513393 367970 513426 368004
rect 513460 367970 513492 368004
rect 513393 367935 513492 367970
rect 512204 367934 513492 367935
rect 512204 367900 512224 367934
rect 512258 367903 513492 367934
rect 512258 367900 512262 367903
rect 512204 367869 512262 367900
rect 512296 367869 512352 367903
rect 512386 367869 512442 367903
rect 512476 367869 512532 367903
rect 512566 367869 512622 367903
rect 512656 367869 512712 367903
rect 512746 367869 512802 367903
rect 512836 367869 512892 367903
rect 512926 367869 512982 367903
rect 513016 367869 513072 367903
rect 513106 367869 513162 367903
rect 513196 367869 513252 367903
rect 513286 367869 513342 367903
rect 513376 367869 513492 367903
rect 512204 367764 513492 367869
rect 512204 367730 512224 367764
rect 512258 367750 513492 367764
rect 512258 367730 512262 367750
rect 512204 367716 512262 367730
rect 512296 367716 512352 367750
rect 512386 367716 512442 367750
rect 512476 367716 512532 367750
rect 512566 367716 512622 367750
rect 512656 367716 512712 367750
rect 512746 367716 512802 367750
rect 512836 367716 512892 367750
rect 512926 367716 512982 367750
rect 513016 367716 513072 367750
rect 513106 367716 513162 367750
rect 513196 367716 513252 367750
rect 513286 367716 513342 367750
rect 513376 367716 513492 367750
rect 512204 367685 513492 367716
rect 512204 367674 512303 367685
rect 512204 367640 512224 367674
rect 512258 367654 512303 367674
rect 512204 367620 512239 367640
rect 512273 367620 512303 367654
rect 513393 367654 513492 367685
rect 512204 367584 512303 367620
rect 512204 367550 512224 367584
rect 512258 367564 512303 367584
rect 512204 367530 512239 367550
rect 512273 367530 512303 367564
rect 512204 367494 512303 367530
rect 512204 367460 512224 367494
rect 512258 367474 512303 367494
rect 512204 367440 512239 367460
rect 512273 367440 512303 367474
rect 512204 367404 512303 367440
rect 512204 367370 512224 367404
rect 512258 367384 512303 367404
rect 512204 367350 512239 367370
rect 512273 367350 512303 367384
rect 512204 367314 512303 367350
rect 512204 367280 512224 367314
rect 512258 367294 512303 367314
rect 512204 367260 512239 367280
rect 512273 367260 512303 367294
rect 512204 367224 512303 367260
rect 512204 367190 512224 367224
rect 512258 367204 512303 367224
rect 512204 367170 512239 367190
rect 512273 367170 512303 367204
rect 512204 367134 512303 367170
rect 512204 367100 512224 367134
rect 512258 367114 512303 367134
rect 512204 367080 512239 367100
rect 512273 367080 512303 367114
rect 512204 367044 512303 367080
rect 512204 367010 512224 367044
rect 512258 367024 512303 367044
rect 512204 366990 512239 367010
rect 512273 366990 512303 367024
rect 512204 366954 512303 366990
rect 512204 366920 512224 366954
rect 512258 366934 512303 366954
rect 512204 366900 512239 366920
rect 512273 366900 512303 366934
rect 512204 366864 512303 366900
rect 512204 366830 512224 366864
rect 512258 366844 512303 366864
rect 512204 366810 512239 366830
rect 512273 366810 512303 366844
rect 512204 366774 512303 366810
rect 512204 366740 512224 366774
rect 512258 366754 512303 366774
rect 512204 366720 512239 366740
rect 512273 366720 512303 366754
rect 512204 366684 512303 366720
rect 512204 366650 512224 366684
rect 512258 366664 512303 366684
rect 512204 366630 512239 366650
rect 512273 366630 512303 366664
rect 512367 367602 513329 367621
rect 512367 367600 512443 367602
rect 512367 367566 512384 367600
rect 512418 367568 512443 367600
rect 512477 367568 512533 367602
rect 512567 367568 512623 367602
rect 512657 367568 512713 367602
rect 512747 367568 512803 367602
rect 512837 367568 512893 367602
rect 512927 367568 512983 367602
rect 513017 367568 513073 367602
rect 513107 367568 513163 367602
rect 513197 367568 513329 367602
rect 512418 367566 513329 367568
rect 512367 367549 513329 367566
rect 512367 367510 512439 367549
rect 512367 367476 512384 367510
rect 512418 367490 512439 367510
rect 512367 367456 512386 367476
rect 512420 367456 512439 367490
rect 513257 367524 513329 367549
rect 513257 367490 513276 367524
rect 513310 367490 513329 367524
rect 512367 367420 512439 367456
rect 512367 367386 512384 367420
rect 512418 367400 512439 367420
rect 512367 367366 512386 367386
rect 512420 367366 512439 367400
rect 512367 367330 512439 367366
rect 512367 367296 512384 367330
rect 512418 367310 512439 367330
rect 512367 367276 512386 367296
rect 512420 367276 512439 367310
rect 512367 367240 512439 367276
rect 512367 367206 512384 367240
rect 512418 367220 512439 367240
rect 512367 367186 512386 367206
rect 512420 367186 512439 367220
rect 512367 367150 512439 367186
rect 512367 367116 512384 367150
rect 512418 367130 512439 367150
rect 512367 367096 512386 367116
rect 512420 367096 512439 367130
rect 512367 367060 512439 367096
rect 512367 367026 512384 367060
rect 512418 367040 512439 367060
rect 512367 367006 512386 367026
rect 512420 367006 512439 367040
rect 512367 366970 512439 367006
rect 512367 366936 512384 366970
rect 512418 366950 512439 366970
rect 512367 366916 512386 366936
rect 512420 366916 512439 366950
rect 512367 366880 512439 366916
rect 512367 366846 512384 366880
rect 512418 366860 512439 366880
rect 512367 366826 512386 366846
rect 512420 366826 512439 366860
rect 512367 366790 512439 366826
rect 512501 367426 513195 367487
rect 512501 367392 512560 367426
rect 512594 367414 512650 367426
rect 512622 367392 512650 367414
rect 512684 367414 512740 367426
rect 512684 367392 512688 367414
rect 512501 367380 512588 367392
rect 512622 367380 512688 367392
rect 512722 367392 512740 367414
rect 512774 367414 512830 367426
rect 512774 367392 512788 367414
rect 512722 367380 512788 367392
rect 512822 367392 512830 367414
rect 512864 367414 512920 367426
rect 512954 367414 513010 367426
rect 513044 367414 513100 367426
rect 512864 367392 512888 367414
rect 512954 367392 512988 367414
rect 513044 367392 513088 367414
rect 513134 367392 513195 367426
rect 512822 367380 512888 367392
rect 512922 367380 512988 367392
rect 513022 367380 513088 367392
rect 513122 367380 513195 367392
rect 512501 367336 513195 367380
rect 512501 367302 512560 367336
rect 512594 367314 512650 367336
rect 512622 367302 512650 367314
rect 512684 367314 512740 367336
rect 512684 367302 512688 367314
rect 512501 367280 512588 367302
rect 512622 367280 512688 367302
rect 512722 367302 512740 367314
rect 512774 367314 512830 367336
rect 512774 367302 512788 367314
rect 512722 367280 512788 367302
rect 512822 367302 512830 367314
rect 512864 367314 512920 367336
rect 512954 367314 513010 367336
rect 513044 367314 513100 367336
rect 512864 367302 512888 367314
rect 512954 367302 512988 367314
rect 513044 367302 513088 367314
rect 513134 367302 513195 367336
rect 512822 367280 512888 367302
rect 512922 367280 512988 367302
rect 513022 367280 513088 367302
rect 513122 367280 513195 367302
rect 512501 367246 513195 367280
rect 512501 367212 512560 367246
rect 512594 367214 512650 367246
rect 512622 367212 512650 367214
rect 512684 367214 512740 367246
rect 512684 367212 512688 367214
rect 512501 367180 512588 367212
rect 512622 367180 512688 367212
rect 512722 367212 512740 367214
rect 512774 367214 512830 367246
rect 512774 367212 512788 367214
rect 512722 367180 512788 367212
rect 512822 367212 512830 367214
rect 512864 367214 512920 367246
rect 512954 367214 513010 367246
rect 513044 367214 513100 367246
rect 512864 367212 512888 367214
rect 512954 367212 512988 367214
rect 513044 367212 513088 367214
rect 513134 367212 513195 367246
rect 512822 367180 512888 367212
rect 512922 367180 512988 367212
rect 513022 367180 513088 367212
rect 513122 367180 513195 367212
rect 512501 367156 513195 367180
rect 512501 367122 512560 367156
rect 512594 367122 512650 367156
rect 512684 367122 512740 367156
rect 512774 367122 512830 367156
rect 512864 367122 512920 367156
rect 512954 367122 513010 367156
rect 513044 367122 513100 367156
rect 513134 367122 513195 367156
rect 512501 367114 513195 367122
rect 512501 367080 512588 367114
rect 512622 367080 512688 367114
rect 512722 367080 512788 367114
rect 512822 367080 512888 367114
rect 512922 367080 512988 367114
rect 513022 367080 513088 367114
rect 513122 367080 513195 367114
rect 512501 367066 513195 367080
rect 512501 367032 512560 367066
rect 512594 367032 512650 367066
rect 512684 367032 512740 367066
rect 512774 367032 512830 367066
rect 512864 367032 512920 367066
rect 512954 367032 513010 367066
rect 513044 367032 513100 367066
rect 513134 367032 513195 367066
rect 512501 367014 513195 367032
rect 512501 366980 512588 367014
rect 512622 366980 512688 367014
rect 512722 366980 512788 367014
rect 512822 366980 512888 367014
rect 512922 366980 512988 367014
rect 513022 366980 513088 367014
rect 513122 366980 513195 367014
rect 512501 366976 513195 366980
rect 512501 366942 512560 366976
rect 512594 366942 512650 366976
rect 512684 366942 512740 366976
rect 512774 366942 512830 366976
rect 512864 366942 512920 366976
rect 512954 366942 513010 366976
rect 513044 366942 513100 366976
rect 513134 366942 513195 366976
rect 512501 366914 513195 366942
rect 512501 366886 512588 366914
rect 512622 366886 512688 366914
rect 512501 366852 512560 366886
rect 512622 366880 512650 366886
rect 512594 366852 512650 366880
rect 512684 366880 512688 366886
rect 512722 366886 512788 366914
rect 512722 366880 512740 366886
rect 512684 366852 512740 366880
rect 512774 366880 512788 366886
rect 512822 366886 512888 366914
rect 512922 366886 512988 366914
rect 513022 366886 513088 366914
rect 513122 366886 513195 366914
rect 512822 366880 512830 366886
rect 512774 366852 512830 366880
rect 512864 366880 512888 366886
rect 512954 366880 512988 366886
rect 513044 366880 513088 366886
rect 512864 366852 512920 366880
rect 512954 366852 513010 366880
rect 513044 366852 513100 366880
rect 513134 366852 513195 366886
rect 512501 366793 513195 366852
rect 513257 367434 513329 367490
rect 513257 367400 513276 367434
rect 513310 367400 513329 367434
rect 513257 367344 513329 367400
rect 513257 367310 513276 367344
rect 513310 367310 513329 367344
rect 513257 367254 513329 367310
rect 513257 367220 513276 367254
rect 513310 367220 513329 367254
rect 513257 367164 513329 367220
rect 513257 367130 513276 367164
rect 513310 367130 513329 367164
rect 513257 367074 513329 367130
rect 513257 367040 513276 367074
rect 513310 367040 513329 367074
rect 513257 366984 513329 367040
rect 513257 366950 513276 366984
rect 513310 366950 513329 366984
rect 513257 366894 513329 366950
rect 513257 366860 513276 366894
rect 513310 366860 513329 366894
rect 513257 366804 513329 366860
rect 512367 366756 512384 366790
rect 512418 366770 512439 366790
rect 512367 366736 512386 366756
rect 512420 366736 512439 366770
rect 512367 366731 512439 366736
rect 513257 366770 513276 366804
rect 513310 366770 513329 366804
rect 513257 366731 513329 366770
rect 512367 366712 513329 366731
rect 512367 366700 512462 366712
rect 512367 366666 512384 366700
rect 512418 366678 512462 366700
rect 512496 366678 512552 366712
rect 512586 366678 512642 366712
rect 512676 366678 512732 366712
rect 512766 366678 512822 366712
rect 512856 366678 512912 366712
rect 512946 366678 513002 366712
rect 513036 366678 513092 366712
rect 513126 366678 513182 366712
rect 513216 366678 513329 366712
rect 512418 366666 513329 366678
rect 512367 366659 513329 366666
rect 513393 367620 513426 367654
rect 513460 367620 513492 367654
rect 513393 367564 513492 367620
rect 513393 367530 513426 367564
rect 513460 367530 513492 367564
rect 513393 367474 513492 367530
rect 513393 367440 513426 367474
rect 513460 367440 513492 367474
rect 513393 367384 513492 367440
rect 513393 367350 513426 367384
rect 513460 367350 513492 367384
rect 513393 367294 513492 367350
rect 513393 367260 513426 367294
rect 513460 367260 513492 367294
rect 513393 367204 513492 367260
rect 513393 367170 513426 367204
rect 513460 367170 513492 367204
rect 513393 367114 513492 367170
rect 513393 367080 513426 367114
rect 513460 367080 513492 367114
rect 513393 367024 513492 367080
rect 513393 366990 513426 367024
rect 513460 366990 513492 367024
rect 513393 366934 513492 366990
rect 513393 366900 513426 366934
rect 513460 366900 513492 366934
rect 513393 366844 513492 366900
rect 513393 366810 513426 366844
rect 513460 366810 513492 366844
rect 513393 366754 513492 366810
rect 513393 366720 513426 366754
rect 513460 366720 513492 366754
rect 513393 366664 513492 366720
rect 512204 366595 512303 366630
rect 513393 366630 513426 366664
rect 513460 366630 513492 366664
rect 513393 366595 513492 366630
rect 512204 366594 513492 366595
rect 512204 366560 512224 366594
rect 512258 366563 513492 366594
rect 512258 366560 512262 366563
rect 512204 366529 512262 366560
rect 512296 366529 512352 366563
rect 512386 366529 512442 366563
rect 512476 366529 512532 366563
rect 512566 366529 512622 366563
rect 512656 366529 512712 366563
rect 512746 366529 512802 366563
rect 512836 366529 512892 366563
rect 512926 366529 512982 366563
rect 513016 366529 513072 366563
rect 513106 366529 513162 366563
rect 513196 366529 513252 366563
rect 513286 366529 513342 366563
rect 513376 366529 513492 366563
rect 512204 366424 513492 366529
rect 512204 366390 512224 366424
rect 512258 366410 513492 366424
rect 512258 366390 512262 366410
rect 512204 366376 512262 366390
rect 512296 366376 512352 366410
rect 512386 366376 512442 366410
rect 512476 366376 512532 366410
rect 512566 366376 512622 366410
rect 512656 366376 512712 366410
rect 512746 366376 512802 366410
rect 512836 366376 512892 366410
rect 512926 366376 512982 366410
rect 513016 366376 513072 366410
rect 513106 366376 513162 366410
rect 513196 366376 513252 366410
rect 513286 366376 513342 366410
rect 513376 366376 513492 366410
rect 512204 366345 513492 366376
rect 512204 366334 512303 366345
rect 512204 366300 512224 366334
rect 512258 366314 512303 366334
rect 512204 366280 512239 366300
rect 512273 366280 512303 366314
rect 513393 366314 513492 366345
rect 512204 366244 512303 366280
rect 512204 366210 512224 366244
rect 512258 366224 512303 366244
rect 512204 366190 512239 366210
rect 512273 366190 512303 366224
rect 512204 366154 512303 366190
rect 512204 366120 512224 366154
rect 512258 366134 512303 366154
rect 512204 366100 512239 366120
rect 512273 366100 512303 366134
rect 512204 366064 512303 366100
rect 512204 366030 512224 366064
rect 512258 366044 512303 366064
rect 512204 366010 512239 366030
rect 512273 366010 512303 366044
rect 512204 365974 512303 366010
rect 512204 365940 512224 365974
rect 512258 365954 512303 365974
rect 512204 365920 512239 365940
rect 512273 365920 512303 365954
rect 512204 365884 512303 365920
rect 512204 365850 512224 365884
rect 512258 365864 512303 365884
rect 512204 365830 512239 365850
rect 512273 365830 512303 365864
rect 512204 365794 512303 365830
rect 512204 365760 512224 365794
rect 512258 365774 512303 365794
rect 512204 365740 512239 365760
rect 512273 365740 512303 365774
rect 512204 365704 512303 365740
rect 512204 365670 512224 365704
rect 512258 365684 512303 365704
rect 512204 365650 512239 365670
rect 512273 365650 512303 365684
rect 512204 365614 512303 365650
rect 512204 365580 512224 365614
rect 512258 365594 512303 365614
rect 512204 365560 512239 365580
rect 512273 365560 512303 365594
rect 512204 365524 512303 365560
rect 512204 365490 512224 365524
rect 512258 365504 512303 365524
rect 512204 365470 512239 365490
rect 512273 365470 512303 365504
rect 512204 365434 512303 365470
rect 512204 365400 512224 365434
rect 512258 365414 512303 365434
rect 512204 365380 512239 365400
rect 512273 365380 512303 365414
rect 512204 365344 512303 365380
rect 512204 365310 512224 365344
rect 512258 365324 512303 365344
rect 512204 365290 512239 365310
rect 512273 365290 512303 365324
rect 512367 366262 513329 366281
rect 512367 366260 512443 366262
rect 512367 366226 512384 366260
rect 512418 366228 512443 366260
rect 512477 366228 512533 366262
rect 512567 366228 512623 366262
rect 512657 366228 512713 366262
rect 512747 366228 512803 366262
rect 512837 366228 512893 366262
rect 512927 366228 512983 366262
rect 513017 366228 513073 366262
rect 513107 366228 513163 366262
rect 513197 366228 513329 366262
rect 512418 366226 513329 366228
rect 512367 366209 513329 366226
rect 512367 366170 512439 366209
rect 512367 366136 512384 366170
rect 512418 366150 512439 366170
rect 512367 366116 512386 366136
rect 512420 366116 512439 366150
rect 513257 366184 513329 366209
rect 513257 366150 513276 366184
rect 513310 366150 513329 366184
rect 512367 366080 512439 366116
rect 512367 366046 512384 366080
rect 512418 366060 512439 366080
rect 512367 366026 512386 366046
rect 512420 366026 512439 366060
rect 512367 365990 512439 366026
rect 512367 365956 512384 365990
rect 512418 365970 512439 365990
rect 512367 365936 512386 365956
rect 512420 365936 512439 365970
rect 512367 365900 512439 365936
rect 512367 365866 512384 365900
rect 512418 365880 512439 365900
rect 512367 365846 512386 365866
rect 512420 365846 512439 365880
rect 512367 365810 512439 365846
rect 512367 365776 512384 365810
rect 512418 365790 512439 365810
rect 512367 365756 512386 365776
rect 512420 365756 512439 365790
rect 512367 365720 512439 365756
rect 512367 365686 512384 365720
rect 512418 365700 512439 365720
rect 512367 365666 512386 365686
rect 512420 365666 512439 365700
rect 512367 365630 512439 365666
rect 512367 365596 512384 365630
rect 512418 365610 512439 365630
rect 512367 365576 512386 365596
rect 512420 365576 512439 365610
rect 512367 365540 512439 365576
rect 512367 365506 512384 365540
rect 512418 365520 512439 365540
rect 512367 365486 512386 365506
rect 512420 365486 512439 365520
rect 512367 365450 512439 365486
rect 512501 366086 513195 366147
rect 512501 366052 512560 366086
rect 512594 366074 512650 366086
rect 512622 366052 512650 366074
rect 512684 366074 512740 366086
rect 512684 366052 512688 366074
rect 512501 366040 512588 366052
rect 512622 366040 512688 366052
rect 512722 366052 512740 366074
rect 512774 366074 512830 366086
rect 512774 366052 512788 366074
rect 512722 366040 512788 366052
rect 512822 366052 512830 366074
rect 512864 366074 512920 366086
rect 512954 366074 513010 366086
rect 513044 366074 513100 366086
rect 512864 366052 512888 366074
rect 512954 366052 512988 366074
rect 513044 366052 513088 366074
rect 513134 366052 513195 366086
rect 512822 366040 512888 366052
rect 512922 366040 512988 366052
rect 513022 366040 513088 366052
rect 513122 366040 513195 366052
rect 512501 365996 513195 366040
rect 512501 365962 512560 365996
rect 512594 365974 512650 365996
rect 512622 365962 512650 365974
rect 512684 365974 512740 365996
rect 512684 365962 512688 365974
rect 512501 365940 512588 365962
rect 512622 365940 512688 365962
rect 512722 365962 512740 365974
rect 512774 365974 512830 365996
rect 512774 365962 512788 365974
rect 512722 365940 512788 365962
rect 512822 365962 512830 365974
rect 512864 365974 512920 365996
rect 512954 365974 513010 365996
rect 513044 365974 513100 365996
rect 512864 365962 512888 365974
rect 512954 365962 512988 365974
rect 513044 365962 513088 365974
rect 513134 365962 513195 365996
rect 512822 365940 512888 365962
rect 512922 365940 512988 365962
rect 513022 365940 513088 365962
rect 513122 365940 513195 365962
rect 512501 365906 513195 365940
rect 512501 365872 512560 365906
rect 512594 365874 512650 365906
rect 512622 365872 512650 365874
rect 512684 365874 512740 365906
rect 512684 365872 512688 365874
rect 512501 365840 512588 365872
rect 512622 365840 512688 365872
rect 512722 365872 512740 365874
rect 512774 365874 512830 365906
rect 512774 365872 512788 365874
rect 512722 365840 512788 365872
rect 512822 365872 512830 365874
rect 512864 365874 512920 365906
rect 512954 365874 513010 365906
rect 513044 365874 513100 365906
rect 512864 365872 512888 365874
rect 512954 365872 512988 365874
rect 513044 365872 513088 365874
rect 513134 365872 513195 365906
rect 512822 365840 512888 365872
rect 512922 365840 512988 365872
rect 513022 365840 513088 365872
rect 513122 365840 513195 365872
rect 512501 365816 513195 365840
rect 512501 365782 512560 365816
rect 512594 365782 512650 365816
rect 512684 365782 512740 365816
rect 512774 365782 512830 365816
rect 512864 365782 512920 365816
rect 512954 365782 513010 365816
rect 513044 365782 513100 365816
rect 513134 365782 513195 365816
rect 512501 365774 513195 365782
rect 512501 365740 512588 365774
rect 512622 365740 512688 365774
rect 512722 365740 512788 365774
rect 512822 365740 512888 365774
rect 512922 365740 512988 365774
rect 513022 365740 513088 365774
rect 513122 365740 513195 365774
rect 512501 365726 513195 365740
rect 512501 365692 512560 365726
rect 512594 365692 512650 365726
rect 512684 365692 512740 365726
rect 512774 365692 512830 365726
rect 512864 365692 512920 365726
rect 512954 365692 513010 365726
rect 513044 365692 513100 365726
rect 513134 365692 513195 365726
rect 512501 365674 513195 365692
rect 512501 365640 512588 365674
rect 512622 365640 512688 365674
rect 512722 365640 512788 365674
rect 512822 365640 512888 365674
rect 512922 365640 512988 365674
rect 513022 365640 513088 365674
rect 513122 365640 513195 365674
rect 512501 365636 513195 365640
rect 512501 365602 512560 365636
rect 512594 365602 512650 365636
rect 512684 365602 512740 365636
rect 512774 365602 512830 365636
rect 512864 365602 512920 365636
rect 512954 365602 513010 365636
rect 513044 365602 513100 365636
rect 513134 365602 513195 365636
rect 512501 365574 513195 365602
rect 512501 365546 512588 365574
rect 512622 365546 512688 365574
rect 512501 365512 512560 365546
rect 512622 365540 512650 365546
rect 512594 365512 512650 365540
rect 512684 365540 512688 365546
rect 512722 365546 512788 365574
rect 512722 365540 512740 365546
rect 512684 365512 512740 365540
rect 512774 365540 512788 365546
rect 512822 365546 512888 365574
rect 512922 365546 512988 365574
rect 513022 365546 513088 365574
rect 513122 365546 513195 365574
rect 512822 365540 512830 365546
rect 512774 365512 512830 365540
rect 512864 365540 512888 365546
rect 512954 365540 512988 365546
rect 513044 365540 513088 365546
rect 512864 365512 512920 365540
rect 512954 365512 513010 365540
rect 513044 365512 513100 365540
rect 513134 365512 513195 365546
rect 512501 365453 513195 365512
rect 513257 366094 513329 366150
rect 513257 366060 513276 366094
rect 513310 366060 513329 366094
rect 513257 366004 513329 366060
rect 513257 365970 513276 366004
rect 513310 365970 513329 366004
rect 513257 365914 513329 365970
rect 513257 365880 513276 365914
rect 513310 365880 513329 365914
rect 513257 365824 513329 365880
rect 513257 365790 513276 365824
rect 513310 365790 513329 365824
rect 513257 365734 513329 365790
rect 513257 365700 513276 365734
rect 513310 365700 513329 365734
rect 513257 365644 513329 365700
rect 513257 365610 513276 365644
rect 513310 365610 513329 365644
rect 513257 365554 513329 365610
rect 513257 365520 513276 365554
rect 513310 365520 513329 365554
rect 513257 365464 513329 365520
rect 512367 365416 512384 365450
rect 512418 365430 512439 365450
rect 512367 365396 512386 365416
rect 512420 365396 512439 365430
rect 512367 365391 512439 365396
rect 513257 365430 513276 365464
rect 513310 365430 513329 365464
rect 513257 365391 513329 365430
rect 512367 365372 513329 365391
rect 512367 365360 512462 365372
rect 512367 365326 512384 365360
rect 512418 365338 512462 365360
rect 512496 365338 512552 365372
rect 512586 365338 512642 365372
rect 512676 365338 512732 365372
rect 512766 365338 512822 365372
rect 512856 365338 512912 365372
rect 512946 365338 513002 365372
rect 513036 365338 513092 365372
rect 513126 365338 513182 365372
rect 513216 365338 513329 365372
rect 512418 365326 513329 365338
rect 512367 365319 513329 365326
rect 513393 366280 513426 366314
rect 513460 366280 513492 366314
rect 513393 366224 513492 366280
rect 513393 366190 513426 366224
rect 513460 366190 513492 366224
rect 513393 366134 513492 366190
rect 513393 366100 513426 366134
rect 513460 366100 513492 366134
rect 513393 366044 513492 366100
rect 513393 366010 513426 366044
rect 513460 366010 513492 366044
rect 513393 365954 513492 366010
rect 513393 365920 513426 365954
rect 513460 365920 513492 365954
rect 513393 365864 513492 365920
rect 513393 365830 513426 365864
rect 513460 365830 513492 365864
rect 513393 365774 513492 365830
rect 513393 365740 513426 365774
rect 513460 365740 513492 365774
rect 513393 365684 513492 365740
rect 513393 365650 513426 365684
rect 513460 365650 513492 365684
rect 513393 365594 513492 365650
rect 513393 365560 513426 365594
rect 513460 365560 513492 365594
rect 513393 365504 513492 365560
rect 513393 365470 513426 365504
rect 513460 365470 513492 365504
rect 513393 365414 513492 365470
rect 513393 365380 513426 365414
rect 513460 365380 513492 365414
rect 513393 365324 513492 365380
rect 512204 365255 512303 365290
rect 513393 365290 513426 365324
rect 513460 365290 513492 365324
rect 513393 365255 513492 365290
rect 512204 365254 513492 365255
rect 512204 365220 512224 365254
rect 512258 365223 513492 365254
rect 512258 365220 512262 365223
rect 512204 365189 512262 365220
rect 512296 365189 512352 365223
rect 512386 365189 512442 365223
rect 512476 365189 512532 365223
rect 512566 365189 512622 365223
rect 512656 365189 512712 365223
rect 512746 365189 512802 365223
rect 512836 365189 512892 365223
rect 512926 365189 512982 365223
rect 513016 365189 513072 365223
rect 513106 365189 513162 365223
rect 513196 365189 513252 365223
rect 513286 365189 513342 365223
rect 513376 365189 513492 365223
rect 512204 365084 513492 365189
rect 512204 365050 512224 365084
rect 512258 365070 513492 365084
rect 512258 365050 512262 365070
rect 512204 365036 512262 365050
rect 512296 365036 512352 365070
rect 512386 365036 512442 365070
rect 512476 365036 512532 365070
rect 512566 365036 512622 365070
rect 512656 365036 512712 365070
rect 512746 365036 512802 365070
rect 512836 365036 512892 365070
rect 512926 365036 512982 365070
rect 513016 365036 513072 365070
rect 513106 365036 513162 365070
rect 513196 365036 513252 365070
rect 513286 365036 513342 365070
rect 513376 365036 513492 365070
rect 512204 365005 513492 365036
rect 512204 364994 512303 365005
rect 512204 364960 512224 364994
rect 512258 364974 512303 364994
rect 512204 364940 512239 364960
rect 512273 364940 512303 364974
rect 513393 364974 513492 365005
rect 512204 364904 512303 364940
rect 512204 364870 512224 364904
rect 512258 364884 512303 364904
rect 512204 364850 512239 364870
rect 512273 364850 512303 364884
rect 512204 364814 512303 364850
rect 512204 364780 512224 364814
rect 512258 364794 512303 364814
rect 512204 364760 512239 364780
rect 512273 364760 512303 364794
rect 512204 364724 512303 364760
rect 512204 364690 512224 364724
rect 512258 364704 512303 364724
rect 512204 364670 512239 364690
rect 512273 364670 512303 364704
rect 512204 364634 512303 364670
rect 512204 364600 512224 364634
rect 512258 364614 512303 364634
rect 512204 364580 512239 364600
rect 512273 364580 512303 364614
rect 512204 364544 512303 364580
rect 512204 364510 512224 364544
rect 512258 364524 512303 364544
rect 512204 364490 512239 364510
rect 512273 364490 512303 364524
rect 512204 364454 512303 364490
rect 512204 364420 512224 364454
rect 512258 364434 512303 364454
rect 512204 364400 512239 364420
rect 512273 364400 512303 364434
rect 512204 364364 512303 364400
rect 512204 364330 512224 364364
rect 512258 364344 512303 364364
rect 512204 364310 512239 364330
rect 512273 364310 512303 364344
rect 512204 364274 512303 364310
rect 512204 364240 512224 364274
rect 512258 364254 512303 364274
rect 512204 364220 512239 364240
rect 512273 364220 512303 364254
rect 512204 364184 512303 364220
rect 512204 364150 512224 364184
rect 512258 364164 512303 364184
rect 512204 364130 512239 364150
rect 512273 364130 512303 364164
rect 512204 364094 512303 364130
rect 512204 364060 512224 364094
rect 512258 364074 512303 364094
rect 512204 364040 512239 364060
rect 512273 364040 512303 364074
rect 512204 364004 512303 364040
rect 512204 363970 512224 364004
rect 512258 363984 512303 364004
rect 512204 363950 512239 363970
rect 512273 363950 512303 363984
rect 512367 364922 513329 364941
rect 512367 364920 512443 364922
rect 512367 364886 512384 364920
rect 512418 364888 512443 364920
rect 512477 364888 512533 364922
rect 512567 364888 512623 364922
rect 512657 364888 512713 364922
rect 512747 364888 512803 364922
rect 512837 364888 512893 364922
rect 512927 364888 512983 364922
rect 513017 364888 513073 364922
rect 513107 364888 513163 364922
rect 513197 364888 513329 364922
rect 512418 364886 513329 364888
rect 512367 364869 513329 364886
rect 512367 364830 512439 364869
rect 512367 364796 512384 364830
rect 512418 364810 512439 364830
rect 512367 364776 512386 364796
rect 512420 364776 512439 364810
rect 513257 364844 513329 364869
rect 513257 364810 513276 364844
rect 513310 364810 513329 364844
rect 512367 364740 512439 364776
rect 512367 364706 512384 364740
rect 512418 364720 512439 364740
rect 512367 364686 512386 364706
rect 512420 364686 512439 364720
rect 512367 364650 512439 364686
rect 512367 364616 512384 364650
rect 512418 364630 512439 364650
rect 512367 364596 512386 364616
rect 512420 364596 512439 364630
rect 512367 364560 512439 364596
rect 512367 364526 512384 364560
rect 512418 364540 512439 364560
rect 512367 364506 512386 364526
rect 512420 364506 512439 364540
rect 512367 364470 512439 364506
rect 512367 364436 512384 364470
rect 512418 364450 512439 364470
rect 512367 364416 512386 364436
rect 512420 364416 512439 364450
rect 512367 364380 512439 364416
rect 512367 364346 512384 364380
rect 512418 364360 512439 364380
rect 512367 364326 512386 364346
rect 512420 364326 512439 364360
rect 512367 364290 512439 364326
rect 512367 364256 512384 364290
rect 512418 364270 512439 364290
rect 512367 364236 512386 364256
rect 512420 364236 512439 364270
rect 512367 364200 512439 364236
rect 512367 364166 512384 364200
rect 512418 364180 512439 364200
rect 512367 364146 512386 364166
rect 512420 364146 512439 364180
rect 512367 364110 512439 364146
rect 512501 364746 513195 364807
rect 512501 364712 512560 364746
rect 512594 364734 512650 364746
rect 512622 364712 512650 364734
rect 512684 364734 512740 364746
rect 512684 364712 512688 364734
rect 512501 364700 512588 364712
rect 512622 364700 512688 364712
rect 512722 364712 512740 364734
rect 512774 364734 512830 364746
rect 512774 364712 512788 364734
rect 512722 364700 512788 364712
rect 512822 364712 512830 364734
rect 512864 364734 512920 364746
rect 512954 364734 513010 364746
rect 513044 364734 513100 364746
rect 512864 364712 512888 364734
rect 512954 364712 512988 364734
rect 513044 364712 513088 364734
rect 513134 364712 513195 364746
rect 512822 364700 512888 364712
rect 512922 364700 512988 364712
rect 513022 364700 513088 364712
rect 513122 364700 513195 364712
rect 512501 364656 513195 364700
rect 512501 364622 512560 364656
rect 512594 364634 512650 364656
rect 512622 364622 512650 364634
rect 512684 364634 512740 364656
rect 512684 364622 512688 364634
rect 512501 364600 512588 364622
rect 512622 364600 512688 364622
rect 512722 364622 512740 364634
rect 512774 364634 512830 364656
rect 512774 364622 512788 364634
rect 512722 364600 512788 364622
rect 512822 364622 512830 364634
rect 512864 364634 512920 364656
rect 512954 364634 513010 364656
rect 513044 364634 513100 364656
rect 512864 364622 512888 364634
rect 512954 364622 512988 364634
rect 513044 364622 513088 364634
rect 513134 364622 513195 364656
rect 512822 364600 512888 364622
rect 512922 364600 512988 364622
rect 513022 364600 513088 364622
rect 513122 364600 513195 364622
rect 512501 364566 513195 364600
rect 512501 364532 512560 364566
rect 512594 364534 512650 364566
rect 512622 364532 512650 364534
rect 512684 364534 512740 364566
rect 512684 364532 512688 364534
rect 512501 364500 512588 364532
rect 512622 364500 512688 364532
rect 512722 364532 512740 364534
rect 512774 364534 512830 364566
rect 512774 364532 512788 364534
rect 512722 364500 512788 364532
rect 512822 364532 512830 364534
rect 512864 364534 512920 364566
rect 512954 364534 513010 364566
rect 513044 364534 513100 364566
rect 512864 364532 512888 364534
rect 512954 364532 512988 364534
rect 513044 364532 513088 364534
rect 513134 364532 513195 364566
rect 512822 364500 512888 364532
rect 512922 364500 512988 364532
rect 513022 364500 513088 364532
rect 513122 364500 513195 364532
rect 512501 364476 513195 364500
rect 512501 364442 512560 364476
rect 512594 364442 512650 364476
rect 512684 364442 512740 364476
rect 512774 364442 512830 364476
rect 512864 364442 512920 364476
rect 512954 364442 513010 364476
rect 513044 364442 513100 364476
rect 513134 364442 513195 364476
rect 512501 364434 513195 364442
rect 512501 364400 512588 364434
rect 512622 364400 512688 364434
rect 512722 364400 512788 364434
rect 512822 364400 512888 364434
rect 512922 364400 512988 364434
rect 513022 364400 513088 364434
rect 513122 364400 513195 364434
rect 512501 364386 513195 364400
rect 512501 364352 512560 364386
rect 512594 364352 512650 364386
rect 512684 364352 512740 364386
rect 512774 364352 512830 364386
rect 512864 364352 512920 364386
rect 512954 364352 513010 364386
rect 513044 364352 513100 364386
rect 513134 364352 513195 364386
rect 512501 364334 513195 364352
rect 512501 364300 512588 364334
rect 512622 364300 512688 364334
rect 512722 364300 512788 364334
rect 512822 364300 512888 364334
rect 512922 364300 512988 364334
rect 513022 364300 513088 364334
rect 513122 364300 513195 364334
rect 512501 364296 513195 364300
rect 512501 364262 512560 364296
rect 512594 364262 512650 364296
rect 512684 364262 512740 364296
rect 512774 364262 512830 364296
rect 512864 364262 512920 364296
rect 512954 364262 513010 364296
rect 513044 364262 513100 364296
rect 513134 364262 513195 364296
rect 512501 364234 513195 364262
rect 512501 364206 512588 364234
rect 512622 364206 512688 364234
rect 512501 364172 512560 364206
rect 512622 364200 512650 364206
rect 512594 364172 512650 364200
rect 512684 364200 512688 364206
rect 512722 364206 512788 364234
rect 512722 364200 512740 364206
rect 512684 364172 512740 364200
rect 512774 364200 512788 364206
rect 512822 364206 512888 364234
rect 512922 364206 512988 364234
rect 513022 364206 513088 364234
rect 513122 364206 513195 364234
rect 512822 364200 512830 364206
rect 512774 364172 512830 364200
rect 512864 364200 512888 364206
rect 512954 364200 512988 364206
rect 513044 364200 513088 364206
rect 512864 364172 512920 364200
rect 512954 364172 513010 364200
rect 513044 364172 513100 364200
rect 513134 364172 513195 364206
rect 512501 364113 513195 364172
rect 513257 364754 513329 364810
rect 513257 364720 513276 364754
rect 513310 364720 513329 364754
rect 513257 364664 513329 364720
rect 513257 364630 513276 364664
rect 513310 364630 513329 364664
rect 513257 364574 513329 364630
rect 513257 364540 513276 364574
rect 513310 364540 513329 364574
rect 513257 364484 513329 364540
rect 513257 364450 513276 364484
rect 513310 364450 513329 364484
rect 513257 364394 513329 364450
rect 513257 364360 513276 364394
rect 513310 364360 513329 364394
rect 513257 364304 513329 364360
rect 513257 364270 513276 364304
rect 513310 364270 513329 364304
rect 513257 364214 513329 364270
rect 513257 364180 513276 364214
rect 513310 364180 513329 364214
rect 513257 364124 513329 364180
rect 512367 364076 512384 364110
rect 512418 364090 512439 364110
rect 512367 364056 512386 364076
rect 512420 364056 512439 364090
rect 512367 364051 512439 364056
rect 513257 364090 513276 364124
rect 513310 364090 513329 364124
rect 513257 364051 513329 364090
rect 512367 364032 513329 364051
rect 512367 364020 512462 364032
rect 512367 363986 512384 364020
rect 512418 363998 512462 364020
rect 512496 363998 512552 364032
rect 512586 363998 512642 364032
rect 512676 363998 512732 364032
rect 512766 363998 512822 364032
rect 512856 363998 512912 364032
rect 512946 363998 513002 364032
rect 513036 363998 513092 364032
rect 513126 363998 513182 364032
rect 513216 363998 513329 364032
rect 512418 363986 513329 363998
rect 512367 363979 513329 363986
rect 513393 364940 513426 364974
rect 513460 364940 513492 364974
rect 513393 364884 513492 364940
rect 513393 364850 513426 364884
rect 513460 364850 513492 364884
rect 513393 364794 513492 364850
rect 513393 364760 513426 364794
rect 513460 364760 513492 364794
rect 513393 364704 513492 364760
rect 513393 364670 513426 364704
rect 513460 364670 513492 364704
rect 513393 364614 513492 364670
rect 513393 364580 513426 364614
rect 513460 364580 513492 364614
rect 513393 364524 513492 364580
rect 513393 364490 513426 364524
rect 513460 364490 513492 364524
rect 513393 364434 513492 364490
rect 513393 364400 513426 364434
rect 513460 364400 513492 364434
rect 513393 364344 513492 364400
rect 513393 364310 513426 364344
rect 513460 364310 513492 364344
rect 513393 364254 513492 364310
rect 513393 364220 513426 364254
rect 513460 364220 513492 364254
rect 513393 364164 513492 364220
rect 513393 364130 513426 364164
rect 513460 364130 513492 364164
rect 513393 364074 513492 364130
rect 513393 364040 513426 364074
rect 513460 364040 513492 364074
rect 513393 363984 513492 364040
rect 512204 363915 512303 363950
rect 513393 363950 513426 363984
rect 513460 363950 513492 363984
rect 513393 363915 513492 363950
rect 512204 363914 513492 363915
rect 512204 363880 512224 363914
rect 512258 363883 513492 363914
rect 512258 363880 512262 363883
rect 512204 363849 512262 363880
rect 512296 363849 512352 363883
rect 512386 363849 512442 363883
rect 512476 363849 512532 363883
rect 512566 363849 512622 363883
rect 512656 363849 512712 363883
rect 512746 363849 512802 363883
rect 512836 363849 512892 363883
rect 512926 363849 512982 363883
rect 513016 363849 513072 363883
rect 513106 363849 513162 363883
rect 513196 363849 513252 363883
rect 513286 363849 513342 363883
rect 513376 363849 513492 363883
rect 512204 363744 513492 363849
rect 512204 363710 512224 363744
rect 512258 363730 513492 363744
rect 512258 363710 512262 363730
rect 512204 363696 512262 363710
rect 512296 363696 512352 363730
rect 512386 363696 512442 363730
rect 512476 363696 512532 363730
rect 512566 363696 512622 363730
rect 512656 363696 512712 363730
rect 512746 363696 512802 363730
rect 512836 363696 512892 363730
rect 512926 363696 512982 363730
rect 513016 363696 513072 363730
rect 513106 363696 513162 363730
rect 513196 363696 513252 363730
rect 513286 363696 513342 363730
rect 513376 363696 513492 363730
rect 512204 363665 513492 363696
rect 512204 363654 512303 363665
rect 512204 363620 512224 363654
rect 512258 363634 512303 363654
rect 512204 363600 512239 363620
rect 512273 363600 512303 363634
rect 513393 363634 513492 363665
rect 512204 363564 512303 363600
rect 512204 363530 512224 363564
rect 512258 363544 512303 363564
rect 512204 363510 512239 363530
rect 512273 363510 512303 363544
rect 512204 363474 512303 363510
rect 512204 363440 512224 363474
rect 512258 363454 512303 363474
rect 512204 363420 512239 363440
rect 512273 363420 512303 363454
rect 512204 363384 512303 363420
rect 512204 363350 512224 363384
rect 512258 363364 512303 363384
rect 512204 363330 512239 363350
rect 512273 363330 512303 363364
rect 512204 363294 512303 363330
rect 512204 363260 512224 363294
rect 512258 363274 512303 363294
rect 512204 363240 512239 363260
rect 512273 363240 512303 363274
rect 512204 363204 512303 363240
rect 512204 363170 512224 363204
rect 512258 363184 512303 363204
rect 512204 363150 512239 363170
rect 512273 363150 512303 363184
rect 512204 363114 512303 363150
rect 512204 363080 512224 363114
rect 512258 363094 512303 363114
rect 512204 363060 512239 363080
rect 512273 363060 512303 363094
rect 512204 363024 512303 363060
rect 512204 362990 512224 363024
rect 512258 363004 512303 363024
rect 512204 362970 512239 362990
rect 512273 362970 512303 363004
rect 512204 362934 512303 362970
rect 512204 362900 512224 362934
rect 512258 362914 512303 362934
rect 512204 362880 512239 362900
rect 512273 362880 512303 362914
rect 512204 362844 512303 362880
rect 512204 362810 512224 362844
rect 512258 362824 512303 362844
rect 512204 362790 512239 362810
rect 512273 362790 512303 362824
rect 512204 362754 512303 362790
rect 512204 362720 512224 362754
rect 512258 362734 512303 362754
rect 512204 362700 512239 362720
rect 512273 362700 512303 362734
rect 512204 362664 512303 362700
rect 512204 362630 512224 362664
rect 512258 362644 512303 362664
rect 512204 362610 512239 362630
rect 512273 362610 512303 362644
rect 512367 363582 513329 363601
rect 512367 363580 512443 363582
rect 512367 363546 512384 363580
rect 512418 363548 512443 363580
rect 512477 363548 512533 363582
rect 512567 363548 512623 363582
rect 512657 363548 512713 363582
rect 512747 363548 512803 363582
rect 512837 363548 512893 363582
rect 512927 363548 512983 363582
rect 513017 363548 513073 363582
rect 513107 363548 513163 363582
rect 513197 363548 513329 363582
rect 512418 363546 513329 363548
rect 512367 363529 513329 363546
rect 512367 363490 512439 363529
rect 512367 363456 512384 363490
rect 512418 363470 512439 363490
rect 512367 363436 512386 363456
rect 512420 363436 512439 363470
rect 513257 363504 513329 363529
rect 513257 363470 513276 363504
rect 513310 363470 513329 363504
rect 512367 363400 512439 363436
rect 512367 363366 512384 363400
rect 512418 363380 512439 363400
rect 512367 363346 512386 363366
rect 512420 363346 512439 363380
rect 512367 363310 512439 363346
rect 512367 363276 512384 363310
rect 512418 363290 512439 363310
rect 512367 363256 512386 363276
rect 512420 363256 512439 363290
rect 512367 363220 512439 363256
rect 512367 363186 512384 363220
rect 512418 363200 512439 363220
rect 512367 363166 512386 363186
rect 512420 363166 512439 363200
rect 512367 363130 512439 363166
rect 512367 363096 512384 363130
rect 512418 363110 512439 363130
rect 512367 363076 512386 363096
rect 512420 363076 512439 363110
rect 512367 363040 512439 363076
rect 512367 363006 512384 363040
rect 512418 363020 512439 363040
rect 512367 362986 512386 363006
rect 512420 362986 512439 363020
rect 512367 362950 512439 362986
rect 512367 362916 512384 362950
rect 512418 362930 512439 362950
rect 512367 362896 512386 362916
rect 512420 362896 512439 362930
rect 512367 362860 512439 362896
rect 512367 362826 512384 362860
rect 512418 362840 512439 362860
rect 512367 362806 512386 362826
rect 512420 362806 512439 362840
rect 512367 362770 512439 362806
rect 512501 363406 513195 363467
rect 512501 363372 512560 363406
rect 512594 363394 512650 363406
rect 512622 363372 512650 363394
rect 512684 363394 512740 363406
rect 512684 363372 512688 363394
rect 512501 363360 512588 363372
rect 512622 363360 512688 363372
rect 512722 363372 512740 363394
rect 512774 363394 512830 363406
rect 512774 363372 512788 363394
rect 512722 363360 512788 363372
rect 512822 363372 512830 363394
rect 512864 363394 512920 363406
rect 512954 363394 513010 363406
rect 513044 363394 513100 363406
rect 512864 363372 512888 363394
rect 512954 363372 512988 363394
rect 513044 363372 513088 363394
rect 513134 363372 513195 363406
rect 512822 363360 512888 363372
rect 512922 363360 512988 363372
rect 513022 363360 513088 363372
rect 513122 363360 513195 363372
rect 512501 363316 513195 363360
rect 512501 363282 512560 363316
rect 512594 363294 512650 363316
rect 512622 363282 512650 363294
rect 512684 363294 512740 363316
rect 512684 363282 512688 363294
rect 512501 363260 512588 363282
rect 512622 363260 512688 363282
rect 512722 363282 512740 363294
rect 512774 363294 512830 363316
rect 512774 363282 512788 363294
rect 512722 363260 512788 363282
rect 512822 363282 512830 363294
rect 512864 363294 512920 363316
rect 512954 363294 513010 363316
rect 513044 363294 513100 363316
rect 512864 363282 512888 363294
rect 512954 363282 512988 363294
rect 513044 363282 513088 363294
rect 513134 363282 513195 363316
rect 512822 363260 512888 363282
rect 512922 363260 512988 363282
rect 513022 363260 513088 363282
rect 513122 363260 513195 363282
rect 512501 363226 513195 363260
rect 512501 363192 512560 363226
rect 512594 363194 512650 363226
rect 512622 363192 512650 363194
rect 512684 363194 512740 363226
rect 512684 363192 512688 363194
rect 512501 363160 512588 363192
rect 512622 363160 512688 363192
rect 512722 363192 512740 363194
rect 512774 363194 512830 363226
rect 512774 363192 512788 363194
rect 512722 363160 512788 363192
rect 512822 363192 512830 363194
rect 512864 363194 512920 363226
rect 512954 363194 513010 363226
rect 513044 363194 513100 363226
rect 512864 363192 512888 363194
rect 512954 363192 512988 363194
rect 513044 363192 513088 363194
rect 513134 363192 513195 363226
rect 512822 363160 512888 363192
rect 512922 363160 512988 363192
rect 513022 363160 513088 363192
rect 513122 363160 513195 363192
rect 512501 363136 513195 363160
rect 512501 363102 512560 363136
rect 512594 363102 512650 363136
rect 512684 363102 512740 363136
rect 512774 363102 512830 363136
rect 512864 363102 512920 363136
rect 512954 363102 513010 363136
rect 513044 363102 513100 363136
rect 513134 363102 513195 363136
rect 512501 363094 513195 363102
rect 512501 363060 512588 363094
rect 512622 363060 512688 363094
rect 512722 363060 512788 363094
rect 512822 363060 512888 363094
rect 512922 363060 512988 363094
rect 513022 363060 513088 363094
rect 513122 363060 513195 363094
rect 512501 363046 513195 363060
rect 512501 363012 512560 363046
rect 512594 363012 512650 363046
rect 512684 363012 512740 363046
rect 512774 363012 512830 363046
rect 512864 363012 512920 363046
rect 512954 363012 513010 363046
rect 513044 363012 513100 363046
rect 513134 363012 513195 363046
rect 512501 362994 513195 363012
rect 512501 362960 512588 362994
rect 512622 362960 512688 362994
rect 512722 362960 512788 362994
rect 512822 362960 512888 362994
rect 512922 362960 512988 362994
rect 513022 362960 513088 362994
rect 513122 362960 513195 362994
rect 512501 362956 513195 362960
rect 512501 362922 512560 362956
rect 512594 362922 512650 362956
rect 512684 362922 512740 362956
rect 512774 362922 512830 362956
rect 512864 362922 512920 362956
rect 512954 362922 513010 362956
rect 513044 362922 513100 362956
rect 513134 362922 513195 362956
rect 512501 362894 513195 362922
rect 512501 362866 512588 362894
rect 512622 362866 512688 362894
rect 512501 362832 512560 362866
rect 512622 362860 512650 362866
rect 512594 362832 512650 362860
rect 512684 362860 512688 362866
rect 512722 362866 512788 362894
rect 512722 362860 512740 362866
rect 512684 362832 512740 362860
rect 512774 362860 512788 362866
rect 512822 362866 512888 362894
rect 512922 362866 512988 362894
rect 513022 362866 513088 362894
rect 513122 362866 513195 362894
rect 512822 362860 512830 362866
rect 512774 362832 512830 362860
rect 512864 362860 512888 362866
rect 512954 362860 512988 362866
rect 513044 362860 513088 362866
rect 512864 362832 512920 362860
rect 512954 362832 513010 362860
rect 513044 362832 513100 362860
rect 513134 362832 513195 362866
rect 512501 362773 513195 362832
rect 513257 363414 513329 363470
rect 513257 363380 513276 363414
rect 513310 363380 513329 363414
rect 513257 363324 513329 363380
rect 513257 363290 513276 363324
rect 513310 363290 513329 363324
rect 513257 363234 513329 363290
rect 513257 363200 513276 363234
rect 513310 363200 513329 363234
rect 513257 363144 513329 363200
rect 513257 363110 513276 363144
rect 513310 363110 513329 363144
rect 513257 363054 513329 363110
rect 513257 363020 513276 363054
rect 513310 363020 513329 363054
rect 513257 362964 513329 363020
rect 513257 362930 513276 362964
rect 513310 362930 513329 362964
rect 513257 362874 513329 362930
rect 513257 362840 513276 362874
rect 513310 362840 513329 362874
rect 513257 362784 513329 362840
rect 512367 362736 512384 362770
rect 512418 362750 512439 362770
rect 512367 362716 512386 362736
rect 512420 362716 512439 362750
rect 512367 362711 512439 362716
rect 513257 362750 513276 362784
rect 513310 362750 513329 362784
rect 513257 362711 513329 362750
rect 512367 362692 513329 362711
rect 512367 362680 512462 362692
rect 512367 362646 512384 362680
rect 512418 362658 512462 362680
rect 512496 362658 512552 362692
rect 512586 362658 512642 362692
rect 512676 362658 512732 362692
rect 512766 362658 512822 362692
rect 512856 362658 512912 362692
rect 512946 362658 513002 362692
rect 513036 362658 513092 362692
rect 513126 362658 513182 362692
rect 513216 362658 513329 362692
rect 512418 362646 513329 362658
rect 512367 362639 513329 362646
rect 513393 363600 513426 363634
rect 513460 363600 513492 363634
rect 513393 363544 513492 363600
rect 513393 363510 513426 363544
rect 513460 363510 513492 363544
rect 513393 363454 513492 363510
rect 513393 363420 513426 363454
rect 513460 363420 513492 363454
rect 513393 363364 513492 363420
rect 513393 363330 513426 363364
rect 513460 363330 513492 363364
rect 513393 363274 513492 363330
rect 513393 363240 513426 363274
rect 513460 363240 513492 363274
rect 513393 363184 513492 363240
rect 513393 363150 513426 363184
rect 513460 363150 513492 363184
rect 513393 363094 513492 363150
rect 513393 363060 513426 363094
rect 513460 363060 513492 363094
rect 513393 363004 513492 363060
rect 513393 362970 513426 363004
rect 513460 362970 513492 363004
rect 513393 362914 513492 362970
rect 513393 362880 513426 362914
rect 513460 362880 513492 362914
rect 513393 362824 513492 362880
rect 513393 362790 513426 362824
rect 513460 362790 513492 362824
rect 513393 362734 513492 362790
rect 513393 362700 513426 362734
rect 513460 362700 513492 362734
rect 513393 362644 513492 362700
rect 512204 362575 512303 362610
rect 513393 362610 513426 362644
rect 513460 362610 513492 362644
rect 513393 362575 513492 362610
rect 512204 362574 513492 362575
rect 512204 362540 512224 362574
rect 512258 362543 513492 362574
rect 512258 362540 512262 362543
rect 512204 362509 512262 362540
rect 512296 362509 512352 362543
rect 512386 362509 512442 362543
rect 512476 362509 512532 362543
rect 512566 362509 512622 362543
rect 512656 362509 512712 362543
rect 512746 362509 512802 362543
rect 512836 362509 512892 362543
rect 512926 362509 512982 362543
rect 513016 362509 513072 362543
rect 513106 362509 513162 362543
rect 513196 362509 513252 362543
rect 513286 362509 513342 362543
rect 513376 362509 513492 362543
rect 512204 362476 513492 362509
rect 513758 372987 513818 373170
rect 513758 372953 513771 372987
rect 513805 372953 513818 372987
rect 513758 372787 513818 372953
rect 513758 372753 513771 372787
rect 513805 372753 513818 372787
rect 513758 372587 513818 372753
rect 513758 372553 513771 372587
rect 513805 372553 513818 372587
rect 513758 372387 513818 372553
rect 513758 372353 513771 372387
rect 513805 372353 513818 372387
rect 515638 373033 515698 373199
rect 515638 372999 515651 373033
rect 515685 372999 515698 373033
rect 515638 372833 515698 372999
rect 515638 372799 515651 372833
rect 515685 372799 515698 372833
rect 517518 373233 517578 373288
rect 517518 373199 517531 373233
rect 517565 373199 517578 373233
rect 517518 373033 517578 373199
rect 517518 372999 517531 373033
rect 517565 372999 517578 373033
rect 517518 372833 517578 372999
rect 515638 372633 515698 372799
rect 515638 372599 515651 372633
rect 515685 372599 515698 372633
rect 515638 372376 515698 372599
rect 516473 372376 516863 372808
rect 517518 372799 517531 372833
rect 517565 372799 517578 372833
rect 517518 372633 517578 372799
rect 517518 372599 517531 372633
rect 517565 372599 517578 372633
rect 517518 372376 517578 372599
rect 519398 374633 519458 374816
rect 519398 374599 519411 374633
rect 519445 374599 519458 374633
rect 519398 374433 519458 374599
rect 519398 374399 519411 374433
rect 519445 374399 519458 374433
rect 519398 374233 519458 374399
rect 521278 374633 521338 374816
rect 521278 374599 521291 374633
rect 521325 374599 521338 374633
rect 521278 374433 521338 374599
rect 521278 374399 521291 374433
rect 521325 374399 521338 374433
rect 519398 374199 519411 374233
rect 519445 374199 519458 374233
rect 519398 374033 519458 374199
rect 519398 373999 519411 374033
rect 519445 373999 519458 374033
rect 519398 373833 519458 373999
rect 521278 374233 521338 374399
rect 521278 374199 521291 374233
rect 521325 374199 521338 374233
rect 521278 374033 521338 374199
rect 521278 373999 521291 374033
rect 521325 373999 521338 374033
rect 521278 373904 521338 373999
rect 519398 373799 519411 373833
rect 519445 373799 519458 373833
rect 519398 373633 519458 373799
rect 519398 373599 519411 373633
rect 519445 373599 519458 373633
rect 519398 373433 519458 373599
rect 519398 373399 519411 373433
rect 519445 373399 519458 373433
rect 519398 373233 519458 373399
rect 520338 373833 521338 373904
rect 520338 373817 521291 373833
rect 520338 373375 520377 373817
rect 520479 373799 521291 373817
rect 521325 373799 521338 373833
rect 520479 373633 521338 373799
rect 520479 373599 521291 373633
rect 521325 373599 521338 373633
rect 520479 373433 521338 373599
rect 520479 373399 521291 373433
rect 521325 373399 521338 373433
rect 520479 373375 521338 373399
rect 520338 373288 521338 373375
rect 519398 373199 519411 373233
rect 519445 373199 519458 373233
rect 519398 373033 519458 373199
rect 519398 372999 519411 373033
rect 519445 372999 519458 373033
rect 519398 372833 519458 372999
rect 519398 372799 519411 372833
rect 519445 372799 519458 372833
rect 521278 373233 521338 373288
rect 521278 373199 521291 373233
rect 521325 373199 521338 373233
rect 521278 373033 521338 373199
rect 521278 372999 521291 373033
rect 521325 372999 521338 373033
rect 521278 372833 521338 372999
rect 519398 372633 519458 372799
rect 519398 372599 519411 372633
rect 519445 372599 519458 372633
rect 519398 372376 519458 372599
rect 520233 372376 520623 372808
rect 521278 372799 521291 372833
rect 521325 372799 521338 372833
rect 521278 372633 521338 372799
rect 521278 372599 521291 372633
rect 521325 372599 521338 372633
rect 521278 372376 521338 372599
rect 523158 374781 523298 374846
rect 523158 374747 523261 374781
rect 523295 374747 523298 374781
rect 523158 374741 523298 374747
rect 523158 374707 523171 374741
rect 523205 374707 523298 374741
rect 523158 374686 523298 374707
rect 523158 374341 523218 374686
rect 523158 374307 523171 374341
rect 523205 374307 523218 374341
rect 523158 373941 523218 374307
rect 523158 373907 523171 373941
rect 523205 373907 523218 373941
rect 523158 373546 523218 373907
rect 523338 374047 523378 374929
rect 524798 374505 524858 375387
rect 523419 374471 523439 374505
rect 523473 374471 523507 374505
rect 523545 374471 523575 374505
rect 523617 374471 523643 374505
rect 523689 374471 523711 374505
rect 523761 374471 523779 374505
rect 523833 374471 523847 374505
rect 523905 374471 523915 374505
rect 523977 374471 523983 374505
rect 524049 374471 524051 374505
rect 524085 374471 524087 374505
rect 524153 374471 524159 374505
rect 524221 374471 524231 374505
rect 524289 374471 524303 374505
rect 524357 374471 524375 374505
rect 524425 374471 524447 374505
rect 524493 374471 524519 374505
rect 524561 374471 524591 374505
rect 524629 374471 524663 374505
rect 524697 374471 524858 374505
rect 523338 374013 523439 374047
rect 523473 374013 523507 374047
rect 523545 374013 523575 374047
rect 523617 374013 523643 374047
rect 523689 374013 523711 374047
rect 523761 374013 523779 374047
rect 523833 374013 523847 374047
rect 523905 374013 523915 374047
rect 523977 374013 523983 374047
rect 524049 374013 524051 374047
rect 524085 374013 524087 374047
rect 524153 374013 524159 374047
rect 524221 374013 524231 374047
rect 524289 374013 524303 374047
rect 524357 374013 524375 374047
rect 524425 374013 524447 374047
rect 524493 374013 524519 374047
rect 524561 374013 524591 374047
rect 524629 374013 524663 374047
rect 524697 374013 524717 374047
rect 523158 373541 523298 373546
rect 523158 373507 523171 373541
rect 523205 373507 523298 373541
rect 523158 373481 523298 373507
rect 523158 373447 523261 373481
rect 523295 373447 523298 373481
rect 523158 373386 523298 373447
rect 523158 373141 523218 373386
rect 523158 373107 523171 373141
rect 523205 373107 523218 373141
rect 523158 372741 523218 373107
rect 523158 372707 523171 372741
rect 523205 372707 523218 372741
rect 513758 372187 513818 372353
rect 513758 372153 513771 372187
rect 513805 372153 513818 372187
rect 513758 371987 513818 372153
rect 523158 372341 523218 372707
rect 523158 372307 523171 372341
rect 523205 372307 523218 372341
rect 523158 372246 523218 372307
rect 523338 373131 523378 374013
rect 524798 373589 524858 374471
rect 523419 373555 523439 373589
rect 523473 373555 523507 373589
rect 523545 373555 523575 373589
rect 523617 373555 523643 373589
rect 523689 373555 523711 373589
rect 523761 373555 523779 373589
rect 523833 373555 523847 373589
rect 523905 373555 523915 373589
rect 523977 373555 523983 373589
rect 524049 373555 524051 373589
rect 524085 373555 524087 373589
rect 524153 373555 524159 373589
rect 524221 373555 524231 373589
rect 524289 373555 524303 373589
rect 524357 373555 524375 373589
rect 524425 373555 524447 373589
rect 524493 373555 524519 373589
rect 524561 373555 524591 373589
rect 524629 373555 524663 373589
rect 524697 373555 524858 373589
rect 523338 373097 523439 373131
rect 523473 373097 523507 373131
rect 523545 373097 523575 373131
rect 523617 373097 523643 373131
rect 523689 373097 523711 373131
rect 523761 373097 523779 373131
rect 523833 373097 523847 373131
rect 523905 373097 523915 373131
rect 523977 373097 523983 373131
rect 524049 373097 524051 373131
rect 524085 373097 524087 373131
rect 524153 373097 524159 373131
rect 524221 373097 524231 373131
rect 524289 373097 524303 373131
rect 524357 373097 524375 373131
rect 524425 373097 524447 373131
rect 524493 373097 524519 373131
rect 524561 373097 524591 373131
rect 524629 373097 524663 373131
rect 524697 373097 524717 373131
rect 523158 372181 523298 372246
rect 523158 372147 523261 372181
rect 523295 372147 523298 372181
rect 523158 372086 523298 372147
rect 523338 372215 523378 373097
rect 524798 372673 524858 373555
rect 523419 372639 523439 372673
rect 523473 372639 523507 372673
rect 523545 372639 523575 372673
rect 523617 372639 523643 372673
rect 523689 372639 523711 372673
rect 523761 372639 523779 372673
rect 523833 372639 523847 372673
rect 523905 372639 523915 372673
rect 523977 372639 523983 372673
rect 524049 372639 524051 372673
rect 524085 372639 524087 372673
rect 524153 372639 524159 372673
rect 524221 372639 524231 372673
rect 524289 372639 524303 372673
rect 524357 372639 524375 372673
rect 524425 372639 524447 372673
rect 524493 372639 524519 372673
rect 524561 372639 524591 372673
rect 524629 372639 524663 372673
rect 524697 372639 524858 372673
rect 523338 372181 523439 372215
rect 523473 372181 523507 372215
rect 523545 372181 523575 372215
rect 523617 372181 523643 372215
rect 523689 372181 523711 372215
rect 523761 372181 523779 372215
rect 523833 372181 523847 372215
rect 523905 372181 523915 372215
rect 523977 372181 523983 372215
rect 524049 372181 524051 372215
rect 524085 372181 524087 372215
rect 524153 372181 524159 372215
rect 524221 372181 524231 372215
rect 524289 372181 524303 372215
rect 524357 372181 524375 372215
rect 524425 372181 524447 372215
rect 524493 372181 524519 372215
rect 524561 372181 524591 372215
rect 524629 372181 524663 372215
rect 524697 372181 524717 372215
rect 513758 371953 513771 371987
rect 513805 371953 513818 371987
rect 513758 371787 513818 371953
rect 513758 371753 513771 371787
rect 513805 371753 513818 371787
rect 513758 371587 513818 371753
rect 513758 371553 513771 371587
rect 513805 371553 513818 371587
rect 513758 371387 513818 371553
rect 513758 371353 513771 371387
rect 513805 371353 513818 371387
rect 513758 371187 513818 371353
rect 513758 371153 513771 371187
rect 513805 371153 513818 371187
rect 513758 370987 513818 371153
rect 513758 370953 513771 370987
rect 513805 370953 513818 370987
rect 513758 370787 513818 370953
rect 513758 370753 513771 370787
rect 513805 370753 513818 370787
rect 513758 370587 513818 370753
rect 513758 370553 513771 370587
rect 513805 370553 513818 370587
rect 513758 370387 513818 370553
rect 513758 370353 513771 370387
rect 513805 370353 513818 370387
rect 513758 370187 513818 370353
rect 513758 370153 513771 370187
rect 513805 370153 513818 370187
rect 513758 369987 513818 370153
rect 513758 369953 513771 369987
rect 513805 369953 513818 369987
rect 513758 369787 513818 369953
rect 513758 369753 513771 369787
rect 513805 369753 513818 369787
rect 513758 369587 513818 369753
rect 515638 371889 515698 372072
rect 515638 371855 515651 371889
rect 515685 371855 515698 371889
rect 515638 371689 515698 371855
rect 515638 371655 515651 371689
rect 515685 371655 515698 371689
rect 515638 371489 515698 371655
rect 517518 371889 517578 372072
rect 517518 371855 517531 371889
rect 517565 371855 517578 371889
rect 517518 371689 517578 371855
rect 517518 371655 517531 371689
rect 517565 371655 517578 371689
rect 515638 371455 515651 371489
rect 515685 371455 515698 371489
rect 515638 371289 515698 371455
rect 515638 371255 515651 371289
rect 515685 371255 515698 371289
rect 515638 371089 515698 371255
rect 517518 371489 517578 371655
rect 517518 371455 517531 371489
rect 517565 371455 517578 371489
rect 517518 371289 517578 371455
rect 517518 371255 517531 371289
rect 517565 371255 517578 371289
rect 517518 371160 517578 371255
rect 515638 371055 515651 371089
rect 515685 371055 515698 371089
rect 515638 370889 515698 371055
rect 515638 370855 515651 370889
rect 515685 370855 515698 370889
rect 515638 370689 515698 370855
rect 515638 370655 515651 370689
rect 515685 370655 515698 370689
rect 515638 370489 515698 370655
rect 516578 371089 517578 371160
rect 516578 371073 517531 371089
rect 516578 370631 516617 371073
rect 516719 371055 517531 371073
rect 517565 371055 517578 371089
rect 516719 370889 517578 371055
rect 516719 370855 517531 370889
rect 517565 370855 517578 370889
rect 516719 370689 517578 370855
rect 516719 370655 517531 370689
rect 517565 370655 517578 370689
rect 516719 370631 517578 370655
rect 516578 370544 517578 370631
rect 515638 370455 515651 370489
rect 515685 370455 515698 370489
rect 515638 370289 515698 370455
rect 515638 370255 515651 370289
rect 515685 370255 515698 370289
rect 515638 370089 515698 370255
rect 515638 370055 515651 370089
rect 515685 370055 515698 370089
rect 517518 370489 517578 370544
rect 517518 370455 517531 370489
rect 517565 370455 517578 370489
rect 517518 370289 517578 370455
rect 517518 370255 517531 370289
rect 517565 370255 517578 370289
rect 517518 370089 517578 370255
rect 515638 369889 515698 370055
rect 515638 369855 515651 369889
rect 515685 369855 515698 369889
rect 515638 369632 515698 369855
rect 516473 369632 516863 370064
rect 517518 370055 517531 370089
rect 517565 370055 517578 370089
rect 517518 369889 517578 370055
rect 517518 369855 517531 369889
rect 517565 369855 517578 369889
rect 517518 369632 517578 369855
rect 523158 371941 523218 372086
rect 523158 371907 523171 371941
rect 523205 371907 523218 371941
rect 523158 371541 523218 371907
rect 523158 371507 523171 371541
rect 523205 371507 523218 371541
rect 523158 371141 523218 371507
rect 523158 371107 523171 371141
rect 523205 371107 523218 371141
rect 523158 370946 523218 371107
rect 523338 371299 523378 372181
rect 524798 371757 524858 372639
rect 523419 371723 523439 371757
rect 523473 371723 523507 371757
rect 523545 371723 523575 371757
rect 523617 371723 523643 371757
rect 523689 371723 523711 371757
rect 523761 371723 523779 371757
rect 523833 371723 523847 371757
rect 523905 371723 523915 371757
rect 523977 371723 523983 371757
rect 524049 371723 524051 371757
rect 524085 371723 524087 371757
rect 524153 371723 524159 371757
rect 524221 371723 524231 371757
rect 524289 371723 524303 371757
rect 524357 371723 524375 371757
rect 524425 371723 524447 371757
rect 524493 371723 524519 371757
rect 524561 371723 524591 371757
rect 524629 371723 524663 371757
rect 524697 371723 524858 371757
rect 523338 371265 523439 371299
rect 523473 371265 523507 371299
rect 523545 371265 523575 371299
rect 523617 371265 523643 371299
rect 523689 371265 523711 371299
rect 523761 371265 523779 371299
rect 523833 371265 523847 371299
rect 523905 371265 523915 371299
rect 523977 371265 523983 371299
rect 524049 371265 524051 371299
rect 524085 371265 524087 371299
rect 524153 371265 524159 371299
rect 524221 371265 524231 371299
rect 524289 371265 524303 371299
rect 524357 371265 524375 371299
rect 524425 371265 524447 371299
rect 524493 371265 524519 371299
rect 524561 371265 524591 371299
rect 524629 371265 524663 371299
rect 524697 371265 524717 371299
rect 523158 370881 523298 370946
rect 523158 370847 523261 370881
rect 523295 370847 523298 370881
rect 523158 370786 523298 370847
rect 523158 370741 523218 370786
rect 523158 370707 523171 370741
rect 523205 370707 523218 370741
rect 523158 370341 523218 370707
rect 523158 370307 523171 370341
rect 523205 370307 523218 370341
rect 523158 369941 523218 370307
rect 523158 369907 523171 369941
rect 523205 369907 523218 369941
rect 523158 369646 523218 369907
rect 523338 370383 523378 371265
rect 524798 370841 524858 371723
rect 523419 370807 523439 370841
rect 523473 370807 523507 370841
rect 523545 370807 523575 370841
rect 523617 370807 523643 370841
rect 523689 370807 523711 370841
rect 523761 370807 523779 370841
rect 523833 370807 523847 370841
rect 523905 370807 523915 370841
rect 523977 370807 523983 370841
rect 524049 370807 524051 370841
rect 524085 370807 524087 370841
rect 524153 370807 524159 370841
rect 524221 370807 524231 370841
rect 524289 370807 524303 370841
rect 524357 370807 524375 370841
rect 524425 370807 524447 370841
rect 524493 370807 524519 370841
rect 524561 370807 524591 370841
rect 524629 370807 524663 370841
rect 524697 370807 524858 370841
rect 523338 370349 523439 370383
rect 523473 370349 523507 370383
rect 523545 370349 523575 370383
rect 523617 370349 523643 370383
rect 523689 370349 523711 370383
rect 523761 370349 523779 370383
rect 523833 370349 523847 370383
rect 523905 370349 523915 370383
rect 523977 370349 523983 370383
rect 524049 370349 524051 370383
rect 524085 370349 524087 370383
rect 524153 370349 524159 370383
rect 524221 370349 524231 370383
rect 524289 370349 524303 370383
rect 524357 370349 524375 370383
rect 524425 370349 524447 370383
rect 524493 370349 524519 370383
rect 524561 370349 524591 370383
rect 524629 370349 524663 370383
rect 524697 370349 524717 370383
rect 513758 369553 513771 369587
rect 513805 369553 513818 369587
rect 513758 369387 513818 369553
rect 513758 369353 513771 369387
rect 513805 369353 513818 369387
rect 513758 369187 513818 369353
rect 523158 369581 523298 369646
rect 523158 369547 523261 369581
rect 523295 369547 523298 369581
rect 523158 369541 523298 369547
rect 523158 369507 523171 369541
rect 523205 369507 523298 369541
rect 523158 369486 523298 369507
rect 513758 369153 513771 369187
rect 513805 369153 513818 369187
rect 513758 368987 513818 369153
rect 513758 368953 513771 368987
rect 513805 368953 513818 368987
rect 513758 368787 513818 368953
rect 513758 368753 513771 368787
rect 513805 368753 513818 368787
rect 513758 368587 513818 368753
rect 513758 368553 513771 368587
rect 513805 368553 513818 368587
rect 513758 368387 513818 368553
rect 513758 368353 513771 368387
rect 513805 368353 513818 368387
rect 513758 368187 513818 368353
rect 513758 368153 513771 368187
rect 513805 368153 513818 368187
rect 513758 367987 513818 368153
rect 513758 367953 513771 367987
rect 513805 367953 513818 367987
rect 513758 367787 513818 367953
rect 513758 367753 513771 367787
rect 513805 367753 513818 367787
rect 513758 367587 513818 367753
rect 513758 367553 513771 367587
rect 513805 367553 513818 367587
rect 513758 367387 513818 367553
rect 513758 367353 513771 367387
rect 513805 367353 513818 367387
rect 513758 367187 513818 367353
rect 513758 367153 513771 367187
rect 513805 367153 513818 367187
rect 513758 366987 513818 367153
rect 513758 366953 513771 366987
rect 513805 366953 513818 366987
rect 513758 366787 513818 366953
rect 515638 369145 515698 369328
rect 515638 369111 515651 369145
rect 515685 369111 515698 369145
rect 515638 368945 515698 369111
rect 515638 368911 515651 368945
rect 515685 368911 515698 368945
rect 515638 368745 515698 368911
rect 517518 369145 517578 369328
rect 517518 369111 517531 369145
rect 517565 369111 517578 369145
rect 517518 368945 517578 369111
rect 517518 368911 517531 368945
rect 517565 368911 517578 368945
rect 515638 368711 515651 368745
rect 515685 368711 515698 368745
rect 515638 368545 515698 368711
rect 515638 368511 515651 368545
rect 515685 368511 515698 368545
rect 515638 368345 515698 368511
rect 517518 368745 517578 368911
rect 517518 368711 517531 368745
rect 517565 368711 517578 368745
rect 517518 368545 517578 368711
rect 517518 368511 517531 368545
rect 517565 368511 517578 368545
rect 517518 368416 517578 368511
rect 515638 368311 515651 368345
rect 515685 368311 515698 368345
rect 515638 368145 515698 368311
rect 515638 368111 515651 368145
rect 515685 368111 515698 368145
rect 515638 367945 515698 368111
rect 515638 367911 515651 367945
rect 515685 367911 515698 367945
rect 515638 367745 515698 367911
rect 516578 368345 517578 368416
rect 516578 368329 517531 368345
rect 516578 367887 516617 368329
rect 516719 368311 517531 368329
rect 517565 368311 517578 368345
rect 516719 368145 517578 368311
rect 516719 368111 517531 368145
rect 517565 368111 517578 368145
rect 516719 367945 517578 368111
rect 516719 367911 517531 367945
rect 517565 367911 517578 367945
rect 516719 367887 517578 367911
rect 516578 367800 517578 367887
rect 515638 367711 515651 367745
rect 515685 367711 515698 367745
rect 515638 367545 515698 367711
rect 515638 367511 515651 367545
rect 515685 367511 515698 367545
rect 515638 367345 515698 367511
rect 515638 367311 515651 367345
rect 515685 367311 515698 367345
rect 517518 367745 517578 367800
rect 517518 367711 517531 367745
rect 517565 367711 517578 367745
rect 517518 367545 517578 367711
rect 517518 367511 517531 367545
rect 517565 367511 517578 367545
rect 517518 367345 517578 367511
rect 515638 367145 515698 367311
rect 515638 367111 515651 367145
rect 515685 367111 515698 367145
rect 515638 366888 515698 367111
rect 516473 366888 516863 367320
rect 517518 367311 517531 367345
rect 517565 367311 517578 367345
rect 517518 367145 517578 367311
rect 517518 367111 517531 367145
rect 517565 367111 517578 367145
rect 517518 366888 517578 367111
rect 523158 369141 523218 369486
rect 523158 369107 523171 369141
rect 523205 369107 523218 369141
rect 523158 368741 523218 369107
rect 523158 368707 523171 368741
rect 523205 368707 523218 368741
rect 523158 368346 523218 368707
rect 523338 369467 523378 370349
rect 524798 369925 524858 370807
rect 523419 369891 523439 369925
rect 523473 369891 523507 369925
rect 523545 369891 523575 369925
rect 523617 369891 523643 369925
rect 523689 369891 523711 369925
rect 523761 369891 523779 369925
rect 523833 369891 523847 369925
rect 523905 369891 523915 369925
rect 523977 369891 523983 369925
rect 524049 369891 524051 369925
rect 524085 369891 524087 369925
rect 524153 369891 524159 369925
rect 524221 369891 524231 369925
rect 524289 369891 524303 369925
rect 524357 369891 524375 369925
rect 524425 369891 524447 369925
rect 524493 369891 524519 369925
rect 524561 369891 524591 369925
rect 524629 369891 524663 369925
rect 524697 369891 524858 369925
rect 523338 369433 523439 369467
rect 523473 369433 523507 369467
rect 523545 369433 523575 369467
rect 523617 369433 523643 369467
rect 523689 369433 523711 369467
rect 523761 369433 523779 369467
rect 523833 369433 523847 369467
rect 523905 369433 523915 369467
rect 523977 369433 523983 369467
rect 524049 369433 524051 369467
rect 524085 369433 524087 369467
rect 524153 369433 524159 369467
rect 524221 369433 524231 369467
rect 524289 369433 524303 369467
rect 524357 369433 524375 369467
rect 524425 369433 524447 369467
rect 524493 369433 524519 369467
rect 524561 369433 524591 369467
rect 524629 369433 524663 369467
rect 524697 369433 524717 369467
rect 523338 368551 523378 369433
rect 524798 369009 524858 369891
rect 523419 368975 523439 369009
rect 523473 368975 523507 369009
rect 523545 368975 523575 369009
rect 523617 368975 523643 369009
rect 523689 368975 523711 369009
rect 523761 368975 523779 369009
rect 523833 368975 523847 369009
rect 523905 368975 523915 369009
rect 523977 368975 523983 369009
rect 524049 368975 524051 369009
rect 524085 368975 524087 369009
rect 524153 368975 524159 369009
rect 524221 368975 524231 369009
rect 524289 368975 524303 369009
rect 524357 368975 524375 369009
rect 524425 368975 524447 369009
rect 524493 368975 524519 369009
rect 524561 368975 524591 369009
rect 524629 368975 524663 369009
rect 524697 368975 524858 369009
rect 523338 368517 523439 368551
rect 523473 368517 523507 368551
rect 523545 368517 523575 368551
rect 523617 368517 523643 368551
rect 523689 368517 523711 368551
rect 523761 368517 523779 368551
rect 523833 368517 523847 368551
rect 523905 368517 523915 368551
rect 523977 368517 523983 368551
rect 524049 368517 524051 368551
rect 524085 368517 524087 368551
rect 524153 368517 524159 368551
rect 524221 368517 524231 368551
rect 524289 368517 524303 368551
rect 524357 368517 524375 368551
rect 524425 368517 524447 368551
rect 524493 368517 524519 368551
rect 524561 368517 524591 368551
rect 524629 368517 524663 368551
rect 524697 368517 524717 368551
rect 523158 368341 523298 368346
rect 523158 368307 523171 368341
rect 523205 368307 523298 368341
rect 523158 368281 523298 368307
rect 523158 368247 523261 368281
rect 523295 368247 523298 368281
rect 523158 368186 523298 368247
rect 523158 367941 523218 368186
rect 523158 367907 523171 367941
rect 523205 367907 523218 367941
rect 523158 367541 523218 367907
rect 523158 367507 523171 367541
rect 523205 367507 523218 367541
rect 523158 367141 523218 367507
rect 523158 367107 523171 367141
rect 523205 367107 523218 367141
rect 523158 367046 523218 367107
rect 523338 367635 523378 368517
rect 524798 368093 524858 368975
rect 523419 368059 523439 368093
rect 523473 368059 523507 368093
rect 523545 368059 523575 368093
rect 523617 368059 523643 368093
rect 523689 368059 523711 368093
rect 523761 368059 523779 368093
rect 523833 368059 523847 368093
rect 523905 368059 523915 368093
rect 523977 368059 523983 368093
rect 524049 368059 524051 368093
rect 524085 368059 524087 368093
rect 524153 368059 524159 368093
rect 524221 368059 524231 368093
rect 524289 368059 524303 368093
rect 524357 368059 524375 368093
rect 524425 368059 524447 368093
rect 524493 368059 524519 368093
rect 524561 368059 524591 368093
rect 524629 368059 524663 368093
rect 524697 368059 524858 368093
rect 523338 367601 523439 367635
rect 523473 367601 523507 367635
rect 523545 367601 523575 367635
rect 523617 367601 523643 367635
rect 523689 367601 523711 367635
rect 523761 367601 523779 367635
rect 523833 367601 523847 367635
rect 523905 367601 523915 367635
rect 523977 367601 523983 367635
rect 524049 367601 524051 367635
rect 524085 367601 524087 367635
rect 524153 367601 524159 367635
rect 524221 367601 524231 367635
rect 524289 367601 524303 367635
rect 524357 367601 524375 367635
rect 524425 367601 524447 367635
rect 524493 367601 524519 367635
rect 524561 367601 524591 367635
rect 524629 367601 524663 367635
rect 524697 367601 524717 367635
rect 523158 366981 523298 367046
rect 523158 366947 523261 366981
rect 523295 366947 523298 366981
rect 513758 366753 513771 366787
rect 513805 366753 513818 366787
rect 513758 366587 513818 366753
rect 513758 366553 513771 366587
rect 513805 366553 513818 366587
rect 523158 366886 523298 366947
rect 523158 366741 523218 366886
rect 523158 366707 523171 366741
rect 523205 366707 523218 366741
rect 513758 366387 513818 366553
rect 513758 366353 513771 366387
rect 513805 366353 513818 366387
rect 513758 366187 513818 366353
rect 513758 366153 513771 366187
rect 513805 366153 513818 366187
rect 513758 365987 513818 366153
rect 513758 365953 513771 365987
rect 513805 365953 513818 365987
rect 513758 365787 513818 365953
rect 513758 365753 513771 365787
rect 513805 365753 513818 365787
rect 513758 365587 513818 365753
rect 513758 365553 513771 365587
rect 513805 365553 513818 365587
rect 513758 365387 513818 365553
rect 513758 365353 513771 365387
rect 513805 365353 513818 365387
rect 513758 365187 513818 365353
rect 513758 365153 513771 365187
rect 513805 365153 513818 365187
rect 513758 364987 513818 365153
rect 513758 364953 513771 364987
rect 513805 364953 513818 364987
rect 513758 364787 513818 364953
rect 513758 364753 513771 364787
rect 513805 364753 513818 364787
rect 513758 364587 513818 364753
rect 513758 364553 513771 364587
rect 513805 364553 513818 364587
rect 513758 364387 513818 364553
rect 513758 364353 513771 364387
rect 513805 364353 513818 364387
rect 513758 364187 513818 364353
rect 513758 364153 513771 364187
rect 513805 364153 513818 364187
rect 513758 363987 513818 364153
rect 515638 366401 515698 366584
rect 515638 366367 515651 366401
rect 515685 366367 515698 366401
rect 515638 366201 515698 366367
rect 515638 366167 515651 366201
rect 515685 366167 515698 366201
rect 515638 366001 515698 366167
rect 517518 366401 517578 366584
rect 517518 366367 517531 366401
rect 517565 366367 517578 366401
rect 517518 366201 517578 366367
rect 517518 366167 517531 366201
rect 517565 366167 517578 366201
rect 515638 365967 515651 366001
rect 515685 365967 515698 366001
rect 515638 365801 515698 365967
rect 515638 365767 515651 365801
rect 515685 365767 515698 365801
rect 515638 365601 515698 365767
rect 517518 366001 517578 366167
rect 517518 365967 517531 366001
rect 517565 365967 517578 366001
rect 517518 365801 517578 365967
rect 517518 365767 517531 365801
rect 517565 365767 517578 365801
rect 517518 365672 517578 365767
rect 515638 365567 515651 365601
rect 515685 365567 515698 365601
rect 515638 365401 515698 365567
rect 515638 365367 515651 365401
rect 515685 365367 515698 365401
rect 515638 365201 515698 365367
rect 515638 365167 515651 365201
rect 515685 365167 515698 365201
rect 515638 365001 515698 365167
rect 516578 365601 517578 365672
rect 516578 365585 517531 365601
rect 516578 365143 516617 365585
rect 516719 365567 517531 365585
rect 517565 365567 517578 365601
rect 516719 365401 517578 365567
rect 516719 365367 517531 365401
rect 517565 365367 517578 365401
rect 516719 365201 517578 365367
rect 516719 365167 517531 365201
rect 517565 365167 517578 365201
rect 516719 365143 517578 365167
rect 516578 365056 517578 365143
rect 515638 364967 515651 365001
rect 515685 364967 515698 365001
rect 515638 364801 515698 364967
rect 515638 364767 515651 364801
rect 515685 364767 515698 364801
rect 515638 364601 515698 364767
rect 515638 364567 515651 364601
rect 515685 364567 515698 364601
rect 517518 365001 517578 365056
rect 517518 364967 517531 365001
rect 517565 364967 517578 365001
rect 517518 364801 517578 364967
rect 517518 364767 517531 364801
rect 517565 364767 517578 364801
rect 517518 364601 517578 364767
rect 515638 364401 515698 364567
rect 515638 364367 515651 364401
rect 515685 364367 515698 364401
rect 515638 364144 515698 364367
rect 516473 364144 516863 364576
rect 517518 364567 517531 364601
rect 517565 364567 517578 364601
rect 517518 364401 517578 364567
rect 517518 364367 517531 364401
rect 517565 364367 517578 364401
rect 517518 364144 517578 364367
rect 519398 366401 519458 366584
rect 519398 366367 519411 366401
rect 519445 366367 519458 366401
rect 519398 366201 519458 366367
rect 519398 366167 519411 366201
rect 519445 366167 519458 366201
rect 519398 366001 519458 366167
rect 521278 366401 521338 366584
rect 521278 366367 521291 366401
rect 521325 366367 521338 366401
rect 521278 366201 521338 366367
rect 521278 366167 521291 366201
rect 521325 366167 521338 366201
rect 519398 365967 519411 366001
rect 519445 365967 519458 366001
rect 519398 365801 519458 365967
rect 519398 365767 519411 365801
rect 519445 365767 519458 365801
rect 519398 365601 519458 365767
rect 521278 366001 521338 366167
rect 521278 365967 521291 366001
rect 521325 365967 521338 366001
rect 521278 365801 521338 365967
rect 521278 365767 521291 365801
rect 521325 365767 521338 365801
rect 521278 365672 521338 365767
rect 519398 365567 519411 365601
rect 519445 365567 519458 365601
rect 519398 365401 519458 365567
rect 519398 365367 519411 365401
rect 519445 365367 519458 365401
rect 519398 365201 519458 365367
rect 519398 365167 519411 365201
rect 519445 365167 519458 365201
rect 519398 365001 519458 365167
rect 520338 365601 521338 365672
rect 520338 365585 521291 365601
rect 520338 365143 520377 365585
rect 520479 365567 521291 365585
rect 521325 365567 521338 365601
rect 520479 365401 521338 365567
rect 520479 365367 521291 365401
rect 521325 365367 521338 365401
rect 520479 365201 521338 365367
rect 520479 365167 521291 365201
rect 521325 365167 521338 365201
rect 520479 365143 521338 365167
rect 520338 365056 521338 365143
rect 519398 364967 519411 365001
rect 519445 364967 519458 365001
rect 519398 364801 519458 364967
rect 519398 364767 519411 364801
rect 519445 364767 519458 364801
rect 519398 364601 519458 364767
rect 519398 364567 519411 364601
rect 519445 364567 519458 364601
rect 521278 365001 521338 365056
rect 521278 364967 521291 365001
rect 521325 364967 521338 365001
rect 521278 364801 521338 364967
rect 521278 364767 521291 364801
rect 521325 364767 521338 364801
rect 521278 364601 521338 364767
rect 519398 364401 519458 364567
rect 519398 364367 519411 364401
rect 519445 364367 519458 364401
rect 519398 364144 519458 364367
rect 520233 364144 520623 364576
rect 521278 364567 521291 364601
rect 521325 364567 521338 364601
rect 521278 364401 521338 364567
rect 521278 364367 521291 364401
rect 521325 364367 521338 364401
rect 521278 364144 521338 364367
rect 523158 366341 523218 366707
rect 523158 366307 523171 366341
rect 523205 366307 523218 366341
rect 523158 365941 523218 366307
rect 523158 365907 523171 365941
rect 523205 365907 523218 365941
rect 523158 365746 523218 365907
rect 523338 366719 523378 367601
rect 524798 367177 524858 368059
rect 523419 367143 523439 367177
rect 523473 367143 523507 367177
rect 523545 367143 523575 367177
rect 523617 367143 523643 367177
rect 523689 367143 523711 367177
rect 523761 367143 523779 367177
rect 523833 367143 523847 367177
rect 523905 367143 523915 367177
rect 523977 367143 523983 367177
rect 524049 367143 524051 367177
rect 524085 367143 524087 367177
rect 524153 367143 524159 367177
rect 524221 367143 524231 367177
rect 524289 367143 524303 367177
rect 524357 367143 524375 367177
rect 524425 367143 524447 367177
rect 524493 367143 524519 367177
rect 524561 367143 524591 367177
rect 524629 367143 524663 367177
rect 524697 367143 524858 367177
rect 523338 366685 523439 366719
rect 523473 366685 523507 366719
rect 523545 366685 523575 366719
rect 523617 366685 523643 366719
rect 523689 366685 523711 366719
rect 523761 366685 523779 366719
rect 523833 366685 523847 366719
rect 523905 366685 523915 366719
rect 523977 366685 523983 366719
rect 524049 366685 524051 366719
rect 524085 366685 524087 366719
rect 524153 366685 524159 366719
rect 524221 366685 524231 366719
rect 524289 366685 524303 366719
rect 524357 366685 524375 366719
rect 524425 366685 524447 366719
rect 524493 366685 524519 366719
rect 524561 366685 524591 366719
rect 524629 366685 524663 366719
rect 524697 366685 524717 366719
rect 523338 365803 523378 366685
rect 524798 366261 524858 367143
rect 523419 366227 523439 366261
rect 523473 366227 523507 366261
rect 523545 366227 523575 366261
rect 523617 366227 523643 366261
rect 523689 366227 523711 366261
rect 523761 366227 523779 366261
rect 523833 366227 523847 366261
rect 523905 366227 523915 366261
rect 523977 366227 523983 366261
rect 524049 366227 524051 366261
rect 524085 366227 524087 366261
rect 524153 366227 524159 366261
rect 524221 366227 524231 366261
rect 524289 366227 524303 366261
rect 524357 366227 524375 366261
rect 524425 366227 524447 366261
rect 524493 366227 524519 366261
rect 524561 366227 524591 366261
rect 524629 366227 524663 366261
rect 524697 366227 524858 366261
rect 523338 365769 523439 365803
rect 523473 365769 523507 365803
rect 523545 365769 523575 365803
rect 523617 365769 523643 365803
rect 523689 365769 523711 365803
rect 523761 365769 523779 365803
rect 523833 365769 523847 365803
rect 523905 365769 523915 365803
rect 523977 365769 523983 365803
rect 524049 365769 524051 365803
rect 524085 365769 524087 365803
rect 524153 365769 524159 365803
rect 524221 365769 524231 365803
rect 524289 365769 524303 365803
rect 524357 365769 524375 365803
rect 524425 365769 524447 365803
rect 524493 365769 524519 365803
rect 524561 365769 524591 365803
rect 524629 365769 524663 365803
rect 524697 365769 524717 365803
rect 523158 365681 523298 365746
rect 523158 365647 523261 365681
rect 523295 365647 523298 365681
rect 523158 365586 523298 365647
rect 523158 365541 523218 365586
rect 523158 365507 523171 365541
rect 523205 365507 523218 365541
rect 523158 365141 523218 365507
rect 523158 365107 523171 365141
rect 523205 365107 523218 365141
rect 523158 364741 523218 365107
rect 523158 364707 523171 364741
rect 523205 364707 523218 364741
rect 523158 364446 523218 364707
rect 523338 364887 523378 365769
rect 524798 365345 524858 366227
rect 523419 365311 523439 365345
rect 523473 365311 523507 365345
rect 523545 365311 523575 365345
rect 523617 365311 523643 365345
rect 523689 365311 523711 365345
rect 523761 365311 523779 365345
rect 523833 365311 523847 365345
rect 523905 365311 523915 365345
rect 523977 365311 523983 365345
rect 524049 365311 524051 365345
rect 524085 365311 524087 365345
rect 524153 365311 524159 365345
rect 524221 365311 524231 365345
rect 524289 365311 524303 365345
rect 524357 365311 524375 365345
rect 524425 365311 524447 365345
rect 524493 365311 524519 365345
rect 524561 365311 524591 365345
rect 524629 365311 524663 365345
rect 524697 365311 524858 365345
rect 523338 364853 523439 364887
rect 523473 364853 523507 364887
rect 523545 364853 523575 364887
rect 523617 364853 523643 364887
rect 523689 364853 523711 364887
rect 523761 364853 523779 364887
rect 523833 364853 523847 364887
rect 523905 364853 523915 364887
rect 523977 364853 523983 364887
rect 524049 364853 524051 364887
rect 524085 364853 524087 364887
rect 524153 364853 524159 364887
rect 524221 364853 524231 364887
rect 524289 364853 524303 364887
rect 524357 364853 524375 364887
rect 524425 364853 524447 364887
rect 524493 364853 524519 364887
rect 524561 364853 524591 364887
rect 524629 364853 524663 364887
rect 524697 364853 524717 364887
rect 523158 364381 523298 364446
rect 523158 364347 523261 364381
rect 523295 364347 523298 364381
rect 523158 364341 523298 364347
rect 523158 364307 523171 364341
rect 523205 364307 523298 364341
rect 523158 364286 523298 364307
rect 513758 363953 513771 363987
rect 513805 363953 513818 363987
rect 513758 363787 513818 363953
rect 513758 363753 513771 363787
rect 513805 363753 513818 363787
rect 513758 363587 513818 363753
rect 513758 363553 513771 363587
rect 513805 363553 513818 363587
rect 513758 363387 513818 363553
rect 513758 363353 513771 363387
rect 513805 363353 513818 363387
rect 513758 363187 513818 363353
rect 513758 363153 513771 363187
rect 513805 363153 513818 363187
rect 513758 362987 513818 363153
rect 513758 362953 513771 362987
rect 513805 362953 513818 362987
rect 513758 362787 513818 362953
rect 513758 362753 513771 362787
rect 513805 362753 513818 362787
rect 513758 362587 513818 362753
rect 513758 362553 513771 362587
rect 513805 362553 513818 362587
rect 513758 362450 513818 362553
rect 523158 363941 523218 364286
rect 523158 363907 523171 363941
rect 523205 363907 523218 363941
rect 523158 363541 523218 363907
rect 523158 363507 523171 363541
rect 523205 363507 523218 363541
rect 523158 363141 523218 363507
rect 523158 363107 523171 363141
rect 523205 363107 523218 363141
rect 523158 362741 523218 363107
rect 523158 362707 523171 362741
rect 523205 362707 523218 362741
rect 523158 362516 523218 362707
rect 523338 363971 523378 364853
rect 524798 364429 524858 365311
rect 523419 364395 523439 364429
rect 523473 364395 523507 364429
rect 523545 364395 523575 364429
rect 523617 364395 523643 364429
rect 523689 364395 523711 364429
rect 523761 364395 523779 364429
rect 523833 364395 523847 364429
rect 523905 364395 523915 364429
rect 523977 364395 523983 364429
rect 524049 364395 524051 364429
rect 524085 364395 524087 364429
rect 524153 364395 524159 364429
rect 524221 364395 524231 364429
rect 524289 364395 524303 364429
rect 524357 364395 524375 364429
rect 524425 364395 524447 364429
rect 524493 364395 524519 364429
rect 524561 364395 524591 364429
rect 524629 364395 524663 364429
rect 524697 364395 524858 364429
rect 523338 363937 523439 363971
rect 523473 363937 523507 363971
rect 523545 363937 523575 363971
rect 523617 363937 523643 363971
rect 523689 363937 523711 363971
rect 523761 363937 523779 363971
rect 523833 363937 523847 363971
rect 523905 363937 523915 363971
rect 523977 363937 523983 363971
rect 524049 363937 524051 363971
rect 524085 363937 524087 363971
rect 524153 363937 524159 363971
rect 524221 363937 524231 363971
rect 524289 363937 524303 363971
rect 524357 363937 524375 363971
rect 524425 363937 524447 363971
rect 524493 363937 524519 363971
rect 524561 363937 524591 363971
rect 524629 363937 524663 363971
rect 524697 363937 524717 363971
rect 523338 363055 523378 363937
rect 524798 363513 524858 364395
rect 523419 363479 523439 363513
rect 523473 363479 523507 363513
rect 523545 363479 523575 363513
rect 523617 363479 523643 363513
rect 523689 363479 523711 363513
rect 523761 363479 523779 363513
rect 523833 363479 523847 363513
rect 523905 363479 523915 363513
rect 523977 363479 523983 363513
rect 524049 363479 524051 363513
rect 524085 363479 524087 363513
rect 524153 363479 524159 363513
rect 524221 363479 524231 363513
rect 524289 363479 524303 363513
rect 524357 363479 524375 363513
rect 524425 363479 524447 363513
rect 524493 363479 524519 363513
rect 524561 363479 524591 363513
rect 524629 363479 524663 363513
rect 524697 363479 524858 363513
rect 523338 363021 523439 363055
rect 523473 363021 523507 363055
rect 523545 363021 523575 363055
rect 523617 363021 523643 363055
rect 523689 363021 523711 363055
rect 523761 363021 523779 363055
rect 523833 363021 523847 363055
rect 523905 363021 523915 363055
rect 523977 363021 523983 363055
rect 524049 363021 524051 363055
rect 524085 363021 524087 363055
rect 524153 363021 524159 363055
rect 524221 363021 524231 363055
rect 524289 363021 524303 363055
rect 524357 363021 524375 363055
rect 524425 363021 524447 363055
rect 524493 363021 524519 363055
rect 524561 363021 524591 363055
rect 524629 363021 524663 363055
rect 524697 363021 524717 363055
rect 523338 362516 523378 363021
rect 524798 362597 524858 363479
rect 523419 362563 523439 362597
rect 523473 362563 523507 362597
rect 523545 362563 523575 362597
rect 523617 362563 523643 362597
rect 523689 362563 523711 362597
rect 523761 362563 523779 362597
rect 523833 362563 523847 362597
rect 523905 362563 523915 362597
rect 523977 362563 523983 362597
rect 524049 362563 524051 362597
rect 524085 362563 524087 362597
rect 524153 362563 524159 362597
rect 524221 362563 524231 362597
rect 524289 362563 524303 362597
rect 524357 362563 524375 362597
rect 524425 362563 524447 362597
rect 524493 362563 524519 362597
rect 524561 362563 524591 362597
rect 524629 362563 524663 362597
rect 524697 362563 524858 362597
rect 524798 362516 524858 362563
rect 524904 389941 524964 390124
rect 524904 389907 524917 389941
rect 524951 389907 524964 389941
rect 524904 389541 524964 389907
rect 524904 389533 524917 389541
rect 524904 389499 524907 389533
rect 524951 389507 524964 389541
rect 524941 389499 524964 389507
rect 524904 389141 524964 389499
rect 524904 389107 524917 389141
rect 524951 389107 524964 389141
rect 524904 388741 524964 389107
rect 524904 388707 524917 388741
rect 524951 388707 524964 388741
rect 524904 388341 524964 388707
rect 524904 388307 524917 388341
rect 524951 388307 524964 388341
rect 524904 387941 524964 388307
rect 524904 387907 524917 387941
rect 524951 387907 524964 387941
rect 524904 387541 524964 387907
rect 524904 387507 524917 387541
rect 524951 387507 524964 387541
rect 524904 387141 524964 387507
rect 524904 387107 524917 387141
rect 524951 387107 524964 387141
rect 524904 386741 524964 387107
rect 524904 386707 524917 386741
rect 524951 386707 524964 386741
rect 524904 386341 524964 386707
rect 524904 386307 524917 386341
rect 524951 386307 524964 386341
rect 524904 385941 524964 386307
rect 524904 385907 524917 385941
rect 524951 385907 524964 385941
rect 524904 385541 524964 385907
rect 524904 385507 524917 385541
rect 524951 385507 524964 385541
rect 524904 385141 524964 385507
rect 524904 385107 524917 385141
rect 524951 385107 524964 385141
rect 524904 384741 524964 385107
rect 524904 384707 524917 384741
rect 524951 384707 524964 384741
rect 524904 384341 524964 384707
rect 524904 384307 524917 384341
rect 524951 384307 524964 384341
rect 524904 383941 524964 384307
rect 524904 383907 524917 383941
rect 524951 383907 524964 383941
rect 524904 383541 524964 383907
rect 524904 383507 524917 383541
rect 524951 383507 524964 383541
rect 524904 383141 524964 383507
rect 524904 383107 524917 383141
rect 524951 383107 524964 383141
rect 524904 382741 524964 383107
rect 524904 382707 524917 382741
rect 524951 382707 524964 382741
rect 524904 382341 524964 382707
rect 524904 382307 524917 382341
rect 524951 382307 524964 382341
rect 524904 381941 524964 382307
rect 524904 381907 524917 381941
rect 524951 381907 524964 381941
rect 524904 381541 524964 381907
rect 524904 381507 524917 381541
rect 524951 381507 524964 381541
rect 524904 381141 524964 381507
rect 524904 381107 524917 381141
rect 524951 381107 524964 381141
rect 524904 380741 524964 381107
rect 524904 380707 524917 380741
rect 524951 380707 524964 380741
rect 524904 380341 524964 380707
rect 524904 380307 524917 380341
rect 524951 380307 524964 380341
rect 524904 379941 524964 380307
rect 524904 379907 524917 379941
rect 524951 379907 524964 379941
rect 524904 379541 524964 379907
rect 524904 379507 524917 379541
rect 524951 379507 524964 379541
rect 524904 379141 524964 379507
rect 524904 379107 524917 379141
rect 524951 379107 524964 379141
rect 524904 378741 524964 379107
rect 524904 378707 524917 378741
rect 524951 378707 524964 378741
rect 524904 378341 524964 378707
rect 524904 378307 524917 378341
rect 524951 378307 524964 378341
rect 524904 377941 524964 378307
rect 524904 377907 524917 377941
rect 524951 377907 524964 377941
rect 524904 377541 524964 377907
rect 524904 377507 524917 377541
rect 524951 377507 524964 377541
rect 524904 377141 524964 377507
rect 524904 377107 524917 377141
rect 524951 377107 524964 377141
rect 524904 376741 524964 377107
rect 524904 376707 524917 376741
rect 524951 376707 524964 376741
rect 524904 376341 524964 376707
rect 524904 376307 524917 376341
rect 524951 376307 524964 376341
rect 524904 375941 524964 376307
rect 524904 375907 524917 375941
rect 524951 375907 524964 375941
rect 524904 375541 524964 375907
rect 524904 375507 524917 375541
rect 524951 375507 524964 375541
rect 524904 375141 524964 375507
rect 524904 375107 524917 375141
rect 524951 375107 524964 375141
rect 524904 374741 524964 375107
rect 524904 374707 524917 374741
rect 524951 374707 524964 374741
rect 524904 374341 524964 374707
rect 524904 374307 524917 374341
rect 524951 374307 524964 374341
rect 524904 373941 524964 374307
rect 524904 373907 524917 373941
rect 524951 373907 524964 373941
rect 524904 373541 524964 373907
rect 524904 373507 524917 373541
rect 524951 373507 524964 373541
rect 524904 373141 524964 373507
rect 524904 373107 524917 373141
rect 524951 373107 524964 373141
rect 524904 372741 524964 373107
rect 524904 372707 524917 372741
rect 524951 372707 524964 372741
rect 524904 372341 524964 372707
rect 524904 372307 524917 372341
rect 524951 372307 524964 372341
rect 524904 371941 524964 372307
rect 524904 371907 524917 371941
rect 524951 371907 524964 371941
rect 524904 371541 524964 371907
rect 524904 371507 524917 371541
rect 524951 371507 524964 371541
rect 524904 371141 524964 371507
rect 524904 371107 524917 371141
rect 524951 371107 524964 371141
rect 524904 370741 524964 371107
rect 524904 370707 524917 370741
rect 524951 370707 524964 370741
rect 524904 370341 524964 370707
rect 524904 370307 524917 370341
rect 524951 370307 524964 370341
rect 524904 369941 524964 370307
rect 524904 369907 524917 369941
rect 524951 369907 524964 369941
rect 524904 369541 524964 369907
rect 524904 369507 524917 369541
rect 524951 369507 524964 369541
rect 524904 369141 524964 369507
rect 524904 369107 524917 369141
rect 524951 369107 524964 369141
rect 524904 368741 524964 369107
rect 524904 368707 524917 368741
rect 524951 368707 524964 368741
rect 524904 368341 524964 368707
rect 524904 368307 524917 368341
rect 524951 368307 524964 368341
rect 524904 367941 524964 368307
rect 524904 367907 524917 367941
rect 524951 367907 524964 367941
rect 524904 367541 524964 367907
rect 524904 367507 524917 367541
rect 524951 367507 524964 367541
rect 524904 367141 524964 367507
rect 524904 367107 524917 367141
rect 524951 367107 524964 367141
rect 524904 366741 524964 367107
rect 524904 366707 524917 366741
rect 524951 366707 524964 366741
rect 524904 366341 524964 366707
rect 524904 366307 524917 366341
rect 524951 366307 524964 366341
rect 524904 365941 524964 366307
rect 524904 365907 524917 365941
rect 524951 365907 524964 365941
rect 524904 365541 524964 365907
rect 524904 365507 524917 365541
rect 524951 365507 524964 365541
rect 524904 365141 524964 365507
rect 524904 365107 524917 365141
rect 524951 365107 524964 365141
rect 524904 364741 524964 365107
rect 524904 364707 524917 364741
rect 524951 364707 524964 364741
rect 524904 364341 524964 364707
rect 524904 364307 524917 364341
rect 524951 364307 524964 364341
rect 524904 363941 524964 364307
rect 524904 363907 524917 363941
rect 524951 363907 524964 363941
rect 524904 363541 524964 363907
rect 524904 363507 524917 363541
rect 524951 363507 524964 363541
rect 524904 363141 524964 363507
rect 524904 363107 524917 363141
rect 524951 363107 524964 363141
rect 524904 362741 524964 363107
rect 524904 362707 524917 362741
rect 524951 362707 524964 362741
rect 524904 362516 524964 362707
rect 525038 389941 525098 390222
rect 525038 389907 525051 389941
rect 525085 389907 525098 389941
rect 525038 389541 525098 389907
rect 525038 389507 525051 389541
rect 525085 389507 525098 389541
rect 525038 389141 525098 389507
rect 525038 389107 525051 389141
rect 525085 389107 525098 389141
rect 525038 388741 525098 389107
rect 525038 388707 525051 388741
rect 525085 388707 525098 388741
rect 525038 388341 525098 388707
rect 525038 388307 525051 388341
rect 525085 388307 525098 388341
rect 525038 387941 525098 388307
rect 525038 387907 525051 387941
rect 525085 387907 525098 387941
rect 525038 387541 525098 387907
rect 525038 387507 525051 387541
rect 525085 387507 525098 387541
rect 525038 387141 525098 387507
rect 525038 387107 525051 387141
rect 525085 387107 525098 387141
rect 525038 386741 525098 387107
rect 525038 386707 525051 386741
rect 525085 386707 525098 386741
rect 525038 386341 525098 386707
rect 525038 386307 525051 386341
rect 525085 386307 525098 386341
rect 525038 385941 525098 386307
rect 525038 385907 525051 385941
rect 525085 385907 525098 385941
rect 525038 385541 525098 385907
rect 525038 385507 525051 385541
rect 525085 385507 525098 385541
rect 525038 385141 525098 385507
rect 525038 385107 525051 385141
rect 525085 385107 525098 385141
rect 525038 384741 525098 385107
rect 525038 384707 525051 384741
rect 525085 384707 525098 384741
rect 525038 384341 525098 384707
rect 525038 384307 525051 384341
rect 525085 384307 525098 384341
rect 525038 383941 525098 384307
rect 525038 383907 525051 383941
rect 525085 383907 525098 383941
rect 525038 383541 525098 383907
rect 525038 383507 525051 383541
rect 525085 383507 525098 383541
rect 525038 383141 525098 383507
rect 525038 383107 525051 383141
rect 525085 383107 525098 383141
rect 525038 382741 525098 383107
rect 525038 382707 525051 382741
rect 525085 382707 525098 382741
rect 525038 382341 525098 382707
rect 525038 382307 525051 382341
rect 525085 382307 525098 382341
rect 525038 381941 525098 382307
rect 525038 381907 525051 381941
rect 525085 381907 525098 381941
rect 525038 381541 525098 381907
rect 525038 381507 525051 381541
rect 525085 381507 525098 381541
rect 525038 381141 525098 381507
rect 525038 381107 525051 381141
rect 525085 381107 525098 381141
rect 525038 380741 525098 381107
rect 525038 380707 525051 380741
rect 525085 380707 525098 380741
rect 525038 380341 525098 380707
rect 525038 380307 525051 380341
rect 525085 380307 525098 380341
rect 525038 379941 525098 380307
rect 525038 379907 525051 379941
rect 525085 379907 525098 379941
rect 525038 379541 525098 379907
rect 525038 379507 525051 379541
rect 525085 379507 525098 379541
rect 525038 379141 525098 379507
rect 525038 379107 525051 379141
rect 525085 379107 525098 379141
rect 525038 378741 525098 379107
rect 525038 378707 525051 378741
rect 525085 378707 525098 378741
rect 525038 378341 525098 378707
rect 525038 378307 525051 378341
rect 525085 378307 525098 378341
rect 525038 377941 525098 378307
rect 525038 377907 525051 377941
rect 525085 377907 525098 377941
rect 525038 377541 525098 377907
rect 525038 377507 525051 377541
rect 525085 377507 525098 377541
rect 525038 377141 525098 377507
rect 525038 377107 525051 377141
rect 525085 377107 525098 377141
rect 525038 376741 525098 377107
rect 525038 376707 525051 376741
rect 525085 376707 525098 376741
rect 525038 376341 525098 376707
rect 525038 376307 525051 376341
rect 525085 376307 525098 376341
rect 525038 375941 525098 376307
rect 525038 375907 525051 375941
rect 525085 375907 525098 375941
rect 525038 375541 525098 375907
rect 525038 375507 525051 375541
rect 525085 375507 525098 375541
rect 525038 375141 525098 375507
rect 525038 375107 525051 375141
rect 525085 375107 525098 375141
rect 525038 374741 525098 375107
rect 525038 374707 525051 374741
rect 525085 374707 525098 374741
rect 525038 374341 525098 374707
rect 525038 374307 525051 374341
rect 525085 374307 525098 374341
rect 525038 373941 525098 374307
rect 525038 373907 525051 373941
rect 525085 373907 525098 373941
rect 525038 373541 525098 373907
rect 525038 373507 525051 373541
rect 525085 373507 525098 373541
rect 525038 373141 525098 373507
rect 525038 373107 525051 373141
rect 525085 373107 525098 373141
rect 525038 372741 525098 373107
rect 525038 372707 525051 372741
rect 525085 372707 525098 372741
rect 525038 372341 525098 372707
rect 525038 372307 525051 372341
rect 525085 372307 525098 372341
rect 525038 371941 525098 372307
rect 525038 371907 525051 371941
rect 525085 371907 525098 371941
rect 525038 371541 525098 371907
rect 525038 371507 525051 371541
rect 525085 371507 525098 371541
rect 525038 371141 525098 371507
rect 525038 371107 525051 371141
rect 525085 371107 525098 371141
rect 525038 370741 525098 371107
rect 525038 370707 525051 370741
rect 525085 370707 525098 370741
rect 525038 370341 525098 370707
rect 525038 370307 525051 370341
rect 525085 370307 525098 370341
rect 525038 369941 525098 370307
rect 525038 369907 525051 369941
rect 525085 369907 525098 369941
rect 525038 369541 525098 369907
rect 525038 369507 525051 369541
rect 525085 369507 525098 369541
rect 525038 369141 525098 369507
rect 525038 369107 525051 369141
rect 525085 369107 525098 369141
rect 525038 368741 525098 369107
rect 525038 368707 525051 368741
rect 525085 368707 525098 368741
rect 525038 368341 525098 368707
rect 526918 370909 526978 371092
rect 526918 370875 526931 370909
rect 526965 370875 526978 370909
rect 526918 370709 526978 370875
rect 526918 370675 526931 370709
rect 526965 370675 526978 370709
rect 526918 370509 526978 370675
rect 528798 370909 528858 371092
rect 528798 370875 528811 370909
rect 528845 370875 528858 370909
rect 528798 370709 528858 370875
rect 528798 370675 528811 370709
rect 528845 370675 528858 370709
rect 526918 370475 526931 370509
rect 526965 370475 526978 370509
rect 526918 370309 526978 370475
rect 526918 370275 526931 370309
rect 526965 370275 526978 370309
rect 526918 370109 526978 370275
rect 528798 370509 528858 370675
rect 528798 370475 528811 370509
rect 528845 370475 528858 370509
rect 528798 370309 528858 370475
rect 528798 370275 528811 370309
rect 528845 370275 528858 370309
rect 528798 370180 528858 370275
rect 526918 370075 526931 370109
rect 526965 370075 526978 370109
rect 526918 369909 526978 370075
rect 526918 369875 526931 369909
rect 526965 369875 526978 369909
rect 526918 369709 526978 369875
rect 526918 369675 526931 369709
rect 526965 369675 526978 369709
rect 526918 369509 526978 369675
rect 527858 370109 528858 370180
rect 527858 370093 528811 370109
rect 527858 369651 527897 370093
rect 527999 370075 528811 370093
rect 528845 370075 528858 370109
rect 527999 369909 528858 370075
rect 527999 369875 528811 369909
rect 528845 369875 528858 369909
rect 527999 369709 528858 369875
rect 527999 369675 528811 369709
rect 528845 369675 528858 369709
rect 527999 369651 528858 369675
rect 527858 369564 528858 369651
rect 526918 369475 526931 369509
rect 526965 369475 526978 369509
rect 526918 369309 526978 369475
rect 526918 369275 526931 369309
rect 526965 369275 526978 369309
rect 526918 369109 526978 369275
rect 526918 369075 526931 369109
rect 526965 369075 526978 369109
rect 528798 369509 528858 369564
rect 528798 369475 528811 369509
rect 528845 369475 528858 369509
rect 528798 369309 528858 369475
rect 528798 369275 528811 369309
rect 528845 369275 528858 369309
rect 528798 369109 528858 369275
rect 526918 368909 526978 369075
rect 526918 368875 526931 368909
rect 526965 368875 526978 368909
rect 526918 368652 526978 368875
rect 527753 368652 528143 369084
rect 528798 369075 528811 369109
rect 528845 369075 528858 369109
rect 528798 368909 528858 369075
rect 528798 368875 528811 368909
rect 528845 368875 528858 368909
rect 528798 368652 528858 368875
rect 530678 371007 530738 371190
rect 530678 370973 530691 371007
rect 530725 370973 530738 371007
rect 530678 370807 530738 370973
rect 530678 370773 530691 370807
rect 530725 370773 530738 370807
rect 530678 370607 530738 370773
rect 532558 371007 532618 371190
rect 532558 370973 532571 371007
rect 532605 370973 532618 371007
rect 532558 370807 532618 370973
rect 532558 370773 532571 370807
rect 532605 370773 532618 370807
rect 530678 370573 530691 370607
rect 530725 370573 530738 370607
rect 530678 370407 530738 370573
rect 530678 370373 530691 370407
rect 530725 370373 530738 370407
rect 530678 370207 530738 370373
rect 532558 370607 532618 370773
rect 532558 370573 532571 370607
rect 532605 370573 532618 370607
rect 532558 370407 532618 370573
rect 532558 370373 532571 370407
rect 532605 370373 532618 370407
rect 532558 370278 532618 370373
rect 530678 370173 530691 370207
rect 530725 370173 530738 370207
rect 530678 370007 530738 370173
rect 530678 369973 530691 370007
rect 530725 369973 530738 370007
rect 530678 369807 530738 369973
rect 530678 369773 530691 369807
rect 530725 369773 530738 369807
rect 530678 369607 530738 369773
rect 531618 370207 532618 370278
rect 531618 370191 532571 370207
rect 531618 369749 531657 370191
rect 531759 370173 532571 370191
rect 532605 370173 532618 370207
rect 531759 370007 532618 370173
rect 531759 369973 532571 370007
rect 532605 369973 532618 370007
rect 531759 369807 532618 369973
rect 531759 369773 532571 369807
rect 532605 369773 532618 369807
rect 531759 369749 532618 369773
rect 531618 369662 532618 369749
rect 530678 369573 530691 369607
rect 530725 369573 530738 369607
rect 530678 369407 530738 369573
rect 530678 369373 530691 369407
rect 530725 369373 530738 369407
rect 530678 369207 530738 369373
rect 530678 369173 530691 369207
rect 530725 369173 530738 369207
rect 532558 369607 532618 369662
rect 532558 369573 532571 369607
rect 532605 369573 532618 369607
rect 532558 369407 532618 369573
rect 532558 369373 532571 369407
rect 532605 369373 532618 369407
rect 532558 369207 532618 369373
rect 530678 369007 530738 369173
rect 530678 368973 530691 369007
rect 530725 368973 530738 369007
rect 530678 368750 530738 368973
rect 531513 368750 531903 369182
rect 532558 369173 532571 369207
rect 532605 369173 532618 369207
rect 532558 369007 532618 369173
rect 532558 368973 532571 369007
rect 532605 368973 532618 369007
rect 532558 368750 532618 368973
rect 534438 370223 534498 370406
rect 534438 370189 534451 370223
rect 534485 370189 534498 370223
rect 534438 370023 534498 370189
rect 534438 369989 534451 370023
rect 534485 369989 534498 370023
rect 534438 369823 534498 369989
rect 536318 370223 536378 370406
rect 536318 370189 536331 370223
rect 536365 370189 536378 370223
rect 536318 370023 536378 370189
rect 536318 369989 536331 370023
rect 536365 369989 536378 370023
rect 534438 369789 534451 369823
rect 534485 369789 534498 369823
rect 534438 369623 534498 369789
rect 534438 369589 534451 369623
rect 534485 369589 534498 369623
rect 534438 369423 534498 369589
rect 536318 369823 536378 369989
rect 536318 369789 536331 369823
rect 536365 369789 536378 369823
rect 536318 369623 536378 369789
rect 536318 369589 536331 369623
rect 536365 369589 536378 369623
rect 536318 369494 536378 369589
rect 534438 369389 534451 369423
rect 534485 369389 534498 369423
rect 534438 369223 534498 369389
rect 534438 369189 534451 369223
rect 534485 369189 534498 369223
rect 534438 369023 534498 369189
rect 534438 368989 534451 369023
rect 534485 368989 534498 369023
rect 534438 368823 534498 368989
rect 535378 369423 536378 369494
rect 535378 369407 536331 369423
rect 535378 368965 535417 369407
rect 535519 369389 536331 369407
rect 536365 369389 536378 369423
rect 535519 369223 536378 369389
rect 535519 369189 536331 369223
rect 536365 369189 536378 369223
rect 535519 369023 536378 369189
rect 535519 368989 536331 369023
rect 536365 368989 536378 369023
rect 535519 368965 536378 368989
rect 535378 368878 536378 368965
rect 534438 368789 534451 368823
rect 534485 368789 534498 368823
rect 534438 368623 534498 368789
rect 534438 368589 534451 368623
rect 534485 368589 534498 368623
rect 525038 368307 525051 368341
rect 525085 368307 525098 368341
rect 525038 367941 525098 368307
rect 525038 367907 525051 367941
rect 525085 367907 525098 367941
rect 525038 367541 525098 367907
rect 525038 367507 525051 367541
rect 525085 367507 525098 367541
rect 525038 367141 525098 367507
rect 525038 367107 525051 367141
rect 525085 367107 525098 367141
rect 525038 366741 525098 367107
rect 525038 366707 525051 366741
rect 525085 366707 525098 366741
rect 525038 366341 525098 366707
rect 525038 366307 525051 366341
rect 525085 366307 525098 366341
rect 525038 365941 525098 366307
rect 525038 365907 525051 365941
rect 525085 365907 525098 365941
rect 526918 368165 526978 368348
rect 526918 368131 526931 368165
rect 526965 368131 526978 368165
rect 526918 367965 526978 368131
rect 526918 367931 526931 367965
rect 526965 367931 526978 367965
rect 526918 367765 526978 367931
rect 528798 368165 528858 368348
rect 528798 368131 528811 368165
rect 528845 368131 528858 368165
rect 528798 367965 528858 368131
rect 528798 367931 528811 367965
rect 528845 367931 528858 367965
rect 526918 367731 526931 367765
rect 526965 367731 526978 367765
rect 526918 367565 526978 367731
rect 526918 367531 526931 367565
rect 526965 367531 526978 367565
rect 526918 367365 526978 367531
rect 528798 367765 528858 367931
rect 528798 367731 528811 367765
rect 528845 367731 528858 367765
rect 528798 367565 528858 367731
rect 528798 367531 528811 367565
rect 528845 367531 528858 367565
rect 528798 367436 528858 367531
rect 526918 367331 526931 367365
rect 526965 367331 526978 367365
rect 526918 367165 526978 367331
rect 526918 367131 526931 367165
rect 526965 367131 526978 367165
rect 526918 366965 526978 367131
rect 526918 366931 526931 366965
rect 526965 366931 526978 366965
rect 526918 366765 526978 366931
rect 527858 367365 528858 367436
rect 527858 367349 528811 367365
rect 527858 366907 527897 367349
rect 527999 367331 528811 367349
rect 528845 367331 528858 367365
rect 527999 367165 528858 367331
rect 527999 367131 528811 367165
rect 528845 367131 528858 367165
rect 527999 366965 528858 367131
rect 527999 366931 528811 366965
rect 528845 366931 528858 366965
rect 527999 366907 528858 366931
rect 527858 366820 528858 366907
rect 526918 366731 526931 366765
rect 526965 366731 526978 366765
rect 526918 366565 526978 366731
rect 526918 366531 526931 366565
rect 526965 366531 526978 366565
rect 526918 366365 526978 366531
rect 526918 366331 526931 366365
rect 526965 366331 526978 366365
rect 528798 366765 528858 366820
rect 528798 366731 528811 366765
rect 528845 366731 528858 366765
rect 528798 366565 528858 366731
rect 528798 366531 528811 366565
rect 528845 366531 528858 366565
rect 528798 366365 528858 366531
rect 526918 366165 526978 366331
rect 526918 366131 526931 366165
rect 526965 366131 526978 366165
rect 526918 365908 526978 366131
rect 527753 365908 528143 366340
rect 528798 366331 528811 366365
rect 528845 366331 528858 366365
rect 528798 366165 528858 366331
rect 528798 366131 528811 366165
rect 528845 366131 528858 366165
rect 528798 365908 528858 366131
rect 530678 368263 530738 368446
rect 530678 368229 530691 368263
rect 530725 368229 530738 368263
rect 530678 368063 530738 368229
rect 530678 368029 530691 368063
rect 530725 368029 530738 368063
rect 530678 367863 530738 368029
rect 532558 368263 532618 368446
rect 532558 368229 532571 368263
rect 532605 368229 532618 368263
rect 532558 368063 532618 368229
rect 532558 368029 532571 368063
rect 532605 368029 532618 368063
rect 530678 367829 530691 367863
rect 530725 367829 530738 367863
rect 530678 367663 530738 367829
rect 530678 367629 530691 367663
rect 530725 367629 530738 367663
rect 530678 367463 530738 367629
rect 532558 367863 532618 368029
rect 534438 368423 534498 368589
rect 534438 368389 534451 368423
rect 534485 368389 534498 368423
rect 536318 368823 536378 368878
rect 536318 368789 536331 368823
rect 536365 368789 536378 368823
rect 536318 368623 536378 368789
rect 536318 368589 536331 368623
rect 536365 368589 536378 368623
rect 536318 368423 536378 368589
rect 534438 368223 534498 368389
rect 534438 368189 534451 368223
rect 534485 368189 534498 368223
rect 534438 367966 534498 368189
rect 535273 367966 535663 368398
rect 536318 368389 536331 368423
rect 536365 368389 536378 368423
rect 536318 368223 536378 368389
rect 536318 368189 536331 368223
rect 536365 368189 536378 368223
rect 536318 367966 536378 368189
rect 532558 367829 532571 367863
rect 532605 367829 532618 367863
rect 532558 367663 532618 367829
rect 532558 367629 532571 367663
rect 532605 367629 532618 367663
rect 532558 367534 532618 367629
rect 530678 367429 530691 367463
rect 530725 367429 530738 367463
rect 530678 367263 530738 367429
rect 530678 367229 530691 367263
rect 530725 367229 530738 367263
rect 530678 367063 530738 367229
rect 530678 367029 530691 367063
rect 530725 367029 530738 367063
rect 530678 366863 530738 367029
rect 531618 367463 532618 367534
rect 531618 367447 532571 367463
rect 531618 367005 531657 367447
rect 531759 367429 532571 367447
rect 532605 367429 532618 367463
rect 531759 367263 532618 367429
rect 531759 367229 532571 367263
rect 532605 367229 532618 367263
rect 531759 367063 532618 367229
rect 531759 367029 532571 367063
rect 532605 367029 532618 367063
rect 531759 367005 532618 367029
rect 531618 366918 532618 367005
rect 530678 366829 530691 366863
rect 530725 366829 530738 366863
rect 530678 366663 530738 366829
rect 530678 366629 530691 366663
rect 530725 366629 530738 366663
rect 530678 366463 530738 366629
rect 530678 366429 530691 366463
rect 530725 366429 530738 366463
rect 532558 366863 532618 366918
rect 532558 366829 532571 366863
rect 532605 366829 532618 366863
rect 532558 366663 532618 366829
rect 532558 366629 532571 366663
rect 532605 366629 532618 366663
rect 532558 366463 532618 366629
rect 530678 366263 530738 366429
rect 530678 366229 530691 366263
rect 530725 366229 530738 366263
rect 530678 366006 530738 366229
rect 531513 366006 531903 366438
rect 532558 366429 532571 366463
rect 532605 366429 532618 366463
rect 532558 366263 532618 366429
rect 532558 366229 532571 366263
rect 532605 366229 532618 366263
rect 532558 366006 532618 366229
rect 534438 367479 534498 367662
rect 534438 367445 534451 367479
rect 534485 367445 534498 367479
rect 534438 367279 534498 367445
rect 534438 367245 534451 367279
rect 534485 367245 534498 367279
rect 534438 367079 534498 367245
rect 536318 367479 536378 367662
rect 536318 367445 536331 367479
rect 536365 367445 536378 367479
rect 536318 367279 536378 367445
rect 536318 367245 536331 367279
rect 536365 367245 536378 367279
rect 534438 367045 534451 367079
rect 534485 367045 534498 367079
rect 534438 366879 534498 367045
rect 534438 366845 534451 366879
rect 534485 366845 534498 366879
rect 534438 366679 534498 366845
rect 536318 367079 536378 367245
rect 536318 367045 536331 367079
rect 536365 367045 536378 367079
rect 536318 366879 536378 367045
rect 536318 366845 536331 366879
rect 536365 366845 536378 366879
rect 536318 366750 536378 366845
rect 534438 366645 534451 366679
rect 534485 366645 534498 366679
rect 534438 366479 534498 366645
rect 534438 366445 534451 366479
rect 534485 366445 534498 366479
rect 534438 366279 534498 366445
rect 534438 366245 534451 366279
rect 534485 366245 534498 366279
rect 534438 366079 534498 366245
rect 535378 366679 536378 366750
rect 535378 366663 536331 366679
rect 535378 366221 535417 366663
rect 535519 366645 536331 366663
rect 536365 366645 536378 366679
rect 535519 366479 536378 366645
rect 535519 366445 536331 366479
rect 536365 366445 536378 366479
rect 535519 366279 536378 366445
rect 535519 366245 536331 366279
rect 536365 366245 536378 366279
rect 535519 366221 536378 366245
rect 535378 366134 536378 366221
rect 534438 366045 534451 366079
rect 534485 366045 534498 366079
rect 525038 365541 525098 365907
rect 534438 365879 534498 366045
rect 534438 365845 534451 365879
rect 534485 365845 534498 365879
rect 525038 365507 525051 365541
rect 525085 365507 525098 365541
rect 525038 365141 525098 365507
rect 525038 365107 525051 365141
rect 525085 365107 525098 365141
rect 525038 364741 525098 365107
rect 525038 364707 525051 364741
rect 525085 364707 525098 364741
rect 525038 364341 525098 364707
rect 525038 364307 525051 364341
rect 525085 364307 525098 364341
rect 525038 363941 525098 364307
rect 525038 363907 525051 363941
rect 525085 363907 525098 363941
rect 525038 363541 525098 363907
rect 525038 363507 525051 363541
rect 525085 363507 525098 363541
rect 525038 363141 525098 363507
rect 526918 365421 526978 365604
rect 526918 365387 526931 365421
rect 526965 365387 526978 365421
rect 526918 365221 526978 365387
rect 526918 365187 526931 365221
rect 526965 365187 526978 365221
rect 526918 365021 526978 365187
rect 528798 365421 528858 365604
rect 528798 365387 528811 365421
rect 528845 365387 528858 365421
rect 528798 365221 528858 365387
rect 528798 365187 528811 365221
rect 528845 365187 528858 365221
rect 526918 364987 526931 365021
rect 526965 364987 526978 365021
rect 526918 364821 526978 364987
rect 526918 364787 526931 364821
rect 526965 364787 526978 364821
rect 526918 364621 526978 364787
rect 528798 365021 528858 365187
rect 528798 364987 528811 365021
rect 528845 364987 528858 365021
rect 528798 364821 528858 364987
rect 528798 364787 528811 364821
rect 528845 364787 528858 364821
rect 528798 364692 528858 364787
rect 526918 364587 526931 364621
rect 526965 364587 526978 364621
rect 526918 364421 526978 364587
rect 526918 364387 526931 364421
rect 526965 364387 526978 364421
rect 526918 364221 526978 364387
rect 526918 364187 526931 364221
rect 526965 364187 526978 364221
rect 526918 364021 526978 364187
rect 527858 364621 528858 364692
rect 527858 364605 528811 364621
rect 527858 364163 527897 364605
rect 527999 364587 528811 364605
rect 528845 364587 528858 364621
rect 527999 364421 528858 364587
rect 527999 364387 528811 364421
rect 528845 364387 528858 364421
rect 527999 364221 528858 364387
rect 527999 364187 528811 364221
rect 528845 364187 528858 364221
rect 527999 364163 528858 364187
rect 527858 364076 528858 364163
rect 526918 363987 526931 364021
rect 526965 363987 526978 364021
rect 526918 363821 526978 363987
rect 526918 363787 526931 363821
rect 526965 363787 526978 363821
rect 526918 363621 526978 363787
rect 526918 363587 526931 363621
rect 526965 363587 526978 363621
rect 528798 364021 528858 364076
rect 528798 363987 528811 364021
rect 528845 363987 528858 364021
rect 528798 363821 528858 363987
rect 528798 363787 528811 363821
rect 528845 363787 528858 363821
rect 528798 363621 528858 363787
rect 526918 363421 526978 363587
rect 526918 363387 526931 363421
rect 526965 363387 526978 363421
rect 526918 363164 526978 363387
rect 527753 363164 528143 363596
rect 528798 363587 528811 363621
rect 528845 363587 528858 363621
rect 528798 363421 528858 363587
rect 528798 363387 528811 363421
rect 528845 363387 528858 363421
rect 528798 363164 528858 363387
rect 530678 365519 530738 365702
rect 530678 365485 530691 365519
rect 530725 365485 530738 365519
rect 530678 365319 530738 365485
rect 530678 365285 530691 365319
rect 530725 365285 530738 365319
rect 530678 365119 530738 365285
rect 532558 365519 532618 365702
rect 532558 365485 532571 365519
rect 532605 365485 532618 365519
rect 532558 365319 532618 365485
rect 532558 365285 532571 365319
rect 532605 365285 532618 365319
rect 530678 365085 530691 365119
rect 530725 365085 530738 365119
rect 530678 364919 530738 365085
rect 530678 364885 530691 364919
rect 530725 364885 530738 364919
rect 530678 364719 530738 364885
rect 532558 365119 532618 365285
rect 534438 365679 534498 365845
rect 534438 365645 534451 365679
rect 534485 365645 534498 365679
rect 536318 366079 536378 366134
rect 536318 366045 536331 366079
rect 536365 366045 536378 366079
rect 536318 365879 536378 366045
rect 536318 365845 536331 365879
rect 536365 365845 536378 365879
rect 536318 365679 536378 365845
rect 534438 365479 534498 365645
rect 534438 365445 534451 365479
rect 534485 365445 534498 365479
rect 534438 365222 534498 365445
rect 535273 365222 535663 365654
rect 536318 365645 536331 365679
rect 536365 365645 536378 365679
rect 536318 365479 536378 365645
rect 536318 365445 536331 365479
rect 536365 365445 536378 365479
rect 536318 365222 536378 365445
rect 532558 365085 532571 365119
rect 532605 365085 532618 365119
rect 532558 364919 532618 365085
rect 532558 364885 532571 364919
rect 532605 364885 532618 364919
rect 532558 364790 532618 364885
rect 530678 364685 530691 364719
rect 530725 364685 530738 364719
rect 530678 364519 530738 364685
rect 530678 364485 530691 364519
rect 530725 364485 530738 364519
rect 530678 364319 530738 364485
rect 530678 364285 530691 364319
rect 530725 364285 530738 364319
rect 530678 364119 530738 364285
rect 531618 364719 532618 364790
rect 531618 364703 532571 364719
rect 531618 364261 531657 364703
rect 531759 364685 532571 364703
rect 532605 364685 532618 364719
rect 531759 364519 532618 364685
rect 531759 364485 532571 364519
rect 532605 364485 532618 364519
rect 531759 364319 532618 364485
rect 531759 364285 532571 364319
rect 532605 364285 532618 364319
rect 531759 364261 532618 364285
rect 531618 364174 532618 364261
rect 530678 364085 530691 364119
rect 530725 364085 530738 364119
rect 530678 363919 530738 364085
rect 530678 363885 530691 363919
rect 530725 363885 530738 363919
rect 530678 363719 530738 363885
rect 530678 363685 530691 363719
rect 530725 363685 530738 363719
rect 532558 364119 532618 364174
rect 532558 364085 532571 364119
rect 532605 364085 532618 364119
rect 532558 363919 532618 364085
rect 532558 363885 532571 363919
rect 532605 363885 532618 363919
rect 532558 363719 532618 363885
rect 530678 363519 530738 363685
rect 530678 363485 530691 363519
rect 530725 363485 530738 363519
rect 530678 363262 530738 363485
rect 531513 363262 531903 363694
rect 532558 363685 532571 363719
rect 532605 363685 532618 363719
rect 532558 363519 532618 363685
rect 532558 363485 532571 363519
rect 532605 363485 532618 363519
rect 532558 363262 532618 363485
rect 534438 364735 534498 364918
rect 534438 364701 534451 364735
rect 534485 364701 534498 364735
rect 534438 364535 534498 364701
rect 534438 364501 534451 364535
rect 534485 364501 534498 364535
rect 534438 364335 534498 364501
rect 536318 364735 536378 364918
rect 536318 364701 536331 364735
rect 536365 364701 536378 364735
rect 536318 364535 536378 364701
rect 536318 364501 536331 364535
rect 536365 364501 536378 364535
rect 534438 364301 534451 364335
rect 534485 364301 534498 364335
rect 534438 364135 534498 364301
rect 534438 364101 534451 364135
rect 534485 364101 534498 364135
rect 534438 363935 534498 364101
rect 536318 364335 536378 364501
rect 536318 364301 536331 364335
rect 536365 364301 536378 364335
rect 536318 364135 536378 364301
rect 536318 364101 536331 364135
rect 536365 364101 536378 364135
rect 536318 364006 536378 364101
rect 534438 363901 534451 363935
rect 534485 363901 534498 363935
rect 534438 363735 534498 363901
rect 534438 363701 534451 363735
rect 534485 363701 534498 363735
rect 534438 363535 534498 363701
rect 534438 363501 534451 363535
rect 534485 363501 534498 363535
rect 534438 363335 534498 363501
rect 535378 363935 536378 364006
rect 535378 363919 536331 363935
rect 535378 363477 535417 363919
rect 535519 363901 536331 363919
rect 536365 363901 536378 363935
rect 535519 363735 536378 363901
rect 535519 363701 536331 363735
rect 536365 363701 536378 363735
rect 535519 363535 536378 363701
rect 535519 363501 536331 363535
rect 536365 363501 536378 363535
rect 535519 363477 536378 363501
rect 535378 363390 536378 363477
rect 534438 363301 534451 363335
rect 534485 363301 534498 363335
rect 525038 363107 525051 363141
rect 525085 363107 525098 363141
rect 525038 362741 525098 363107
rect 525038 362707 525051 362741
rect 525085 362707 525098 362741
rect 525038 362516 525098 362707
rect 534438 363135 534498 363301
rect 534438 363101 534451 363135
rect 534485 363101 534498 363135
rect 534438 362935 534498 363101
rect 534438 362901 534451 362935
rect 534485 362901 534498 362935
rect 536318 363335 536378 363390
rect 536318 363301 536331 363335
rect 536365 363301 536378 363335
rect 536318 363135 536378 363301
rect 536318 363101 536331 363135
rect 536365 363101 536378 363135
rect 536318 362935 536378 363101
rect 534438 362735 534498 362901
rect 534438 362701 534451 362735
rect 534485 362701 534498 362735
rect 534438 362478 534498 362701
rect 535273 362478 535663 362910
rect 536318 362901 536331 362935
rect 536365 362901 536378 362935
rect 536318 362735 536378 362901
rect 536318 362701 536331 362735
rect 536365 362701 536378 362735
rect 536318 362478 536378 362701
rect 560542 359330 560728 359390
rect 560788 359330 560928 359390
rect 560988 359330 561128 359390
rect 561188 359330 561328 359390
rect 561388 359330 561528 359390
rect 561588 359330 561728 359390
rect 561788 359330 561928 359390
rect 561988 359330 562128 359390
rect 562188 359330 562328 359390
rect 562388 359330 562528 359390
rect 562588 359330 562728 359390
rect 562788 359330 562928 359390
rect 562988 359330 563128 359390
rect 563188 359330 563328 359390
rect 563388 359330 563528 359390
rect 563588 359330 563728 359390
rect 563788 359330 563928 359390
rect 563988 359330 564128 359390
rect 564188 359330 564328 359390
rect 564388 359330 564528 359390
rect 564588 359330 564728 359390
rect 564788 359330 564928 359390
rect 564988 359330 565128 359390
rect 565188 359330 565328 359390
rect 565388 359330 565528 359390
rect 565588 359330 565856 359390
rect 574644 359260 574702 359320
rect 574762 359260 574902 359320
rect 574962 359260 575102 359320
rect 575162 359260 575302 359320
rect 575362 359260 575502 359320
rect 575562 359260 575702 359320
rect 575762 359260 575902 359320
rect 575962 359260 576102 359320
rect 576162 359260 576302 359320
rect 576362 359260 576502 359320
rect 576562 359260 576702 359320
rect 576762 359260 576902 359320
rect 576962 359260 577102 359320
rect 577162 359260 577302 359320
rect 577362 359260 577502 359320
rect 577562 359260 577702 359320
rect 577762 359260 577902 359320
rect 577962 359260 578102 359320
rect 578162 359260 578302 359320
rect 578362 359260 578502 359320
rect 578562 359260 578702 359320
rect 578762 359260 578902 359320
rect 578962 359260 579102 359320
rect 579162 359260 579302 359320
rect 579362 359260 579502 359320
rect 579562 359260 579702 359320
rect 579762 359260 580030 359320
rect 560280 359230 560340 359232
rect 560280 359170 565758 359230
rect 576194 359218 576354 359260
rect 576194 359182 576250 359218
rect 576294 359182 576354 359218
rect 576194 359180 576354 359182
rect 577494 359218 577654 359260
rect 577494 359182 577550 359218
rect 577594 359182 577654 359218
rect 577494 359180 577654 359182
rect 578794 359218 578954 359260
rect 578794 359182 578850 359218
rect 578894 359182 578954 359218
rect 578794 359180 578954 359182
rect 579942 359170 580002 359260
rect 560280 358062 560374 359170
rect 560234 358044 560374 358062
rect 560222 358022 560374 358044
rect 560222 357872 560232 358022
rect 560364 357872 560374 358022
rect 560553 358968 560587 358984
rect 560553 357976 560587 357992
rect 560811 358968 560845 359170
rect 560811 357976 560845 357992
rect 561069 358968 561103 358984
rect 561069 357910 561103 357992
rect 561327 358968 561361 359170
rect 561327 357976 561361 357992
rect 561585 358968 561619 358984
rect 561585 357910 561619 357992
rect 561843 358968 561877 359170
rect 561843 357976 561877 357992
rect 562101 358968 562135 358984
rect 562101 357910 562135 357992
rect 562359 358968 562393 359170
rect 562359 357976 562393 357992
rect 562617 358968 562651 358984
rect 562617 357910 562651 357992
rect 562875 358968 562909 359170
rect 562875 357976 562909 357992
rect 563133 358968 563167 358984
rect 563133 357910 563167 357992
rect 563391 358968 563425 359170
rect 563391 357976 563425 357992
rect 563649 358968 563683 358984
rect 563649 357910 563683 357992
rect 563907 358968 563941 359170
rect 563907 357976 563941 357992
rect 564165 358968 564199 358984
rect 564165 357910 564199 357992
rect 564423 358968 564457 359170
rect 564423 357976 564457 357992
rect 564681 358968 564715 358984
rect 564681 357910 564715 357992
rect 564939 358968 564973 359170
rect 564939 357976 564973 357992
rect 565197 358968 565231 358984
rect 565197 357910 565231 357992
rect 565455 358968 565489 359170
rect 574454 359140 574514 359142
rect 574454 359100 579872 359140
rect 579942 359130 579952 359170
rect 579992 359130 580002 359170
rect 574454 359080 579870 359100
rect 565455 357976 565489 357992
rect 565713 358968 565747 358984
rect 565713 357984 565747 357992
rect 565713 357964 565772 357984
rect 565713 357910 565966 357964
rect 560222 357852 560374 357872
rect 560280 357744 560374 357852
rect 560540 357860 565966 357910
rect 566126 357860 566132 357964
rect 560540 357850 566132 357860
rect 560280 357684 560728 357744
rect 560788 357684 560928 357744
rect 560988 357684 561128 357744
rect 561188 357684 561328 357744
rect 561388 357684 561528 357744
rect 561588 357684 561728 357744
rect 561788 357684 561928 357744
rect 561988 357684 562128 357744
rect 562188 357684 562328 357744
rect 562388 357684 562528 357744
rect 562588 357684 562728 357744
rect 562788 357684 562928 357744
rect 562988 357684 563128 357744
rect 563188 357684 563328 357744
rect 563388 357684 563528 357744
rect 563588 357684 563728 357744
rect 563788 357684 563928 357744
rect 563988 357684 564128 357744
rect 564188 357684 564328 357744
rect 564388 357684 564528 357744
rect 564588 357684 564728 357744
rect 564788 357684 564928 357744
rect 564988 357684 565128 357744
rect 565188 357684 565328 357744
rect 565388 357684 565528 357744
rect 565588 357684 565678 357744
rect 574454 357734 574514 359080
rect 574691 358898 574725 358914
rect 574691 357780 574725 357922
rect 574949 358898 574983 359080
rect 574949 357906 574983 357922
rect 575207 358898 575241 358914
rect 575207 357780 575241 357922
rect 575465 358898 575499 359080
rect 575465 357906 575499 357922
rect 575723 358898 575757 358914
rect 575723 357780 575757 357922
rect 575981 358898 576015 359080
rect 575981 357906 576015 357922
rect 576239 358898 576273 358914
rect 576239 357780 576273 357922
rect 576497 358898 576531 359080
rect 576497 357906 576531 357922
rect 576755 358898 576789 358914
rect 576755 357780 576789 357922
rect 577013 358898 577047 359080
rect 577013 357906 577047 357922
rect 577271 358898 577305 358914
rect 577271 357780 577305 357922
rect 577529 358898 577563 359080
rect 577529 357906 577563 357922
rect 577787 358898 577821 358914
rect 577787 357780 577821 357922
rect 578045 358898 578079 359080
rect 578045 357906 578079 357922
rect 578303 358898 578337 358914
rect 578303 357780 578337 357922
rect 578561 358898 578595 359080
rect 578561 357906 578595 357922
rect 578819 358898 578853 358914
rect 578819 357780 578853 357922
rect 579077 358898 579111 359080
rect 579077 357906 579111 357922
rect 579335 358898 579369 358914
rect 579335 357780 579369 357922
rect 579593 358898 579627 359080
rect 579942 359050 580002 359130
rect 579593 357906 579627 357922
rect 579851 358898 579885 358914
rect 579851 357824 579885 357922
rect 579851 357814 580116 357824
rect 579851 357780 580016 357814
rect 565768 357640 565828 357720
rect 562020 357608 562180 357630
rect 562020 357572 562076 357608
rect 562120 357572 562180 357608
rect 562020 357510 562180 357572
rect 563320 357608 563480 357630
rect 563320 357572 563376 357608
rect 563420 357572 563480 357608
rect 563320 357510 563480 357572
rect 564620 357608 564780 357630
rect 564620 357572 564676 357608
rect 564720 357572 564780 357608
rect 564620 357510 564780 357572
rect 565768 357600 565778 357640
rect 565818 357600 565828 357640
rect 565768 357510 565828 357600
rect 574398 357680 574514 357734
rect 574638 357726 580016 357780
rect 580106 357726 580116 357814
rect 574638 357720 580116 357726
rect 574398 357576 574408 357680
rect 574500 357618 574514 357680
rect 574500 357576 574702 357618
rect 574398 357560 574702 357576
rect 574436 357558 574702 357560
rect 574762 357558 574902 357618
rect 574962 357558 575102 357618
rect 575162 357558 575302 357618
rect 575362 357558 575502 357618
rect 575562 357558 575702 357618
rect 575762 357558 575902 357618
rect 575962 357558 576102 357618
rect 576162 357558 576302 357618
rect 576362 357558 576502 357618
rect 576562 357558 576702 357618
rect 576762 357558 576902 357618
rect 576962 357558 577102 357618
rect 577162 357558 577302 357618
rect 577362 357558 577502 357618
rect 577562 357558 577702 357618
rect 577762 357558 577902 357618
rect 577962 357558 578102 357618
rect 578162 357558 578302 357618
rect 578362 357558 578502 357618
rect 578562 357558 578702 357618
rect 578762 357558 578902 357618
rect 578962 357558 579102 357618
rect 579162 357558 579302 357618
rect 579362 357558 579502 357618
rect 579562 357558 579702 357618
rect 579762 357558 579932 357618
rect 560542 357450 560728 357510
rect 560788 357450 560928 357510
rect 560988 357450 561128 357510
rect 561188 357450 561328 357510
rect 561388 357450 561528 357510
rect 561588 357450 561728 357510
rect 561788 357450 561928 357510
rect 561988 357450 562128 357510
rect 562188 357450 562328 357510
rect 562388 357450 562528 357510
rect 562588 357450 562728 357510
rect 562788 357450 562928 357510
rect 562988 357450 563128 357510
rect 563188 357450 563328 357510
rect 563388 357450 563528 357510
rect 563588 357450 563728 357510
rect 563788 357450 563928 357510
rect 563988 357450 564128 357510
rect 564188 357450 564328 357510
rect 564388 357450 564528 357510
rect 564588 357450 564728 357510
rect 564788 357450 564928 357510
rect 564988 357450 565128 357510
rect 565188 357450 565328 357510
rect 565388 357450 565528 357510
rect 565588 357450 565856 357510
rect 574644 357380 574702 357440
rect 574762 357380 574902 357440
rect 574962 357380 575102 357440
rect 575162 357380 575302 357440
rect 575362 357380 575502 357440
rect 575562 357380 575702 357440
rect 575762 357380 575902 357440
rect 575962 357380 576102 357440
rect 576162 357380 576302 357440
rect 576362 357380 576502 357440
rect 576562 357380 576702 357440
rect 576762 357380 576902 357440
rect 576962 357380 577102 357440
rect 577162 357380 577302 357440
rect 577362 357380 577502 357440
rect 577562 357380 577702 357440
rect 577762 357380 577902 357440
rect 577962 357380 578102 357440
rect 578162 357380 578302 357440
rect 578362 357380 578502 357440
rect 578562 357380 578702 357440
rect 578762 357380 578902 357440
rect 578962 357380 579102 357440
rect 579162 357380 579302 357440
rect 579362 357380 579502 357440
rect 579562 357380 579702 357440
rect 579762 357380 580030 357440
rect 575092 313092 575150 313152
rect 575210 313092 575350 313152
rect 575410 313092 575550 313152
rect 575610 313092 575750 313152
rect 575810 313092 575950 313152
rect 576010 313092 576150 313152
rect 576210 313092 576350 313152
rect 576410 313092 576550 313152
rect 576610 313092 576750 313152
rect 576810 313092 576950 313152
rect 577010 313092 577150 313152
rect 577210 313092 577350 313152
rect 577410 313092 577550 313152
rect 577610 313092 577750 313152
rect 577810 313092 577950 313152
rect 578010 313092 578150 313152
rect 578210 313092 578350 313152
rect 578410 313092 578550 313152
rect 578610 313092 578750 313152
rect 578810 313092 578950 313152
rect 579010 313092 579150 313152
rect 579210 313092 579350 313152
rect 579410 313092 579550 313152
rect 579610 313092 579750 313152
rect 579810 313092 579950 313152
rect 580010 313092 580150 313152
rect 580210 313092 580478 313152
rect 560404 313022 560590 313082
rect 560650 313022 560790 313082
rect 560850 313022 560990 313082
rect 561050 313022 561190 313082
rect 561250 313022 561390 313082
rect 561450 313022 561590 313082
rect 561650 313022 561790 313082
rect 561850 313022 561990 313082
rect 562050 313022 562190 313082
rect 562250 313022 562390 313082
rect 562450 313022 562590 313082
rect 562650 313022 562790 313082
rect 562850 313022 562990 313082
rect 563050 313022 563190 313082
rect 563250 313022 563390 313082
rect 563450 313022 563590 313082
rect 563650 313022 563790 313082
rect 563850 313022 563990 313082
rect 564050 313022 564190 313082
rect 564250 313022 564390 313082
rect 564450 313022 564590 313082
rect 564650 313022 564790 313082
rect 564850 313022 564990 313082
rect 565050 313022 565190 313082
rect 565250 313022 565390 313082
rect 565450 313022 565718 313082
rect 576642 313050 576802 313092
rect 576642 313014 576698 313050
rect 576742 313014 576802 313050
rect 576642 313012 576802 313014
rect 577942 313050 578102 313092
rect 577942 313014 577998 313050
rect 578042 313014 578102 313050
rect 577942 313012 578102 313014
rect 579242 313050 579402 313092
rect 579242 313014 579298 313050
rect 579342 313014 579402 313050
rect 579242 313012 579402 313014
rect 580390 313002 580450 313092
rect 574902 312972 574962 312974
rect 574902 312932 580320 312972
rect 580390 312962 580400 313002
rect 580440 312962 580450 313002
rect 560142 312922 560202 312924
rect 560142 312862 565620 312922
rect 574902 312912 580318 312932
rect 560142 311754 560236 312862
rect 560096 311736 560236 311754
rect 560084 311714 560236 311736
rect 560084 311564 560094 311714
rect 560226 311564 560236 311714
rect 560415 312660 560449 312676
rect 560415 311668 560449 311684
rect 560673 312660 560707 312862
rect 560673 311668 560707 311684
rect 560931 312660 560965 312676
rect 560931 311602 560965 311684
rect 561189 312660 561223 312862
rect 561189 311668 561223 311684
rect 561447 312660 561481 312676
rect 561447 311602 561481 311684
rect 561705 312660 561739 312862
rect 561705 311668 561739 311684
rect 561963 312660 561997 312676
rect 561963 311602 561997 311684
rect 562221 312660 562255 312862
rect 562221 311668 562255 311684
rect 562479 312660 562513 312676
rect 562479 311602 562513 311684
rect 562737 312660 562771 312862
rect 562737 311668 562771 311684
rect 562995 312660 563029 312676
rect 562995 311602 563029 311684
rect 563253 312660 563287 312862
rect 563253 311668 563287 311684
rect 563511 312660 563545 312676
rect 563511 311602 563545 311684
rect 563769 312660 563803 312862
rect 563769 311668 563803 311684
rect 564027 312660 564061 312676
rect 564027 311602 564061 311684
rect 564285 312660 564319 312862
rect 564285 311668 564319 311684
rect 564543 312660 564577 312676
rect 564543 311602 564577 311684
rect 564801 312660 564835 312862
rect 564801 311668 564835 311684
rect 565059 312660 565093 312676
rect 565059 311602 565093 311684
rect 565317 312660 565351 312862
rect 565317 311668 565351 311684
rect 565575 312660 565609 312676
rect 565575 311676 565609 311684
rect 565575 311656 565634 311676
rect 565575 311602 565828 311656
rect 560084 311544 560236 311564
rect 560142 311436 560236 311544
rect 560402 311552 565828 311602
rect 565988 311552 565994 311656
rect 574902 311566 574962 312912
rect 575139 312730 575173 312746
rect 575139 311612 575173 311754
rect 575397 312730 575431 312912
rect 575397 311738 575431 311754
rect 575655 312730 575689 312746
rect 575655 311612 575689 311754
rect 575913 312730 575947 312912
rect 575913 311738 575947 311754
rect 576171 312730 576205 312746
rect 576171 311612 576205 311754
rect 576429 312730 576463 312912
rect 576429 311738 576463 311754
rect 576687 312730 576721 312746
rect 576687 311612 576721 311754
rect 576945 312730 576979 312912
rect 576945 311738 576979 311754
rect 577203 312730 577237 312746
rect 577203 311612 577237 311754
rect 577461 312730 577495 312912
rect 577461 311738 577495 311754
rect 577719 312730 577753 312746
rect 577719 311612 577753 311754
rect 577977 312730 578011 312912
rect 577977 311738 578011 311754
rect 578235 312730 578269 312746
rect 578235 311612 578269 311754
rect 578493 312730 578527 312912
rect 578493 311738 578527 311754
rect 578751 312730 578785 312746
rect 578751 311612 578785 311754
rect 579009 312730 579043 312912
rect 579009 311738 579043 311754
rect 579267 312730 579301 312746
rect 579267 311612 579301 311754
rect 579525 312730 579559 312912
rect 579525 311738 579559 311754
rect 579783 312730 579817 312746
rect 579783 311612 579817 311754
rect 580041 312730 580075 312912
rect 580390 312882 580450 312962
rect 580041 311738 580075 311754
rect 580299 312730 580333 312746
rect 580299 311656 580333 311754
rect 580299 311646 580564 311656
rect 580299 311612 580464 311646
rect 560402 311542 565994 311552
rect 574846 311512 574962 311566
rect 575086 311558 580464 311612
rect 580554 311558 580564 311646
rect 575086 311552 580564 311558
rect 560142 311376 560590 311436
rect 560650 311376 560790 311436
rect 560850 311376 560990 311436
rect 561050 311376 561190 311436
rect 561250 311376 561390 311436
rect 561450 311376 561590 311436
rect 561650 311376 561790 311436
rect 561850 311376 561990 311436
rect 562050 311376 562190 311436
rect 562250 311376 562390 311436
rect 562450 311376 562590 311436
rect 562650 311376 562790 311436
rect 562850 311376 562990 311436
rect 563050 311376 563190 311436
rect 563250 311376 563390 311436
rect 563450 311376 563590 311436
rect 563650 311376 563790 311436
rect 563850 311376 563990 311436
rect 564050 311376 564190 311436
rect 564250 311376 564390 311436
rect 564450 311376 564590 311436
rect 564650 311376 564790 311436
rect 564850 311376 564990 311436
rect 565050 311376 565190 311436
rect 565250 311376 565390 311436
rect 565450 311376 565540 311436
rect 565630 311332 565690 311412
rect 574846 311408 574856 311512
rect 574948 311450 574962 311512
rect 574948 311408 575150 311450
rect 574846 311392 575150 311408
rect 574884 311390 575150 311392
rect 575210 311390 575350 311450
rect 575410 311390 575550 311450
rect 575610 311390 575750 311450
rect 575810 311390 575950 311450
rect 576010 311390 576150 311450
rect 576210 311390 576350 311450
rect 576410 311390 576550 311450
rect 576610 311390 576750 311450
rect 576810 311390 576950 311450
rect 577010 311390 577150 311450
rect 577210 311390 577350 311450
rect 577410 311390 577550 311450
rect 577610 311390 577750 311450
rect 577810 311390 577950 311450
rect 578010 311390 578150 311450
rect 578210 311390 578350 311450
rect 578410 311390 578550 311450
rect 578610 311390 578750 311450
rect 578810 311390 578950 311450
rect 579010 311390 579150 311450
rect 579210 311390 579350 311450
rect 579410 311390 579550 311450
rect 579610 311390 579750 311450
rect 579810 311390 579950 311450
rect 580010 311390 580150 311450
rect 580210 311390 580380 311450
rect 561882 311300 562042 311322
rect 561882 311264 561938 311300
rect 561982 311264 562042 311300
rect 561882 311202 562042 311264
rect 563182 311300 563342 311322
rect 563182 311264 563238 311300
rect 563282 311264 563342 311300
rect 563182 311202 563342 311264
rect 564482 311300 564642 311322
rect 564482 311264 564538 311300
rect 564582 311264 564642 311300
rect 564482 311202 564642 311264
rect 565630 311292 565640 311332
rect 565680 311292 565690 311332
rect 565630 311202 565690 311292
rect 575092 311212 575150 311272
rect 575210 311212 575350 311272
rect 575410 311212 575550 311272
rect 575610 311212 575750 311272
rect 575810 311212 575950 311272
rect 576010 311212 576150 311272
rect 576210 311212 576350 311272
rect 576410 311212 576550 311272
rect 576610 311212 576750 311272
rect 576810 311212 576950 311272
rect 577010 311212 577150 311272
rect 577210 311212 577350 311272
rect 577410 311212 577550 311272
rect 577610 311212 577750 311272
rect 577810 311212 577950 311272
rect 578010 311212 578150 311272
rect 578210 311212 578350 311272
rect 578410 311212 578550 311272
rect 578610 311212 578750 311272
rect 578810 311212 578950 311272
rect 579010 311212 579150 311272
rect 579210 311212 579350 311272
rect 579410 311212 579550 311272
rect 579610 311212 579750 311272
rect 579810 311212 579950 311272
rect 580010 311212 580150 311272
rect 580210 311212 580478 311272
rect 560404 311142 560590 311202
rect 560650 311142 560790 311202
rect 560850 311142 560990 311202
rect 561050 311142 561190 311202
rect 561250 311142 561390 311202
rect 561450 311142 561590 311202
rect 561650 311142 561790 311202
rect 561850 311142 561990 311202
rect 562050 311142 562190 311202
rect 562250 311142 562390 311202
rect 562450 311142 562590 311202
rect 562650 311142 562790 311202
rect 562850 311142 562990 311202
rect 563050 311142 563190 311202
rect 563250 311142 563390 311202
rect 563450 311142 563590 311202
rect 563650 311142 563790 311202
rect 563850 311142 563990 311202
rect 564050 311142 564190 311202
rect 564250 311142 564390 311202
rect 564450 311142 564590 311202
rect 564650 311142 564790 311202
rect 564850 311142 564990 311202
rect 565050 311142 565190 311202
rect 565250 311142 565390 311202
rect 565450 311142 565718 311202
<< viali >>
rect 560836 493790 560896 493850
rect 561036 493790 561096 493850
rect 561236 493790 561296 493850
rect 561436 493790 561496 493850
rect 561636 493790 561696 493850
rect 561836 493790 561896 493850
rect 562036 493790 562096 493850
rect 562236 493790 562296 493850
rect 562436 493790 562496 493850
rect 562636 493790 562696 493850
rect 562836 493790 562896 493850
rect 563036 493790 563096 493850
rect 563236 493790 563296 493850
rect 563436 493790 563496 493850
rect 563636 493790 563696 493850
rect 563836 493790 563896 493850
rect 564036 493790 564096 493850
rect 564236 493790 564296 493850
rect 564436 493790 564496 493850
rect 564636 493790 564696 493850
rect 564836 493790 564896 493850
rect 565036 493790 565096 493850
rect 565236 493790 565296 493850
rect 565436 493790 565496 493850
rect 565636 493790 565696 493850
rect 560340 492332 560472 492482
rect 560661 492452 560695 493428
rect 560919 492452 560953 493428
rect 561177 492452 561211 493428
rect 561435 492452 561469 493428
rect 561693 492452 561727 493428
rect 561951 492452 561985 493428
rect 562209 492452 562243 493428
rect 562467 492452 562501 493428
rect 562725 492452 562759 493428
rect 562983 492452 563017 493428
rect 563241 492452 563275 493428
rect 563499 492452 563533 493428
rect 563757 492452 563791 493428
rect 564015 492452 564049 493428
rect 564273 492452 564307 493428
rect 564531 492452 564565 493428
rect 564789 492452 564823 493428
rect 565047 492452 565081 493428
rect 565305 492452 565339 493428
rect 575228 493564 575288 493624
rect 575428 493564 575488 493624
rect 575628 493564 575688 493624
rect 575828 493564 575888 493624
rect 576028 493564 576088 493624
rect 576228 493564 576288 493624
rect 576428 493564 576488 493624
rect 576628 493564 576688 493624
rect 576828 493564 576888 493624
rect 577028 493564 577088 493624
rect 577228 493564 577288 493624
rect 577428 493564 577488 493624
rect 577628 493564 577688 493624
rect 577828 493564 577888 493624
rect 578028 493564 578088 493624
rect 578228 493564 578288 493624
rect 578428 493564 578488 493624
rect 578628 493564 578688 493624
rect 578828 493564 578888 493624
rect 579028 493564 579088 493624
rect 579228 493564 579288 493624
rect 579428 493564 579488 493624
rect 579628 493564 579688 493624
rect 579828 493564 579888 493624
rect 580028 493564 580088 493624
rect 580228 493564 580288 493624
rect 565563 492452 565597 493428
rect 565821 492452 565855 493428
rect 566074 492320 566234 492428
rect 575217 492226 575251 493202
rect 575475 492226 575509 493202
rect 575733 492226 575767 493202
rect 575991 492226 576025 493202
rect 576249 492226 576283 493202
rect 576507 492226 576541 493202
rect 576765 492226 576799 493202
rect 577023 492226 577057 493202
rect 577281 492226 577315 493202
rect 577539 492226 577573 493202
rect 577797 492226 577831 493202
rect 578055 492226 578089 493202
rect 578313 492226 578347 493202
rect 578571 492226 578605 493202
rect 578829 492226 578863 493202
rect 579087 492226 579121 493202
rect 579345 492226 579379 493202
rect 579603 492226 579637 493202
rect 579861 492226 579895 493202
rect 580119 492226 580153 493202
rect 580377 492226 580411 493202
rect 580542 492030 580632 492118
rect 560836 491910 560896 491970
rect 561036 491910 561096 491970
rect 561236 491910 561296 491970
rect 561436 491910 561496 491970
rect 561636 491910 561696 491970
rect 561836 491910 561896 491970
rect 562036 491910 562096 491970
rect 562236 491910 562296 491970
rect 562436 491910 562496 491970
rect 562636 491910 562696 491970
rect 562836 491910 562896 491970
rect 563036 491910 563096 491970
rect 563236 491910 563296 491970
rect 563436 491910 563496 491970
rect 563636 491910 563696 491970
rect 563836 491910 563896 491970
rect 564036 491910 564096 491970
rect 564236 491910 564296 491970
rect 564436 491910 564496 491970
rect 564636 491910 564696 491970
rect 564836 491910 564896 491970
rect 565036 491910 565096 491970
rect 565236 491910 565296 491970
rect 565436 491910 565496 491970
rect 565636 491910 565696 491970
rect 574934 491880 575026 491984
rect 575228 491684 575288 491744
rect 575428 491684 575488 491744
rect 575628 491684 575688 491744
rect 575828 491684 575888 491744
rect 576028 491684 576088 491744
rect 576228 491684 576288 491744
rect 576428 491684 576488 491744
rect 576628 491684 576688 491744
rect 576828 491684 576888 491744
rect 577028 491684 577088 491744
rect 577228 491684 577288 491744
rect 577428 491684 577488 491744
rect 577628 491684 577688 491744
rect 577828 491684 577888 491744
rect 578028 491684 578088 491744
rect 578228 491684 578288 491744
rect 578428 491684 578488 491744
rect 578628 491684 578688 491744
rect 578828 491684 578888 491744
rect 579028 491684 579088 491744
rect 579228 491684 579288 491744
rect 579428 491684 579488 491744
rect 579628 491684 579688 491744
rect 579828 491684 579888 491744
rect 580028 491684 580088 491744
rect 580228 491684 580288 491744
rect 493091 408819 493125 408853
rect 493091 408419 493125 408453
rect 493091 408019 493125 408053
rect 493091 407619 493125 407653
rect 493091 407219 493125 407253
rect 493091 406819 493125 406853
rect 493091 406419 493125 406453
rect 493091 406019 493125 406053
rect 493091 405619 493125 405653
rect 493091 405219 493125 405253
rect 493091 404819 493125 404853
rect 493091 404419 493125 404453
rect 493091 404019 493125 404053
rect 493091 403619 493125 403653
rect 493091 403219 493125 403253
rect 493091 402819 493125 402853
rect 493091 402419 493125 402453
rect 493091 402019 493125 402053
rect 494971 408819 495005 408853
rect 494971 408419 495005 408453
rect 494971 408019 495005 408053
rect 494971 407619 495005 407653
rect 494971 407219 495005 407253
rect 494971 406819 495005 406853
rect 494971 406419 495005 406453
rect 494971 406019 495005 406053
rect 494971 405619 495005 405653
rect 494971 405219 495005 405253
rect 494971 404819 495005 404853
rect 494971 404419 495005 404453
rect 494971 404019 495005 404053
rect 494971 403619 495005 403653
rect 494971 403219 495005 403253
rect 494971 402819 495005 402853
rect 494971 402419 495005 402453
rect 494971 402019 495005 402053
rect 496851 408819 496885 408853
rect 496851 408419 496885 408453
rect 496851 408019 496885 408053
rect 496851 407619 496885 407653
rect 496851 407219 496885 407253
rect 496851 406819 496885 406853
rect 496851 406419 496885 406453
rect 496851 406019 496885 406053
rect 496851 405619 496885 405653
rect 496851 405219 496885 405253
rect 496851 404819 496885 404853
rect 496851 404419 496885 404453
rect 496851 404019 496885 404053
rect 496851 403619 496885 403653
rect 496851 403219 496885 403253
rect 496851 402819 496885 402853
rect 496851 402419 496885 402453
rect 496851 402019 496885 402053
rect 498731 408819 498765 408853
rect 498731 408419 498765 408453
rect 498731 408019 498765 408053
rect 498731 407619 498765 407653
rect 498731 407219 498765 407253
rect 498731 406819 498765 406853
rect 498731 406419 498765 406453
rect 498731 406019 498765 406053
rect 498731 405619 498765 405653
rect 498731 405219 498765 405253
rect 498731 404819 498765 404853
rect 498731 404419 498765 404453
rect 498731 404019 498765 404053
rect 498731 403619 498765 403653
rect 498731 403219 498765 403253
rect 498731 402819 498765 402853
rect 498731 402419 498765 402453
rect 498731 402019 498765 402053
rect 500611 408427 500645 408461
rect 500611 408027 500645 408061
rect 500611 407627 500645 407661
rect 500611 407227 500645 407261
rect 500611 406827 500645 406861
rect 500611 406427 500645 406461
rect 500611 406027 500645 406061
rect 500611 405627 500645 405661
rect 500611 405227 500645 405261
rect 500611 404827 500645 404861
rect 500611 404427 500645 404461
rect 500611 404027 500645 404061
rect 500611 403627 500645 403661
rect 500611 403227 500645 403261
rect 500611 402827 500645 402861
rect 500611 402427 500645 402461
rect 500611 402027 500645 402061
rect 500611 401627 500645 401661
rect 493091 401371 493125 401405
rect 493091 400971 493125 401005
rect 493091 400571 493125 400605
rect 493091 400171 493125 400205
rect 493091 399771 493125 399805
rect 493091 399371 493125 399405
rect 493091 398971 493125 399005
rect 493091 398571 493125 398605
rect 493091 398171 493125 398205
rect 493091 397771 493125 397805
rect 493091 397371 493125 397405
rect 493091 396971 493125 397005
rect 493091 396571 493125 396605
rect 493091 396171 493125 396205
rect 493091 395771 493125 395805
rect 493091 395371 493125 395405
rect 493091 394971 493125 395005
rect 493091 394571 493125 394605
rect 502491 408427 502525 408461
rect 502491 408027 502525 408061
rect 502491 407627 502525 407661
rect 502491 407227 502525 407261
rect 502491 406827 502525 406861
rect 502491 406427 502525 406461
rect 502491 406027 502525 406061
rect 502491 405627 502525 405661
rect 502491 405227 502525 405261
rect 502491 404827 502525 404861
rect 560860 404648 560920 404708
rect 561060 404648 561120 404708
rect 561260 404648 561320 404708
rect 561460 404648 561520 404708
rect 561660 404648 561720 404708
rect 561860 404648 561920 404708
rect 562060 404648 562120 404708
rect 562260 404648 562320 404708
rect 562460 404648 562520 404708
rect 562660 404648 562720 404708
rect 562860 404648 562920 404708
rect 563060 404648 563120 404708
rect 563260 404648 563320 404708
rect 563460 404648 563520 404708
rect 563660 404648 563720 404708
rect 563860 404648 563920 404708
rect 564060 404648 564120 404708
rect 564260 404648 564320 404708
rect 564460 404648 564520 404708
rect 564660 404648 564720 404708
rect 564860 404648 564920 404708
rect 565060 404648 565120 404708
rect 565260 404648 565320 404708
rect 565460 404648 565520 404708
rect 565660 404648 565720 404708
rect 574506 404688 574566 404748
rect 574706 404688 574766 404748
rect 574906 404688 574966 404748
rect 575106 404688 575166 404748
rect 575306 404688 575366 404748
rect 575506 404688 575566 404748
rect 575706 404688 575766 404748
rect 575906 404688 575966 404748
rect 576106 404688 576166 404748
rect 576306 404688 576366 404748
rect 576506 404688 576566 404748
rect 576706 404688 576766 404748
rect 576906 404688 576966 404748
rect 577106 404688 577166 404748
rect 577306 404688 577366 404748
rect 577506 404688 577566 404748
rect 577706 404688 577766 404748
rect 577906 404688 577966 404748
rect 578106 404688 578166 404748
rect 578306 404688 578366 404748
rect 578506 404688 578566 404748
rect 578706 404688 578766 404748
rect 578906 404688 578966 404748
rect 579106 404688 579166 404748
rect 579306 404688 579366 404748
rect 579506 404688 579566 404748
rect 502491 404427 502525 404461
rect 502491 404027 502525 404061
rect 502491 403627 502525 403661
rect 560701 403310 560735 404286
rect 502491 403227 502525 403261
rect 560322 403178 560482 403286
rect 560959 403310 560993 404286
rect 561217 403310 561251 404286
rect 561475 403310 561509 404286
rect 561733 403310 561767 404286
rect 561991 403310 562025 404286
rect 562249 403310 562283 404286
rect 562507 403310 562541 404286
rect 562765 403310 562799 404286
rect 563023 403310 563057 404286
rect 563281 403310 563315 404286
rect 563539 403310 563573 404286
rect 563797 403310 563831 404286
rect 564055 403310 564089 404286
rect 564313 403310 564347 404286
rect 564571 403310 564605 404286
rect 564829 403310 564863 404286
rect 565087 403310 565121 404286
rect 565345 403310 565379 404286
rect 565603 403310 565637 404286
rect 565861 403310 565895 404286
rect 566084 403190 566216 403340
rect 574495 403350 574529 404326
rect 574753 403350 574787 404326
rect 575011 403350 575045 404326
rect 575269 403350 575303 404326
rect 575527 403350 575561 404326
rect 575785 403350 575819 404326
rect 576043 403350 576077 404326
rect 576301 403350 576335 404326
rect 576559 403350 576593 404326
rect 576817 403350 576851 404326
rect 577075 403350 577109 404326
rect 577333 403350 577367 404326
rect 577591 403350 577625 404326
rect 577849 403350 577883 404326
rect 578107 403350 578141 404326
rect 578365 403350 578399 404326
rect 578623 403350 578657 404326
rect 578881 403350 578915 404326
rect 579139 403350 579173 404326
rect 579397 403350 579431 404326
rect 579655 403350 579689 404326
rect 502491 402827 502525 402861
rect 502491 402427 502525 402461
rect 502491 402027 502525 402061
rect 502491 401627 502525 401661
rect 504371 402745 504405 402779
rect 504371 402545 504405 402579
rect 504371 402345 504405 402379
rect 504371 402145 504405 402179
rect 504371 401945 504405 401979
rect 504371 401745 504405 401779
rect 505068 402544 505074 402566
rect 505074 402544 505102 402566
rect 505068 402532 505102 402544
rect 505168 402532 505202 402566
rect 505268 402532 505302 402566
rect 505368 402544 505400 402566
rect 505400 402544 505402 402566
rect 505468 402544 505490 402566
rect 505490 402544 505502 402566
rect 505568 402544 505580 402566
rect 505580 402544 505602 402566
rect 505368 402532 505402 402544
rect 505468 402532 505502 402544
rect 505568 402532 505602 402544
rect 505068 402454 505074 402466
rect 505074 402454 505102 402466
rect 505068 402432 505102 402454
rect 505168 402432 505202 402466
rect 505268 402432 505302 402466
rect 505368 402454 505400 402466
rect 505400 402454 505402 402466
rect 505468 402454 505490 402466
rect 505490 402454 505502 402466
rect 505568 402454 505580 402466
rect 505580 402454 505602 402466
rect 505368 402432 505402 402454
rect 505468 402432 505502 402454
rect 505568 402432 505602 402454
rect 505068 402364 505074 402366
rect 505074 402364 505102 402366
rect 505068 402332 505102 402364
rect 505168 402332 505202 402366
rect 505268 402332 505302 402366
rect 505368 402364 505400 402366
rect 505400 402364 505402 402366
rect 505468 402364 505490 402366
rect 505490 402364 505502 402366
rect 505568 402364 505580 402366
rect 505580 402364 505602 402366
rect 505368 402332 505402 402364
rect 505468 402332 505502 402364
rect 505568 402332 505602 402364
rect 505068 402232 505102 402266
rect 505168 402232 505202 402266
rect 505268 402232 505302 402266
rect 505368 402232 505402 402266
rect 505468 402232 505502 402266
rect 505568 402232 505602 402266
rect 505068 402132 505102 402166
rect 505168 402132 505202 402166
rect 505268 402132 505302 402166
rect 505368 402132 505402 402166
rect 505468 402132 505502 402166
rect 505568 402132 505602 402166
rect 505068 402038 505102 402066
rect 505068 402032 505074 402038
rect 505074 402032 505102 402038
rect 505168 402032 505202 402066
rect 505268 402032 505302 402066
rect 505368 402038 505402 402066
rect 505468 402038 505502 402066
rect 505568 402038 505602 402066
rect 505368 402032 505400 402038
rect 505400 402032 505402 402038
rect 505468 402032 505490 402038
rect 505490 402032 505502 402038
rect 505568 402032 505580 402038
rect 505580 402032 505602 402038
rect 505765 401827 505799 401861
rect 505901 401643 505935 401677
rect 579820 403154 579910 403242
rect 574212 403004 574304 403108
rect 506251 402745 506285 402779
rect 560860 402768 560920 402828
rect 561060 402768 561120 402828
rect 561260 402768 561320 402828
rect 561460 402768 561520 402828
rect 561660 402768 561720 402828
rect 561860 402768 561920 402828
rect 562060 402768 562120 402828
rect 562260 402768 562320 402828
rect 562460 402768 562520 402828
rect 562660 402768 562720 402828
rect 562860 402768 562920 402828
rect 563060 402768 563120 402828
rect 563260 402768 563320 402828
rect 563460 402768 563520 402828
rect 563660 402768 563720 402828
rect 563860 402768 563920 402828
rect 564060 402768 564120 402828
rect 564260 402768 564320 402828
rect 564460 402768 564520 402828
rect 564660 402768 564720 402828
rect 564860 402768 564920 402828
rect 565060 402768 565120 402828
rect 565260 402768 565320 402828
rect 565460 402768 565520 402828
rect 565660 402768 565720 402828
rect 574506 402808 574566 402868
rect 574706 402808 574766 402868
rect 574906 402808 574966 402868
rect 575106 402808 575166 402868
rect 575306 402808 575366 402868
rect 575506 402808 575566 402868
rect 575706 402808 575766 402868
rect 575906 402808 575966 402868
rect 576106 402808 576166 402868
rect 576306 402808 576366 402868
rect 576506 402808 576566 402868
rect 576706 402808 576766 402868
rect 576906 402808 576966 402868
rect 577106 402808 577166 402868
rect 577306 402808 577366 402868
rect 577506 402808 577566 402868
rect 577706 402808 577766 402868
rect 577906 402808 577966 402868
rect 578106 402808 578166 402868
rect 578306 402808 578366 402868
rect 578506 402808 578566 402868
rect 578706 402808 578766 402868
rect 578906 402808 578966 402868
rect 579106 402808 579166 402868
rect 579306 402808 579366 402868
rect 579506 402808 579566 402868
rect 506251 402545 506285 402579
rect 506251 402345 506285 402379
rect 506251 402145 506285 402179
rect 506251 401945 506285 401979
rect 506251 401745 506285 401779
rect 494971 401371 495005 401405
rect 494971 400971 495005 401005
rect 504371 401059 504405 401093
rect 494971 400571 495005 400605
rect 496851 400619 496885 400653
rect 497371 400790 497391 400824
rect 497391 400790 497405 400824
rect 497443 400790 497459 400824
rect 497459 400790 497477 400824
rect 497515 400790 497527 400824
rect 497527 400790 497549 400824
rect 497587 400790 497595 400824
rect 497595 400790 497621 400824
rect 497659 400790 497663 400824
rect 497663 400790 497693 400824
rect 497731 400790 497765 400824
rect 497803 400790 497833 400824
rect 497833 400790 497837 400824
rect 497875 400790 497901 400824
rect 497901 400790 497909 400824
rect 497947 400790 497969 400824
rect 497969 400790 497981 400824
rect 498019 400790 498037 400824
rect 498037 400790 498053 400824
rect 498091 400790 498105 400824
rect 498105 400790 498125 400824
rect 498353 400539 498387 400573
rect 497371 400332 497391 400366
rect 497391 400332 497405 400366
rect 497443 400332 497459 400366
rect 497459 400332 497477 400366
rect 497515 400332 497527 400366
rect 497527 400332 497549 400366
rect 497587 400332 497595 400366
rect 497595 400332 497621 400366
rect 497659 400332 497663 400366
rect 497663 400332 497693 400366
rect 497731 400332 497765 400366
rect 497803 400332 497833 400366
rect 497833 400332 497837 400366
rect 497875 400332 497901 400366
rect 497901 400332 497909 400366
rect 497947 400332 497969 400366
rect 497969 400332 497981 400366
rect 498019 400332 498037 400366
rect 498037 400332 498053 400366
rect 498091 400332 498105 400366
rect 498105 400332 498125 400366
rect 498557 400355 498591 400389
rect 498731 400619 498765 400653
rect 504371 400859 504405 400893
rect 504639 400863 505177 401257
rect 505599 400863 506137 401257
rect 506251 401059 506285 401093
rect 506251 400859 506285 400893
rect 504371 400659 504405 400693
rect 504371 400459 504405 400493
rect 494971 400171 495005 400205
rect 506251 400659 506285 400693
rect 506251 400459 506285 400493
rect 504371 400259 504405 400293
rect 504371 400059 504405 400093
rect 494971 399771 495005 399805
rect 494971 399371 495005 399405
rect 494971 398971 495005 399005
rect 494971 398571 495005 398605
rect 494971 398171 495005 398205
rect 494971 397771 495005 397805
rect 494971 397371 495005 397405
rect 494971 396971 495005 397005
rect 494971 396571 495005 396605
rect 494971 396171 495005 396205
rect 494971 395771 495005 395805
rect 494971 395371 495005 395405
rect 494971 394971 495005 395005
rect 494971 394571 495005 394605
rect 498489 399895 498523 399929
rect 496851 399707 496885 399741
rect 496851 399307 496885 399341
rect 497119 399843 497153 399877
rect 497191 399843 497221 399877
rect 497221 399843 497225 399877
rect 497263 399843 497289 399877
rect 497289 399843 497297 399877
rect 497335 399843 497357 399877
rect 497357 399843 497369 399877
rect 497407 399843 497425 399877
rect 497425 399843 497441 399877
rect 497479 399843 497493 399877
rect 497493 399843 497513 399877
rect 497551 399843 497561 399877
rect 497561 399843 497585 399877
rect 497623 399843 497629 399877
rect 497629 399843 497657 399877
rect 497695 399843 497697 399877
rect 497697 399843 497729 399877
rect 497767 399843 497799 399877
rect 497799 399843 497801 399877
rect 497839 399843 497867 399877
rect 497867 399843 497873 399877
rect 497911 399843 497935 399877
rect 497935 399843 497945 399877
rect 497983 399843 498003 399877
rect 498003 399843 498017 399877
rect 498055 399843 498071 399877
rect 498071 399843 498089 399877
rect 498127 399843 498139 399877
rect 498139 399843 498161 399877
rect 498199 399843 498207 399877
rect 498207 399843 498233 399877
rect 498271 399843 498275 399877
rect 498275 399843 498305 399877
rect 498343 399843 498377 399877
rect 497119 399385 497153 399419
rect 497191 399385 497221 399419
rect 497221 399385 497225 399419
rect 497263 399385 497289 399419
rect 497289 399385 497297 399419
rect 497335 399385 497357 399419
rect 497357 399385 497369 399419
rect 497407 399385 497425 399419
rect 497425 399385 497441 399419
rect 497479 399385 497493 399419
rect 497493 399385 497513 399419
rect 497551 399385 497561 399419
rect 497561 399385 497585 399419
rect 497623 399385 497629 399419
rect 497629 399385 497657 399419
rect 497695 399385 497697 399419
rect 497697 399385 497729 399419
rect 497767 399385 497799 399419
rect 497799 399385 497801 399419
rect 497839 399385 497867 399419
rect 497867 399385 497873 399419
rect 497911 399385 497935 399419
rect 497935 399385 497945 399419
rect 497983 399385 498003 399419
rect 498003 399385 498017 399419
rect 498055 399385 498071 399419
rect 498071 399385 498089 399419
rect 498127 399385 498139 399419
rect 498139 399385 498161 399419
rect 498199 399385 498207 399419
rect 498207 399385 498233 399419
rect 498271 399385 498275 399419
rect 498275 399385 498305 399419
rect 498343 399385 498377 399419
rect 496851 398907 496885 398941
rect 496851 398507 496885 398541
rect 496851 398107 496885 398141
rect 496851 397707 496885 397741
rect 497119 398927 497153 398961
rect 497191 398927 497221 398961
rect 497221 398927 497225 398961
rect 497263 398927 497289 398961
rect 497289 398927 497297 398961
rect 497335 398927 497357 398961
rect 497357 398927 497369 398961
rect 497407 398927 497425 398961
rect 497425 398927 497441 398961
rect 497479 398927 497493 398961
rect 497493 398927 497513 398961
rect 497551 398927 497561 398961
rect 497561 398927 497585 398961
rect 497623 398927 497629 398961
rect 497629 398927 497657 398961
rect 497695 398927 497697 398961
rect 497697 398927 497729 398961
rect 497767 398927 497799 398961
rect 497799 398927 497801 398961
rect 497839 398927 497867 398961
rect 497867 398927 497873 398961
rect 497911 398927 497935 398961
rect 497935 398927 497945 398961
rect 497983 398927 498003 398961
rect 498003 398927 498017 398961
rect 498055 398927 498071 398961
rect 498071 398927 498089 398961
rect 498127 398927 498139 398961
rect 498139 398927 498161 398961
rect 498199 398927 498207 398961
rect 498207 398927 498233 398961
rect 498271 398927 498275 398961
rect 498275 398927 498305 398961
rect 498343 398927 498377 398961
rect 497119 398469 497153 398503
rect 497191 398469 497221 398503
rect 497221 398469 497225 398503
rect 497263 398469 497289 398503
rect 497289 398469 497297 398503
rect 497335 398469 497357 398503
rect 497357 398469 497369 398503
rect 497407 398469 497425 398503
rect 497425 398469 497441 398503
rect 497479 398469 497493 398503
rect 497493 398469 497513 398503
rect 497551 398469 497561 398503
rect 497561 398469 497585 398503
rect 497623 398469 497629 398503
rect 497629 398469 497657 398503
rect 497695 398469 497697 398503
rect 497697 398469 497729 398503
rect 497767 398469 497799 398503
rect 497799 398469 497801 398503
rect 497839 398469 497867 398503
rect 497867 398469 497873 398503
rect 497911 398469 497935 398503
rect 497935 398469 497945 398503
rect 497983 398469 498003 398503
rect 498003 398469 498017 398503
rect 498055 398469 498071 398503
rect 498071 398469 498089 398503
rect 498127 398469 498139 398503
rect 498139 398469 498161 398503
rect 498199 398469 498207 398503
rect 498207 398469 498233 398503
rect 498271 398469 498275 398503
rect 498275 398469 498305 398503
rect 498343 398469 498377 398503
rect 497119 398011 497153 398045
rect 497191 398011 497221 398045
rect 497221 398011 497225 398045
rect 497263 398011 497289 398045
rect 497289 398011 497297 398045
rect 497335 398011 497357 398045
rect 497357 398011 497369 398045
rect 497407 398011 497425 398045
rect 497425 398011 497441 398045
rect 497479 398011 497493 398045
rect 497493 398011 497513 398045
rect 497551 398011 497561 398045
rect 497561 398011 497585 398045
rect 497623 398011 497629 398045
rect 497629 398011 497657 398045
rect 497695 398011 497697 398045
rect 497697 398011 497729 398045
rect 497767 398011 497799 398045
rect 497799 398011 497801 398045
rect 497839 398011 497867 398045
rect 497867 398011 497873 398045
rect 497911 398011 497935 398045
rect 497935 398011 497945 398045
rect 497983 398011 498003 398045
rect 498003 398011 498017 398045
rect 498055 398011 498071 398045
rect 498071 398011 498089 398045
rect 498127 398011 498139 398045
rect 498139 398011 498161 398045
rect 498199 398011 498207 398045
rect 498207 398011 498233 398045
rect 498271 398011 498275 398045
rect 498275 398011 498305 398045
rect 498343 398011 498377 398045
rect 497119 397553 497153 397587
rect 497191 397553 497221 397587
rect 497221 397553 497225 397587
rect 497263 397553 497289 397587
rect 497289 397553 497297 397587
rect 497335 397553 497357 397587
rect 497357 397553 497369 397587
rect 497407 397553 497425 397587
rect 497425 397553 497441 397587
rect 497479 397553 497493 397587
rect 497493 397553 497513 397587
rect 497551 397553 497561 397587
rect 497561 397553 497585 397587
rect 497623 397553 497629 397587
rect 497629 397553 497657 397587
rect 497695 397553 497697 397587
rect 497697 397553 497729 397587
rect 497767 397553 497799 397587
rect 497799 397553 497801 397587
rect 497839 397553 497867 397587
rect 497867 397553 497873 397587
rect 497911 397553 497935 397587
rect 497935 397553 497945 397587
rect 497983 397553 498003 397587
rect 498003 397553 498017 397587
rect 498055 397553 498071 397587
rect 498071 397553 498089 397587
rect 498127 397553 498139 397587
rect 498139 397553 498161 397587
rect 498199 397553 498207 397587
rect 498207 397553 498233 397587
rect 498271 397553 498275 397587
rect 498275 397553 498305 397587
rect 498343 397553 498377 397587
rect 496851 397307 496885 397341
rect 496851 396907 496885 396941
rect 496851 396507 496885 396541
rect 497119 397095 497153 397129
rect 497191 397095 497221 397129
rect 497221 397095 497225 397129
rect 497263 397095 497289 397129
rect 497289 397095 497297 397129
rect 497335 397095 497357 397129
rect 497357 397095 497369 397129
rect 497407 397095 497425 397129
rect 497425 397095 497441 397129
rect 497479 397095 497493 397129
rect 497493 397095 497513 397129
rect 497551 397095 497561 397129
rect 497561 397095 497585 397129
rect 497623 397095 497629 397129
rect 497629 397095 497657 397129
rect 497695 397095 497697 397129
rect 497697 397095 497729 397129
rect 497767 397095 497799 397129
rect 497799 397095 497801 397129
rect 497839 397095 497867 397129
rect 497867 397095 497873 397129
rect 497911 397095 497935 397129
rect 497935 397095 497945 397129
rect 497983 397095 498003 397129
rect 498003 397095 498017 397129
rect 498055 397095 498071 397129
rect 498071 397095 498089 397129
rect 498127 397095 498139 397129
rect 498139 397095 498161 397129
rect 498199 397095 498207 397129
rect 498207 397095 498233 397129
rect 498271 397095 498275 397129
rect 498275 397095 498305 397129
rect 498343 397095 498377 397129
rect 497119 396637 497153 396671
rect 497191 396637 497221 396671
rect 497221 396637 497225 396671
rect 497263 396637 497289 396671
rect 497289 396637 497297 396671
rect 497335 396637 497357 396671
rect 497357 396637 497369 396671
rect 497407 396637 497425 396671
rect 497425 396637 497441 396671
rect 497479 396637 497493 396671
rect 497493 396637 497513 396671
rect 497551 396637 497561 396671
rect 497561 396637 497585 396671
rect 497623 396637 497629 396671
rect 497629 396637 497657 396671
rect 497695 396637 497697 396671
rect 497697 396637 497729 396671
rect 497767 396637 497799 396671
rect 497799 396637 497801 396671
rect 497839 396637 497867 396671
rect 497867 396637 497873 396671
rect 497911 396637 497935 396671
rect 497935 396637 497945 396671
rect 497983 396637 498003 396671
rect 498003 396637 498017 396671
rect 498055 396637 498071 396671
rect 498071 396637 498089 396671
rect 498127 396637 498139 396671
rect 498139 396637 498161 396671
rect 498199 396637 498207 396671
rect 498207 396637 498233 396671
rect 498271 396637 498275 396671
rect 498275 396637 498305 396671
rect 498343 396637 498377 396671
rect 496851 396107 496885 396141
rect 496851 395707 496885 395741
rect 496851 395307 496885 395341
rect 497119 396179 497153 396213
rect 497191 396179 497221 396213
rect 497221 396179 497225 396213
rect 497263 396179 497289 396213
rect 497289 396179 497297 396213
rect 497335 396179 497357 396213
rect 497357 396179 497369 396213
rect 497407 396179 497425 396213
rect 497425 396179 497441 396213
rect 497479 396179 497493 396213
rect 497493 396179 497513 396213
rect 497551 396179 497561 396213
rect 497561 396179 497585 396213
rect 497623 396179 497629 396213
rect 497629 396179 497657 396213
rect 497695 396179 497697 396213
rect 497697 396179 497729 396213
rect 497767 396179 497799 396213
rect 497799 396179 497801 396213
rect 497839 396179 497867 396213
rect 497867 396179 497873 396213
rect 497911 396179 497935 396213
rect 497935 396179 497945 396213
rect 497983 396179 498003 396213
rect 498003 396179 498017 396213
rect 498055 396179 498071 396213
rect 498071 396179 498089 396213
rect 498127 396179 498139 396213
rect 498139 396179 498161 396213
rect 498199 396179 498207 396213
rect 498207 396179 498233 396213
rect 498271 396179 498275 396213
rect 498275 396179 498305 396213
rect 498343 396179 498377 396213
rect 497119 395721 497153 395755
rect 497191 395721 497221 395755
rect 497221 395721 497225 395755
rect 497263 395721 497289 395755
rect 497289 395721 497297 395755
rect 497335 395721 497357 395755
rect 497357 395721 497369 395755
rect 497407 395721 497425 395755
rect 497425 395721 497441 395755
rect 497479 395721 497493 395755
rect 497493 395721 497513 395755
rect 497551 395721 497561 395755
rect 497561 395721 497585 395755
rect 497623 395721 497629 395755
rect 497629 395721 497657 395755
rect 497695 395721 497697 395755
rect 497697 395721 497729 395755
rect 497767 395721 497799 395755
rect 497799 395721 497801 395755
rect 497839 395721 497867 395755
rect 497867 395721 497873 395755
rect 497911 395721 497935 395755
rect 497935 395721 497945 395755
rect 497983 395721 498003 395755
rect 498003 395721 498017 395755
rect 498055 395721 498071 395755
rect 498071 395721 498089 395755
rect 498127 395721 498139 395755
rect 498139 395721 498161 395755
rect 498199 395721 498207 395755
rect 498207 395721 498233 395755
rect 498271 395721 498275 395755
rect 498275 395721 498305 395755
rect 498343 395721 498377 395755
rect 496851 394907 496885 394941
rect 496851 394507 496885 394541
rect 493091 393905 493125 393939
rect 493091 393705 493125 393739
rect 493359 393709 493897 394103
rect 494319 393709 494857 394103
rect 494971 393905 495005 393939
rect 494971 393705 495005 393739
rect 493091 393505 493125 393539
rect 493091 393305 493125 393339
rect 494971 393505 495005 393539
rect 494971 393305 495005 393339
rect 493091 393105 493125 393139
rect 493091 392905 493125 392939
rect 493091 392705 493125 392739
rect 494971 393105 495005 393139
rect 494971 392905 495005 392939
rect 494971 392705 495005 392739
rect 493091 392505 493125 392539
rect 493091 392305 493125 392339
rect 493091 392105 493125 392139
rect 494971 392505 495005 392539
rect 494971 392305 495005 392339
rect 493091 391905 493125 391939
rect 493359 391702 493897 392096
rect 494319 391702 494857 392096
rect 494971 392105 495005 392139
rect 494971 391905 495005 391939
rect 496851 394107 496885 394141
rect 497119 395263 497153 395297
rect 497191 395263 497221 395297
rect 497221 395263 497225 395297
rect 497263 395263 497289 395297
rect 497289 395263 497297 395297
rect 497335 395263 497357 395297
rect 497357 395263 497369 395297
rect 497407 395263 497425 395297
rect 497425 395263 497441 395297
rect 497479 395263 497493 395297
rect 497493 395263 497513 395297
rect 497551 395263 497561 395297
rect 497561 395263 497585 395297
rect 497623 395263 497629 395297
rect 497629 395263 497657 395297
rect 497695 395263 497697 395297
rect 497697 395263 497729 395297
rect 497767 395263 497799 395297
rect 497799 395263 497801 395297
rect 497839 395263 497867 395297
rect 497867 395263 497873 395297
rect 497911 395263 497935 395297
rect 497935 395263 497945 395297
rect 497983 395263 498003 395297
rect 498003 395263 498017 395297
rect 498055 395263 498071 395297
rect 498071 395263 498089 395297
rect 498127 395263 498139 395297
rect 498139 395263 498161 395297
rect 498199 395263 498207 395297
rect 498207 395263 498233 395297
rect 498271 395263 498275 395297
rect 498275 395263 498305 395297
rect 498343 395263 498377 395297
rect 497119 394805 497153 394839
rect 497191 394805 497221 394839
rect 497221 394805 497225 394839
rect 497263 394805 497289 394839
rect 497289 394805 497297 394839
rect 497335 394805 497357 394839
rect 497357 394805 497369 394839
rect 497407 394805 497425 394839
rect 497425 394805 497441 394839
rect 497479 394805 497493 394839
rect 497493 394805 497513 394839
rect 497551 394805 497561 394839
rect 497561 394805 497585 394839
rect 497623 394805 497629 394839
rect 497629 394805 497657 394839
rect 497695 394805 497697 394839
rect 497697 394805 497729 394839
rect 497767 394805 497799 394839
rect 497799 394805 497801 394839
rect 497839 394805 497867 394839
rect 497867 394805 497873 394839
rect 497911 394805 497935 394839
rect 497935 394805 497945 394839
rect 497983 394805 498003 394839
rect 498003 394805 498017 394839
rect 498055 394805 498071 394839
rect 498071 394805 498089 394839
rect 498127 394805 498139 394839
rect 498139 394805 498161 394839
rect 498199 394805 498207 394839
rect 498207 394805 498233 394839
rect 498271 394805 498275 394839
rect 498275 394805 498305 394839
rect 498343 394805 498377 394839
rect 497119 394347 497153 394381
rect 497191 394347 497221 394381
rect 497221 394347 497225 394381
rect 497263 394347 497289 394381
rect 497289 394347 497297 394381
rect 497335 394347 497357 394381
rect 497357 394347 497369 394381
rect 497407 394347 497425 394381
rect 497425 394347 497441 394381
rect 497479 394347 497493 394381
rect 497493 394347 497513 394381
rect 497551 394347 497561 394381
rect 497561 394347 497585 394381
rect 497623 394347 497629 394381
rect 497629 394347 497657 394381
rect 497695 394347 497697 394381
rect 497697 394347 497729 394381
rect 497767 394347 497799 394381
rect 497799 394347 497801 394381
rect 497839 394347 497867 394381
rect 497867 394347 497873 394381
rect 497911 394347 497935 394381
rect 497935 394347 497945 394381
rect 497983 394347 498003 394381
rect 498003 394347 498017 394381
rect 498055 394347 498071 394381
rect 498071 394347 498089 394381
rect 498127 394347 498139 394381
rect 498139 394347 498161 394381
rect 498199 394347 498207 394381
rect 498207 394347 498233 394381
rect 498271 394347 498275 394381
rect 498275 394347 498305 394381
rect 498343 394347 498377 394381
rect 497119 393889 497153 393923
rect 497191 393889 497221 393923
rect 497221 393889 497225 393923
rect 497263 393889 497289 393923
rect 497289 393889 497297 393923
rect 497335 393889 497357 393923
rect 497357 393889 497369 393923
rect 497407 393889 497425 393923
rect 497425 393889 497441 393923
rect 497479 393889 497493 393923
rect 497493 393889 497513 393923
rect 497551 393889 497561 393923
rect 497561 393889 497585 393923
rect 497623 393889 497629 393923
rect 497629 393889 497657 393923
rect 497695 393889 497697 393923
rect 497697 393889 497729 393923
rect 497767 393889 497799 393923
rect 497799 393889 497801 393923
rect 497839 393889 497867 393923
rect 497867 393889 497873 393923
rect 497911 393889 497935 393923
rect 497935 393889 497945 393923
rect 497983 393889 498003 393923
rect 498003 393889 498017 393923
rect 498055 393889 498071 393923
rect 498071 393889 498089 393923
rect 498127 393889 498139 393923
rect 498139 393889 498161 393923
rect 498199 393889 498207 393923
rect 498207 393889 498233 393923
rect 498271 393889 498275 393923
rect 498275 393889 498305 393923
rect 498343 393889 498377 393923
rect 496851 393707 496885 393741
rect 496851 393307 496885 393341
rect 496851 392907 496885 392941
rect 496851 392507 496885 392541
rect 497119 393431 497153 393465
rect 497191 393431 497221 393465
rect 497221 393431 497225 393465
rect 497263 393431 497289 393465
rect 497289 393431 497297 393465
rect 497335 393431 497357 393465
rect 497357 393431 497369 393465
rect 497407 393431 497425 393465
rect 497425 393431 497441 393465
rect 497479 393431 497493 393465
rect 497493 393431 497513 393465
rect 497551 393431 497561 393465
rect 497561 393431 497585 393465
rect 497623 393431 497629 393465
rect 497629 393431 497657 393465
rect 497695 393431 497697 393465
rect 497697 393431 497729 393465
rect 497767 393431 497799 393465
rect 497799 393431 497801 393465
rect 497839 393431 497867 393465
rect 497867 393431 497873 393465
rect 497911 393431 497935 393465
rect 497935 393431 497945 393465
rect 497983 393431 498003 393465
rect 498003 393431 498017 393465
rect 498055 393431 498071 393465
rect 498071 393431 498089 393465
rect 498127 393431 498139 393465
rect 498139 393431 498161 393465
rect 498199 393431 498207 393465
rect 498207 393431 498233 393465
rect 498271 393431 498275 393465
rect 498275 393431 498305 393465
rect 498343 393431 498377 393465
rect 497119 392973 497153 393007
rect 497191 392973 497221 393007
rect 497221 392973 497225 393007
rect 497263 392973 497289 393007
rect 497289 392973 497297 393007
rect 497335 392973 497357 393007
rect 497357 392973 497369 393007
rect 497407 392973 497425 393007
rect 497425 392973 497441 393007
rect 497479 392973 497493 393007
rect 497493 392973 497513 393007
rect 497551 392973 497561 393007
rect 497561 392973 497585 393007
rect 497623 392973 497629 393007
rect 497629 392973 497657 393007
rect 497695 392973 497697 393007
rect 497697 392973 497729 393007
rect 497767 392973 497799 393007
rect 497799 392973 497801 393007
rect 497839 392973 497867 393007
rect 497867 392973 497873 393007
rect 497911 392973 497935 393007
rect 497935 392973 497945 393007
rect 497983 392973 498003 393007
rect 498003 392973 498017 393007
rect 498055 392973 498071 393007
rect 498071 392973 498089 393007
rect 498127 392973 498139 393007
rect 498139 392973 498161 393007
rect 498199 392973 498207 393007
rect 498207 392973 498233 393007
rect 498271 392973 498275 393007
rect 498275 392973 498305 393007
rect 498343 392973 498377 393007
rect 496851 392107 496885 392141
rect 496851 391707 496885 391741
rect 496851 391307 496885 391341
rect 497119 392515 497153 392549
rect 497191 392515 497221 392549
rect 497221 392515 497225 392549
rect 497263 392515 497289 392549
rect 497289 392515 497297 392549
rect 497335 392515 497357 392549
rect 497357 392515 497369 392549
rect 497407 392515 497425 392549
rect 497425 392515 497441 392549
rect 497479 392515 497493 392549
rect 497493 392515 497513 392549
rect 497551 392515 497561 392549
rect 497561 392515 497585 392549
rect 497623 392515 497629 392549
rect 497629 392515 497657 392549
rect 497695 392515 497697 392549
rect 497697 392515 497729 392549
rect 497767 392515 497799 392549
rect 497799 392515 497801 392549
rect 497839 392515 497867 392549
rect 497867 392515 497873 392549
rect 497911 392515 497935 392549
rect 497935 392515 497945 392549
rect 497983 392515 498003 392549
rect 498003 392515 498017 392549
rect 498055 392515 498071 392549
rect 498071 392515 498089 392549
rect 498127 392515 498139 392549
rect 498139 392515 498161 392549
rect 498199 392515 498207 392549
rect 498207 392515 498233 392549
rect 498271 392515 498275 392549
rect 498275 392515 498305 392549
rect 498343 392515 498377 392549
rect 497119 392057 497153 392091
rect 497191 392057 497221 392091
rect 497221 392057 497225 392091
rect 497263 392057 497289 392091
rect 497289 392057 497297 392091
rect 497335 392057 497357 392091
rect 497357 392057 497369 392091
rect 497407 392057 497425 392091
rect 497425 392057 497441 392091
rect 497479 392057 497493 392091
rect 497493 392057 497513 392091
rect 497551 392057 497561 392091
rect 497561 392057 497585 392091
rect 497623 392057 497629 392091
rect 497629 392057 497657 392091
rect 497695 392057 497697 392091
rect 497697 392057 497729 392091
rect 497767 392057 497799 392091
rect 497799 392057 497801 392091
rect 497839 392057 497867 392091
rect 497867 392057 497873 392091
rect 497911 392057 497935 392091
rect 497935 392057 497945 392091
rect 497983 392057 498003 392091
rect 498003 392057 498017 392091
rect 498055 392057 498071 392091
rect 498071 392057 498089 392091
rect 498127 392057 498139 392091
rect 498139 392057 498161 392091
rect 498199 392057 498207 392091
rect 498207 392057 498233 392091
rect 498271 392057 498275 392091
rect 498275 392057 498305 392091
rect 498343 392057 498377 392091
rect 497119 391599 497153 391633
rect 497191 391599 497221 391633
rect 497221 391599 497225 391633
rect 497263 391599 497289 391633
rect 497289 391599 497297 391633
rect 497335 391599 497357 391633
rect 497357 391599 497369 391633
rect 497407 391599 497425 391633
rect 497425 391599 497441 391633
rect 497479 391599 497493 391633
rect 497493 391599 497513 391633
rect 497551 391599 497561 391633
rect 497561 391599 497585 391633
rect 497623 391599 497629 391633
rect 497629 391599 497657 391633
rect 497695 391599 497697 391633
rect 497697 391599 497729 391633
rect 497767 391599 497799 391633
rect 497799 391599 497801 391633
rect 497839 391599 497867 391633
rect 497867 391599 497873 391633
rect 497911 391599 497935 391633
rect 497935 391599 497945 391633
rect 497983 391599 498003 391633
rect 498003 391599 498017 391633
rect 498055 391599 498071 391633
rect 498071 391599 498089 391633
rect 498127 391599 498139 391633
rect 498139 391599 498161 391633
rect 498199 391599 498207 391633
rect 498207 391599 498233 391633
rect 498271 391599 498275 391633
rect 498275 391599 498305 391633
rect 498343 391599 498377 391633
rect 493091 390819 493125 390853
rect 493611 390990 493631 391024
rect 493631 390990 493645 391024
rect 493683 390990 493699 391024
rect 493699 390990 493717 391024
rect 493755 390990 493767 391024
rect 493767 390990 493789 391024
rect 493827 390990 493835 391024
rect 493835 390990 493861 391024
rect 493899 390990 493903 391024
rect 493903 390990 493933 391024
rect 493971 390990 494005 391024
rect 494043 390990 494073 391024
rect 494073 390990 494077 391024
rect 494115 390990 494141 391024
rect 494141 390990 494149 391024
rect 494187 390990 494209 391024
rect 494209 390990 494221 391024
rect 494259 390990 494277 391024
rect 494277 390990 494293 391024
rect 494331 390990 494345 391024
rect 494345 390990 494365 391024
rect 493611 390532 493631 390566
rect 493631 390532 493645 390566
rect 493683 390532 493699 390566
rect 493699 390532 493717 390566
rect 493755 390532 493767 390566
rect 493767 390532 493789 390566
rect 493827 390532 493835 390566
rect 493835 390532 493861 390566
rect 493899 390532 493903 390566
rect 493903 390532 493933 390566
rect 493971 390532 494005 390566
rect 494043 390532 494073 390566
rect 494073 390532 494077 390566
rect 494115 390532 494141 390566
rect 494141 390532 494149 390566
rect 494187 390532 494209 390566
rect 494209 390532 494221 390566
rect 494259 390532 494277 390566
rect 494277 390532 494293 390566
rect 494331 390532 494345 390566
rect 494345 390532 494365 390566
rect 494817 390879 494851 390913
rect 494971 390819 495005 390853
rect 497119 391141 497153 391175
rect 497191 391141 497221 391175
rect 497221 391141 497225 391175
rect 497263 391141 497289 391175
rect 497289 391141 497297 391175
rect 497335 391141 497357 391175
rect 497357 391141 497369 391175
rect 497407 391141 497425 391175
rect 497425 391141 497441 391175
rect 497479 391141 497493 391175
rect 497493 391141 497513 391175
rect 497551 391141 497561 391175
rect 497561 391141 497585 391175
rect 497623 391141 497629 391175
rect 497629 391141 497657 391175
rect 497695 391141 497697 391175
rect 497697 391141 497729 391175
rect 497767 391141 497799 391175
rect 497799 391141 497801 391175
rect 497839 391141 497867 391175
rect 497867 391141 497873 391175
rect 497911 391141 497935 391175
rect 497935 391141 497945 391175
rect 497983 391141 498003 391175
rect 498003 391141 498017 391175
rect 498055 391141 498071 391175
rect 498071 391141 498089 391175
rect 498127 391141 498139 391175
rect 498139 391141 498161 391175
rect 498199 391141 498207 391175
rect 498207 391141 498233 391175
rect 498271 391141 498275 391175
rect 498275 391141 498305 391175
rect 498343 391141 498377 391175
rect 496851 390907 496885 390941
rect 496851 390507 496885 390541
rect 493091 389907 493125 389941
rect 493091 389507 493125 389541
rect 493359 390043 493393 390077
rect 493431 390043 493461 390077
rect 493461 390043 493465 390077
rect 493503 390043 493529 390077
rect 493529 390043 493537 390077
rect 493575 390043 493597 390077
rect 493597 390043 493609 390077
rect 493647 390043 493665 390077
rect 493665 390043 493681 390077
rect 493719 390043 493733 390077
rect 493733 390043 493753 390077
rect 493791 390043 493801 390077
rect 493801 390043 493825 390077
rect 493863 390043 493869 390077
rect 493869 390043 493897 390077
rect 493935 390043 493937 390077
rect 493937 390043 493969 390077
rect 494007 390043 494039 390077
rect 494039 390043 494041 390077
rect 494079 390043 494107 390077
rect 494107 390043 494113 390077
rect 494151 390043 494175 390077
rect 494175 390043 494185 390077
rect 494223 390043 494243 390077
rect 494243 390043 494257 390077
rect 494295 390043 494311 390077
rect 494311 390043 494329 390077
rect 494367 390043 494379 390077
rect 494379 390043 494401 390077
rect 494439 390043 494447 390077
rect 494447 390043 494473 390077
rect 494511 390043 494515 390077
rect 494515 390043 494545 390077
rect 494583 390043 494617 390077
rect 493359 389585 493393 389619
rect 493431 389585 493461 389619
rect 493461 389585 493465 389619
rect 493503 389585 493529 389619
rect 493529 389585 493537 389619
rect 493575 389585 493597 389619
rect 493597 389585 493609 389619
rect 493647 389585 493665 389619
rect 493665 389585 493681 389619
rect 493719 389585 493733 389619
rect 493733 389585 493753 389619
rect 493791 389585 493801 389619
rect 493801 389585 493825 389619
rect 493863 389585 493869 389619
rect 493869 389585 493897 389619
rect 493935 389585 493937 389619
rect 493937 389585 493969 389619
rect 494007 389585 494039 389619
rect 494039 389585 494041 389619
rect 494079 389585 494107 389619
rect 494107 389585 494113 389619
rect 494151 389585 494175 389619
rect 494175 389585 494185 389619
rect 494223 389585 494243 389619
rect 494243 389585 494257 389619
rect 494295 389585 494311 389619
rect 494311 389585 494329 389619
rect 494367 389585 494379 389619
rect 494379 389585 494401 389619
rect 494439 389585 494447 389619
rect 494447 389585 494473 389619
rect 494511 389585 494515 389619
rect 494515 389585 494545 389619
rect 494583 389585 494617 389619
rect 493091 389107 493125 389141
rect 493091 388707 493125 388741
rect 493091 388307 493125 388341
rect 493091 387907 493125 387941
rect 493359 389127 493393 389161
rect 493431 389127 493461 389161
rect 493461 389127 493465 389161
rect 493503 389127 493529 389161
rect 493529 389127 493537 389161
rect 493575 389127 493597 389161
rect 493597 389127 493609 389161
rect 493647 389127 493665 389161
rect 493665 389127 493681 389161
rect 493719 389127 493733 389161
rect 493733 389127 493753 389161
rect 493791 389127 493801 389161
rect 493801 389127 493825 389161
rect 493863 389127 493869 389161
rect 493869 389127 493897 389161
rect 493935 389127 493937 389161
rect 493937 389127 493969 389161
rect 494007 389127 494039 389161
rect 494039 389127 494041 389161
rect 494079 389127 494107 389161
rect 494107 389127 494113 389161
rect 494151 389127 494175 389161
rect 494175 389127 494185 389161
rect 494223 389127 494243 389161
rect 494243 389127 494257 389161
rect 494295 389127 494311 389161
rect 494311 389127 494329 389161
rect 494367 389127 494379 389161
rect 494379 389127 494401 389161
rect 494439 389127 494447 389161
rect 494447 389127 494473 389161
rect 494511 389127 494515 389161
rect 494515 389127 494545 389161
rect 494583 389127 494617 389161
rect 493359 388669 493393 388703
rect 493431 388669 493461 388703
rect 493461 388669 493465 388703
rect 493503 388669 493529 388703
rect 493529 388669 493537 388703
rect 493575 388669 493597 388703
rect 493597 388669 493609 388703
rect 493647 388669 493665 388703
rect 493665 388669 493681 388703
rect 493719 388669 493733 388703
rect 493733 388669 493753 388703
rect 493791 388669 493801 388703
rect 493801 388669 493825 388703
rect 493863 388669 493869 388703
rect 493869 388669 493897 388703
rect 493935 388669 493937 388703
rect 493937 388669 493969 388703
rect 494007 388669 494039 388703
rect 494039 388669 494041 388703
rect 494079 388669 494107 388703
rect 494107 388669 494113 388703
rect 494151 388669 494175 388703
rect 494175 388669 494185 388703
rect 494223 388669 494243 388703
rect 494243 388669 494257 388703
rect 494295 388669 494311 388703
rect 494311 388669 494329 388703
rect 494367 388669 494379 388703
rect 494379 388669 494401 388703
rect 494439 388669 494447 388703
rect 494447 388669 494473 388703
rect 494511 388669 494515 388703
rect 494515 388669 494545 388703
rect 494583 388669 494617 388703
rect 493359 388211 493393 388245
rect 493431 388211 493461 388245
rect 493461 388211 493465 388245
rect 493503 388211 493529 388245
rect 493529 388211 493537 388245
rect 493575 388211 493597 388245
rect 493597 388211 493609 388245
rect 493647 388211 493665 388245
rect 493665 388211 493681 388245
rect 493719 388211 493733 388245
rect 493733 388211 493753 388245
rect 493791 388211 493801 388245
rect 493801 388211 493825 388245
rect 493863 388211 493869 388245
rect 493869 388211 493897 388245
rect 493935 388211 493937 388245
rect 493937 388211 493969 388245
rect 494007 388211 494039 388245
rect 494039 388211 494041 388245
rect 494079 388211 494107 388245
rect 494107 388211 494113 388245
rect 494151 388211 494175 388245
rect 494175 388211 494185 388245
rect 494223 388211 494243 388245
rect 494243 388211 494257 388245
rect 494295 388211 494311 388245
rect 494311 388211 494329 388245
rect 494367 388211 494379 388245
rect 494379 388211 494401 388245
rect 494439 388211 494447 388245
rect 494447 388211 494473 388245
rect 494511 388211 494515 388245
rect 494515 388211 494545 388245
rect 494583 388211 494617 388245
rect 493359 387753 493393 387787
rect 493431 387753 493461 387787
rect 493461 387753 493465 387787
rect 493503 387753 493529 387787
rect 493529 387753 493537 387787
rect 493575 387753 493597 387787
rect 493597 387753 493609 387787
rect 493647 387753 493665 387787
rect 493665 387753 493681 387787
rect 493719 387753 493733 387787
rect 493733 387753 493753 387787
rect 493791 387753 493801 387787
rect 493801 387753 493825 387787
rect 493863 387753 493869 387787
rect 493869 387753 493897 387787
rect 493935 387753 493937 387787
rect 493937 387753 493969 387787
rect 494007 387753 494039 387787
rect 494039 387753 494041 387787
rect 494079 387753 494107 387787
rect 494107 387753 494113 387787
rect 494151 387753 494175 387787
rect 494175 387753 494185 387787
rect 494223 387753 494243 387787
rect 494243 387753 494257 387787
rect 494295 387753 494311 387787
rect 494311 387753 494329 387787
rect 494367 387753 494379 387787
rect 494379 387753 494401 387787
rect 494439 387753 494447 387787
rect 494447 387753 494473 387787
rect 494511 387753 494515 387787
rect 494515 387753 494545 387787
rect 494583 387753 494617 387787
rect 493091 387507 493125 387541
rect 493091 387107 493125 387141
rect 493091 386707 493125 386741
rect 493359 387295 493393 387329
rect 493431 387295 493461 387329
rect 493461 387295 493465 387329
rect 493503 387295 493529 387329
rect 493529 387295 493537 387329
rect 493575 387295 493597 387329
rect 493597 387295 493609 387329
rect 493647 387295 493665 387329
rect 493665 387295 493681 387329
rect 493719 387295 493733 387329
rect 493733 387295 493753 387329
rect 493791 387295 493801 387329
rect 493801 387295 493825 387329
rect 493863 387295 493869 387329
rect 493869 387295 493897 387329
rect 493935 387295 493937 387329
rect 493937 387295 493969 387329
rect 494007 387295 494039 387329
rect 494039 387295 494041 387329
rect 494079 387295 494107 387329
rect 494107 387295 494113 387329
rect 494151 387295 494175 387329
rect 494175 387295 494185 387329
rect 494223 387295 494243 387329
rect 494243 387295 494257 387329
rect 494295 387295 494311 387329
rect 494311 387295 494329 387329
rect 494367 387295 494379 387329
rect 494379 387295 494401 387329
rect 494439 387295 494447 387329
rect 494447 387295 494473 387329
rect 494511 387295 494515 387329
rect 494515 387295 494545 387329
rect 494583 387295 494617 387329
rect 493359 386837 493393 386871
rect 493431 386837 493461 386871
rect 493461 386837 493465 386871
rect 493503 386837 493529 386871
rect 493529 386837 493537 386871
rect 493575 386837 493597 386871
rect 493597 386837 493609 386871
rect 493647 386837 493665 386871
rect 493665 386837 493681 386871
rect 493719 386837 493733 386871
rect 493733 386837 493753 386871
rect 493791 386837 493801 386871
rect 493801 386837 493825 386871
rect 493863 386837 493869 386871
rect 493869 386837 493897 386871
rect 493935 386837 493937 386871
rect 493937 386837 493969 386871
rect 494007 386837 494039 386871
rect 494039 386837 494041 386871
rect 494079 386837 494107 386871
rect 494107 386837 494113 386871
rect 494151 386837 494175 386871
rect 494175 386837 494185 386871
rect 494223 386837 494243 386871
rect 494243 386837 494257 386871
rect 494295 386837 494311 386871
rect 494311 386837 494329 386871
rect 494367 386837 494379 386871
rect 494379 386837 494401 386871
rect 494439 386837 494447 386871
rect 494447 386837 494473 386871
rect 494511 386837 494515 386871
rect 494515 386837 494545 386871
rect 494583 386837 494617 386871
rect 493091 386307 493125 386341
rect 493091 385907 493125 385941
rect 493091 385507 493125 385541
rect 493359 386379 493393 386413
rect 493431 386379 493461 386413
rect 493461 386379 493465 386413
rect 493503 386379 493529 386413
rect 493529 386379 493537 386413
rect 493575 386379 493597 386413
rect 493597 386379 493609 386413
rect 493647 386379 493665 386413
rect 493665 386379 493681 386413
rect 493719 386379 493733 386413
rect 493733 386379 493753 386413
rect 493791 386379 493801 386413
rect 493801 386379 493825 386413
rect 493863 386379 493869 386413
rect 493869 386379 493897 386413
rect 493935 386379 493937 386413
rect 493937 386379 493969 386413
rect 494007 386379 494039 386413
rect 494039 386379 494041 386413
rect 494079 386379 494107 386413
rect 494107 386379 494113 386413
rect 494151 386379 494175 386413
rect 494175 386379 494185 386413
rect 494223 386379 494243 386413
rect 494243 386379 494257 386413
rect 494295 386379 494311 386413
rect 494311 386379 494329 386413
rect 494367 386379 494379 386413
rect 494379 386379 494401 386413
rect 494439 386379 494447 386413
rect 494447 386379 494473 386413
rect 494511 386379 494515 386413
rect 494515 386379 494545 386413
rect 494583 386379 494617 386413
rect 493359 385921 493393 385955
rect 493431 385921 493461 385955
rect 493461 385921 493465 385955
rect 493503 385921 493529 385955
rect 493529 385921 493537 385955
rect 493575 385921 493597 385955
rect 493597 385921 493609 385955
rect 493647 385921 493665 385955
rect 493665 385921 493681 385955
rect 493719 385921 493733 385955
rect 493733 385921 493753 385955
rect 493791 385921 493801 385955
rect 493801 385921 493825 385955
rect 493863 385921 493869 385955
rect 493869 385921 493897 385955
rect 493935 385921 493937 385955
rect 493937 385921 493969 385955
rect 494007 385921 494039 385955
rect 494039 385921 494041 385955
rect 494079 385921 494107 385955
rect 494107 385921 494113 385955
rect 494151 385921 494175 385955
rect 494175 385921 494185 385955
rect 494223 385921 494243 385955
rect 494243 385921 494257 385955
rect 494295 385921 494311 385955
rect 494311 385921 494329 385955
rect 494367 385921 494379 385955
rect 494379 385921 494401 385955
rect 494439 385921 494447 385955
rect 494447 385921 494473 385955
rect 494511 385921 494515 385955
rect 494515 385921 494545 385955
rect 494583 385921 494617 385955
rect 493091 385107 493125 385141
rect 493091 384707 493125 384741
rect 493091 384307 493125 384341
rect 493359 385463 493393 385497
rect 493431 385463 493461 385497
rect 493461 385463 493465 385497
rect 493503 385463 493529 385497
rect 493529 385463 493537 385497
rect 493575 385463 493597 385497
rect 493597 385463 493609 385497
rect 493647 385463 493665 385497
rect 493665 385463 493681 385497
rect 493719 385463 493733 385497
rect 493733 385463 493753 385497
rect 493791 385463 493801 385497
rect 493801 385463 493825 385497
rect 493863 385463 493869 385497
rect 493869 385463 493897 385497
rect 493935 385463 493937 385497
rect 493937 385463 493969 385497
rect 494007 385463 494039 385497
rect 494039 385463 494041 385497
rect 494079 385463 494107 385497
rect 494107 385463 494113 385497
rect 494151 385463 494175 385497
rect 494175 385463 494185 385497
rect 494223 385463 494243 385497
rect 494243 385463 494257 385497
rect 494295 385463 494311 385497
rect 494311 385463 494329 385497
rect 494367 385463 494379 385497
rect 494379 385463 494401 385497
rect 494439 385463 494447 385497
rect 494447 385463 494473 385497
rect 494511 385463 494515 385497
rect 494515 385463 494545 385497
rect 494583 385463 494617 385497
rect 493359 385005 493393 385039
rect 493431 385005 493461 385039
rect 493461 385005 493465 385039
rect 493503 385005 493529 385039
rect 493529 385005 493537 385039
rect 493575 385005 493597 385039
rect 493597 385005 493609 385039
rect 493647 385005 493665 385039
rect 493665 385005 493681 385039
rect 493719 385005 493733 385039
rect 493733 385005 493753 385039
rect 493791 385005 493801 385039
rect 493801 385005 493825 385039
rect 493863 385005 493869 385039
rect 493869 385005 493897 385039
rect 493935 385005 493937 385039
rect 493937 385005 493969 385039
rect 494007 385005 494039 385039
rect 494039 385005 494041 385039
rect 494079 385005 494107 385039
rect 494107 385005 494113 385039
rect 494151 385005 494175 385039
rect 494175 385005 494185 385039
rect 494223 385005 494243 385039
rect 494243 385005 494257 385039
rect 494295 385005 494311 385039
rect 494311 385005 494329 385039
rect 494367 385005 494379 385039
rect 494379 385005 494401 385039
rect 494439 385005 494447 385039
rect 494447 385005 494473 385039
rect 494511 385005 494515 385039
rect 494515 385005 494545 385039
rect 494583 385005 494617 385039
rect 494817 385451 494851 385485
rect 493359 384547 493393 384581
rect 493431 384547 493461 384581
rect 493461 384547 493465 384581
rect 493503 384547 493529 384581
rect 493529 384547 493537 384581
rect 493575 384547 493597 384581
rect 493597 384547 493609 384581
rect 493647 384547 493665 384581
rect 493665 384547 493681 384581
rect 493719 384547 493733 384581
rect 493733 384547 493753 384581
rect 493791 384547 493801 384581
rect 493801 384547 493825 384581
rect 493863 384547 493869 384581
rect 493869 384547 493897 384581
rect 493935 384547 493937 384581
rect 493937 384547 493969 384581
rect 494007 384547 494039 384581
rect 494039 384547 494041 384581
rect 494079 384547 494107 384581
rect 494107 384547 494113 384581
rect 494151 384547 494175 384581
rect 494175 384547 494185 384581
rect 494223 384547 494243 384581
rect 494243 384547 494257 384581
rect 494295 384547 494311 384581
rect 494311 384547 494329 384581
rect 494367 384547 494379 384581
rect 494379 384547 494401 384581
rect 494439 384547 494447 384581
rect 494447 384547 494473 384581
rect 494511 384547 494515 384581
rect 494515 384547 494545 384581
rect 494583 384547 494617 384581
rect 493359 384089 493393 384123
rect 493431 384089 493461 384123
rect 493461 384089 493465 384123
rect 493503 384089 493529 384123
rect 493529 384089 493537 384123
rect 493575 384089 493597 384123
rect 493597 384089 493609 384123
rect 493647 384089 493665 384123
rect 493665 384089 493681 384123
rect 493719 384089 493733 384123
rect 493733 384089 493753 384123
rect 493791 384089 493801 384123
rect 493801 384089 493825 384123
rect 493863 384089 493869 384123
rect 493869 384089 493897 384123
rect 493935 384089 493937 384123
rect 493937 384089 493969 384123
rect 494007 384089 494039 384123
rect 494039 384089 494041 384123
rect 494079 384089 494107 384123
rect 494107 384089 494113 384123
rect 494151 384089 494175 384123
rect 494175 384089 494185 384123
rect 494223 384089 494243 384123
rect 494243 384089 494257 384123
rect 494295 384089 494311 384123
rect 494311 384089 494329 384123
rect 494367 384089 494379 384123
rect 494379 384089 494401 384123
rect 494439 384089 494447 384123
rect 494447 384089 494473 384123
rect 494511 384089 494515 384123
rect 494515 384089 494545 384123
rect 494583 384089 494617 384123
rect 493091 383907 493125 383941
rect 493091 383507 493125 383541
rect 493091 383107 493125 383141
rect 493091 382707 493125 382741
rect 493359 383631 493393 383665
rect 493431 383631 493461 383665
rect 493461 383631 493465 383665
rect 493503 383631 493529 383665
rect 493529 383631 493537 383665
rect 493575 383631 493597 383665
rect 493597 383631 493609 383665
rect 493647 383631 493665 383665
rect 493665 383631 493681 383665
rect 493719 383631 493733 383665
rect 493733 383631 493753 383665
rect 493791 383631 493801 383665
rect 493801 383631 493825 383665
rect 493863 383631 493869 383665
rect 493869 383631 493897 383665
rect 493935 383631 493937 383665
rect 493937 383631 493969 383665
rect 494007 383631 494039 383665
rect 494039 383631 494041 383665
rect 494079 383631 494107 383665
rect 494107 383631 494113 383665
rect 494151 383631 494175 383665
rect 494175 383631 494185 383665
rect 494223 383631 494243 383665
rect 494243 383631 494257 383665
rect 494295 383631 494311 383665
rect 494311 383631 494329 383665
rect 494367 383631 494379 383665
rect 494379 383631 494401 383665
rect 494439 383631 494447 383665
rect 494447 383631 494473 383665
rect 494511 383631 494515 383665
rect 494515 383631 494545 383665
rect 494583 383631 494617 383665
rect 493359 383173 493393 383207
rect 493431 383173 493461 383207
rect 493461 383173 493465 383207
rect 493503 383173 493529 383207
rect 493529 383173 493537 383207
rect 493575 383173 493597 383207
rect 493597 383173 493609 383207
rect 493647 383173 493665 383207
rect 493665 383173 493681 383207
rect 493719 383173 493733 383207
rect 493733 383173 493753 383207
rect 493791 383173 493801 383207
rect 493801 383173 493825 383207
rect 493863 383173 493869 383207
rect 493869 383173 493897 383207
rect 493935 383173 493937 383207
rect 493937 383173 493969 383207
rect 494007 383173 494039 383207
rect 494039 383173 494041 383207
rect 494079 383173 494107 383207
rect 494107 383173 494113 383207
rect 494151 383173 494175 383207
rect 494175 383173 494185 383207
rect 494223 383173 494243 383207
rect 494243 383173 494257 383207
rect 494295 383173 494311 383207
rect 494311 383173 494329 383207
rect 494367 383173 494379 383207
rect 494379 383173 494401 383207
rect 494439 383173 494447 383207
rect 494447 383173 494473 383207
rect 494511 383173 494515 383207
rect 494515 383173 494545 383207
rect 494583 383173 494617 383207
rect 493091 382307 493125 382341
rect 493091 381907 493125 381941
rect 493091 381507 493125 381541
rect 493359 382715 493393 382749
rect 493431 382715 493461 382749
rect 493461 382715 493465 382749
rect 493503 382715 493529 382749
rect 493529 382715 493537 382749
rect 493575 382715 493597 382749
rect 493597 382715 493609 382749
rect 493647 382715 493665 382749
rect 493665 382715 493681 382749
rect 493719 382715 493733 382749
rect 493733 382715 493753 382749
rect 493791 382715 493801 382749
rect 493801 382715 493825 382749
rect 493863 382715 493869 382749
rect 493869 382715 493897 382749
rect 493935 382715 493937 382749
rect 493937 382715 493969 382749
rect 494007 382715 494039 382749
rect 494039 382715 494041 382749
rect 494079 382715 494107 382749
rect 494107 382715 494113 382749
rect 494151 382715 494175 382749
rect 494175 382715 494185 382749
rect 494223 382715 494243 382749
rect 494243 382715 494257 382749
rect 494295 382715 494311 382749
rect 494311 382715 494329 382749
rect 494367 382715 494379 382749
rect 494379 382715 494401 382749
rect 494439 382715 494447 382749
rect 494447 382715 494473 382749
rect 494511 382715 494515 382749
rect 494515 382715 494545 382749
rect 494583 382715 494617 382749
rect 493359 382257 493393 382291
rect 493431 382257 493461 382291
rect 493461 382257 493465 382291
rect 493503 382257 493529 382291
rect 493529 382257 493537 382291
rect 493575 382257 493597 382291
rect 493597 382257 493609 382291
rect 493647 382257 493665 382291
rect 493665 382257 493681 382291
rect 493719 382257 493733 382291
rect 493733 382257 493753 382291
rect 493791 382257 493801 382291
rect 493801 382257 493825 382291
rect 493863 382257 493869 382291
rect 493869 382257 493897 382291
rect 493935 382257 493937 382291
rect 493937 382257 493969 382291
rect 494007 382257 494039 382291
rect 494039 382257 494041 382291
rect 494079 382257 494107 382291
rect 494107 382257 494113 382291
rect 494151 382257 494175 382291
rect 494175 382257 494185 382291
rect 494223 382257 494243 382291
rect 494243 382257 494257 382291
rect 494295 382257 494311 382291
rect 494311 382257 494329 382291
rect 494367 382257 494379 382291
rect 494379 382257 494401 382291
rect 494439 382257 494447 382291
rect 494447 382257 494473 382291
rect 494511 382257 494515 382291
rect 494515 382257 494545 382291
rect 494583 382257 494617 382291
rect 493359 381799 493393 381833
rect 493431 381799 493461 381833
rect 493461 381799 493465 381833
rect 493503 381799 493529 381833
rect 493529 381799 493537 381833
rect 493575 381799 493597 381833
rect 493597 381799 493609 381833
rect 493647 381799 493665 381833
rect 493665 381799 493681 381833
rect 493719 381799 493733 381833
rect 493733 381799 493753 381833
rect 493791 381799 493801 381833
rect 493801 381799 493825 381833
rect 493863 381799 493869 381833
rect 493869 381799 493897 381833
rect 493935 381799 493937 381833
rect 493937 381799 493969 381833
rect 494007 381799 494039 381833
rect 494039 381799 494041 381833
rect 494079 381799 494107 381833
rect 494107 381799 494113 381833
rect 494151 381799 494175 381833
rect 494175 381799 494185 381833
rect 494223 381799 494243 381833
rect 494243 381799 494257 381833
rect 494295 381799 494311 381833
rect 494311 381799 494329 381833
rect 494367 381799 494379 381833
rect 494379 381799 494401 381833
rect 494439 381799 494447 381833
rect 494447 381799 494473 381833
rect 494511 381799 494515 381833
rect 494515 381799 494545 381833
rect 494583 381799 494617 381833
rect 493359 381341 493393 381375
rect 493431 381341 493461 381375
rect 493461 381341 493465 381375
rect 493503 381341 493529 381375
rect 493529 381341 493537 381375
rect 493575 381341 493597 381375
rect 493597 381341 493609 381375
rect 493647 381341 493665 381375
rect 493665 381341 493681 381375
rect 493719 381341 493733 381375
rect 493733 381341 493753 381375
rect 493791 381341 493801 381375
rect 493801 381341 493825 381375
rect 493863 381341 493869 381375
rect 493869 381341 493897 381375
rect 493935 381341 493937 381375
rect 493937 381341 493969 381375
rect 494007 381341 494039 381375
rect 494039 381341 494041 381375
rect 494079 381341 494107 381375
rect 494107 381341 494113 381375
rect 494151 381341 494175 381375
rect 494175 381341 494185 381375
rect 494223 381341 494243 381375
rect 494243 381341 494257 381375
rect 494295 381341 494311 381375
rect 494311 381341 494329 381375
rect 494367 381341 494379 381375
rect 494379 381341 494401 381375
rect 494439 381341 494447 381375
rect 494447 381341 494473 381375
rect 494511 381341 494515 381375
rect 494515 381341 494545 381375
rect 494583 381341 494617 381375
rect 493091 381107 493125 381141
rect 493091 380707 493125 380741
rect 493091 380307 493125 380341
rect 493359 380883 493393 380917
rect 493431 380883 493461 380917
rect 493461 380883 493465 380917
rect 493503 380883 493529 380917
rect 493529 380883 493537 380917
rect 493575 380883 493597 380917
rect 493597 380883 493609 380917
rect 493647 380883 493665 380917
rect 493665 380883 493681 380917
rect 493719 380883 493733 380917
rect 493733 380883 493753 380917
rect 493791 380883 493801 380917
rect 493801 380883 493825 380917
rect 493863 380883 493869 380917
rect 493869 380883 493897 380917
rect 493935 380883 493937 380917
rect 493937 380883 493969 380917
rect 494007 380883 494039 380917
rect 494039 380883 494041 380917
rect 494079 380883 494107 380917
rect 494107 380883 494113 380917
rect 494151 380883 494175 380917
rect 494175 380883 494185 380917
rect 494223 380883 494243 380917
rect 494243 380883 494257 380917
rect 494295 380883 494311 380917
rect 494311 380883 494329 380917
rect 494367 380883 494379 380917
rect 494379 380883 494401 380917
rect 494439 380883 494447 380917
rect 494447 380883 494473 380917
rect 494511 380883 494515 380917
rect 494515 380883 494545 380917
rect 494583 380883 494617 380917
rect 493359 380425 493393 380459
rect 493431 380425 493461 380459
rect 493461 380425 493465 380459
rect 493503 380425 493529 380459
rect 493529 380425 493537 380459
rect 493575 380425 493597 380459
rect 493597 380425 493609 380459
rect 493647 380425 493665 380459
rect 493665 380425 493681 380459
rect 493719 380425 493733 380459
rect 493733 380425 493753 380459
rect 493791 380425 493801 380459
rect 493801 380425 493825 380459
rect 493863 380425 493869 380459
rect 493869 380425 493897 380459
rect 493935 380425 493937 380459
rect 493937 380425 493969 380459
rect 494007 380425 494039 380459
rect 494039 380425 494041 380459
rect 494079 380425 494107 380459
rect 494107 380425 494113 380459
rect 494151 380425 494175 380459
rect 494175 380425 494185 380459
rect 494223 380425 494243 380459
rect 494243 380425 494257 380459
rect 494295 380425 494311 380459
rect 494311 380425 494329 380459
rect 494367 380425 494379 380459
rect 494379 380425 494401 380459
rect 494439 380425 494447 380459
rect 494447 380425 494473 380459
rect 494511 380425 494515 380459
rect 494515 380425 494545 380459
rect 494583 380425 494617 380459
rect 493091 379907 493125 379941
rect 493091 379507 493125 379541
rect 493091 379107 493125 379141
rect 493359 379967 493393 380001
rect 493431 379967 493461 380001
rect 493461 379967 493465 380001
rect 493503 379967 493529 380001
rect 493529 379967 493537 380001
rect 493575 379967 493597 380001
rect 493597 379967 493609 380001
rect 493647 379967 493665 380001
rect 493665 379967 493681 380001
rect 493719 379967 493733 380001
rect 493733 379967 493753 380001
rect 493791 379967 493801 380001
rect 493801 379967 493825 380001
rect 493863 379967 493869 380001
rect 493869 379967 493897 380001
rect 493935 379967 493937 380001
rect 493937 379967 493969 380001
rect 494007 379967 494039 380001
rect 494039 379967 494041 380001
rect 494079 379967 494107 380001
rect 494107 379967 494113 380001
rect 494151 379967 494175 380001
rect 494175 379967 494185 380001
rect 494223 379967 494243 380001
rect 494243 379967 494257 380001
rect 494295 379967 494311 380001
rect 494311 379967 494329 380001
rect 494367 379967 494379 380001
rect 494379 379967 494401 380001
rect 494439 379967 494447 380001
rect 494447 379967 494473 380001
rect 494511 379967 494515 380001
rect 494515 379967 494545 380001
rect 494583 379967 494617 380001
rect 493359 379509 493393 379543
rect 493431 379509 493461 379543
rect 493461 379509 493465 379543
rect 493503 379509 493529 379543
rect 493529 379509 493537 379543
rect 493575 379509 493597 379543
rect 493597 379509 493609 379543
rect 493647 379509 493665 379543
rect 493665 379509 493681 379543
rect 493719 379509 493733 379543
rect 493733 379509 493753 379543
rect 493791 379509 493801 379543
rect 493801 379509 493825 379543
rect 493863 379509 493869 379543
rect 493869 379509 493897 379543
rect 493935 379509 493937 379543
rect 493937 379509 493969 379543
rect 494007 379509 494039 379543
rect 494039 379509 494041 379543
rect 494079 379509 494107 379543
rect 494107 379509 494113 379543
rect 494151 379509 494175 379543
rect 494175 379509 494185 379543
rect 494223 379509 494243 379543
rect 494243 379509 494257 379543
rect 494295 379509 494311 379543
rect 494311 379509 494329 379543
rect 494367 379509 494379 379543
rect 494379 379509 494401 379543
rect 494439 379509 494447 379543
rect 494447 379509 494473 379543
rect 494511 379509 494515 379543
rect 494515 379509 494545 379543
rect 494583 379509 494617 379543
rect 493091 378707 493125 378741
rect 493359 379051 493393 379085
rect 493431 379051 493461 379085
rect 493461 379051 493465 379085
rect 493503 379051 493529 379085
rect 493529 379051 493537 379085
rect 493575 379051 493597 379085
rect 493597 379051 493609 379085
rect 493647 379051 493665 379085
rect 493665 379051 493681 379085
rect 493719 379051 493733 379085
rect 493733 379051 493753 379085
rect 493791 379051 493801 379085
rect 493801 379051 493825 379085
rect 493863 379051 493869 379085
rect 493869 379051 493897 379085
rect 493935 379051 493937 379085
rect 493937 379051 493969 379085
rect 494007 379051 494039 379085
rect 494039 379051 494041 379085
rect 494079 379051 494107 379085
rect 494107 379051 494113 379085
rect 494151 379051 494175 379085
rect 494175 379051 494185 379085
rect 494223 379051 494243 379085
rect 494243 379051 494257 379085
rect 494295 379051 494311 379085
rect 494311 379051 494329 379085
rect 494367 379051 494379 379085
rect 494379 379051 494401 379085
rect 494439 379051 494447 379085
rect 494447 379051 494473 379085
rect 494511 379051 494515 379085
rect 494515 379051 494545 379085
rect 494583 379051 494617 379085
rect 493359 378593 493393 378627
rect 493431 378593 493461 378627
rect 493461 378593 493465 378627
rect 493503 378593 493529 378627
rect 493529 378593 493537 378627
rect 493575 378593 493597 378627
rect 493597 378593 493609 378627
rect 493647 378593 493665 378627
rect 493665 378593 493681 378627
rect 493719 378593 493733 378627
rect 493733 378593 493753 378627
rect 493791 378593 493801 378627
rect 493801 378593 493825 378627
rect 493863 378593 493869 378627
rect 493869 378593 493897 378627
rect 493935 378593 493937 378627
rect 493937 378593 493969 378627
rect 494007 378593 494039 378627
rect 494039 378593 494041 378627
rect 494079 378593 494107 378627
rect 494107 378593 494113 378627
rect 494151 378593 494175 378627
rect 494175 378593 494185 378627
rect 494223 378593 494243 378627
rect 494243 378593 494257 378627
rect 494295 378593 494311 378627
rect 494311 378593 494329 378627
rect 494367 378593 494379 378627
rect 494379 378593 494401 378627
rect 494439 378593 494447 378627
rect 494447 378593 494473 378627
rect 494511 378593 494515 378627
rect 494515 378593 494545 378627
rect 494583 378593 494617 378627
rect 493091 378307 493125 378341
rect 493091 377907 493125 377941
rect 493091 377507 493125 377541
rect 493359 378135 493393 378169
rect 493431 378135 493461 378169
rect 493461 378135 493465 378169
rect 493503 378135 493529 378169
rect 493529 378135 493537 378169
rect 493575 378135 493597 378169
rect 493597 378135 493609 378169
rect 493647 378135 493665 378169
rect 493665 378135 493681 378169
rect 493719 378135 493733 378169
rect 493733 378135 493753 378169
rect 493791 378135 493801 378169
rect 493801 378135 493825 378169
rect 493863 378135 493869 378169
rect 493869 378135 493897 378169
rect 493935 378135 493937 378169
rect 493937 378135 493969 378169
rect 494007 378135 494039 378169
rect 494039 378135 494041 378169
rect 494079 378135 494107 378169
rect 494107 378135 494113 378169
rect 494151 378135 494175 378169
rect 494175 378135 494185 378169
rect 494223 378135 494243 378169
rect 494243 378135 494257 378169
rect 494295 378135 494311 378169
rect 494311 378135 494329 378169
rect 494367 378135 494379 378169
rect 494379 378135 494401 378169
rect 494439 378135 494447 378169
rect 494447 378135 494473 378169
rect 494511 378135 494515 378169
rect 494515 378135 494545 378169
rect 494583 378135 494617 378169
rect 493359 377677 493393 377711
rect 493431 377677 493461 377711
rect 493461 377677 493465 377711
rect 493503 377677 493529 377711
rect 493529 377677 493537 377711
rect 493575 377677 493597 377711
rect 493597 377677 493609 377711
rect 493647 377677 493665 377711
rect 493665 377677 493681 377711
rect 493719 377677 493733 377711
rect 493733 377677 493753 377711
rect 493791 377677 493801 377711
rect 493801 377677 493825 377711
rect 493863 377677 493869 377711
rect 493869 377677 493897 377711
rect 493935 377677 493937 377711
rect 493937 377677 493969 377711
rect 494007 377677 494039 377711
rect 494039 377677 494041 377711
rect 494079 377677 494107 377711
rect 494107 377677 494113 377711
rect 494151 377677 494175 377711
rect 494175 377677 494185 377711
rect 494223 377677 494243 377711
rect 494243 377677 494257 377711
rect 494295 377677 494311 377711
rect 494311 377677 494329 377711
rect 494367 377677 494379 377711
rect 494379 377677 494401 377711
rect 494439 377677 494447 377711
rect 494447 377677 494473 377711
rect 494511 377677 494515 377711
rect 494515 377677 494545 377711
rect 494583 377677 494617 377711
rect 493091 377107 493125 377141
rect 493091 376707 493125 376741
rect 493091 376307 493125 376341
rect 493359 377219 493393 377253
rect 493431 377219 493461 377253
rect 493461 377219 493465 377253
rect 493503 377219 493529 377253
rect 493529 377219 493537 377253
rect 493575 377219 493597 377253
rect 493597 377219 493609 377253
rect 493647 377219 493665 377253
rect 493665 377219 493681 377253
rect 493719 377219 493733 377253
rect 493733 377219 493753 377253
rect 493791 377219 493801 377253
rect 493801 377219 493825 377253
rect 493863 377219 493869 377253
rect 493869 377219 493897 377253
rect 493935 377219 493937 377253
rect 493937 377219 493969 377253
rect 494007 377219 494039 377253
rect 494039 377219 494041 377253
rect 494079 377219 494107 377253
rect 494107 377219 494113 377253
rect 494151 377219 494175 377253
rect 494175 377219 494185 377253
rect 494223 377219 494243 377253
rect 494243 377219 494257 377253
rect 494295 377219 494311 377253
rect 494311 377219 494329 377253
rect 494367 377219 494379 377253
rect 494379 377219 494401 377253
rect 494439 377219 494447 377253
rect 494447 377219 494473 377253
rect 494511 377219 494515 377253
rect 494515 377219 494545 377253
rect 494583 377219 494617 377253
rect 493359 376761 493393 376795
rect 493431 376761 493461 376795
rect 493461 376761 493465 376795
rect 493503 376761 493529 376795
rect 493529 376761 493537 376795
rect 493575 376761 493597 376795
rect 493597 376761 493609 376795
rect 493647 376761 493665 376795
rect 493665 376761 493681 376795
rect 493719 376761 493733 376795
rect 493733 376761 493753 376795
rect 493791 376761 493801 376795
rect 493801 376761 493825 376795
rect 493863 376761 493869 376795
rect 493869 376761 493897 376795
rect 493935 376761 493937 376795
rect 493937 376761 493969 376795
rect 494007 376761 494039 376795
rect 494039 376761 494041 376795
rect 494079 376761 494107 376795
rect 494107 376761 494113 376795
rect 494151 376761 494175 376795
rect 494175 376761 494185 376795
rect 494223 376761 494243 376795
rect 494243 376761 494257 376795
rect 494295 376761 494311 376795
rect 494311 376761 494329 376795
rect 494367 376761 494379 376795
rect 494379 376761 494401 376795
rect 494439 376761 494447 376795
rect 494447 376761 494473 376795
rect 494511 376761 494515 376795
rect 494515 376761 494545 376795
rect 494583 376761 494617 376795
rect 493091 375907 493125 375941
rect 493091 375507 493125 375541
rect 493091 375107 493125 375141
rect 493359 376303 493393 376337
rect 493431 376303 493461 376337
rect 493461 376303 493465 376337
rect 493503 376303 493529 376337
rect 493529 376303 493537 376337
rect 493575 376303 493597 376337
rect 493597 376303 493609 376337
rect 493647 376303 493665 376337
rect 493665 376303 493681 376337
rect 493719 376303 493733 376337
rect 493733 376303 493753 376337
rect 493791 376303 493801 376337
rect 493801 376303 493825 376337
rect 493863 376303 493869 376337
rect 493869 376303 493897 376337
rect 493935 376303 493937 376337
rect 493937 376303 493969 376337
rect 494007 376303 494039 376337
rect 494039 376303 494041 376337
rect 494079 376303 494107 376337
rect 494107 376303 494113 376337
rect 494151 376303 494175 376337
rect 494175 376303 494185 376337
rect 494223 376303 494243 376337
rect 494243 376303 494257 376337
rect 494295 376303 494311 376337
rect 494311 376303 494329 376337
rect 494367 376303 494379 376337
rect 494379 376303 494401 376337
rect 494439 376303 494447 376337
rect 494447 376303 494473 376337
rect 494511 376303 494515 376337
rect 494515 376303 494545 376337
rect 494583 376303 494617 376337
rect 493359 375845 493393 375879
rect 493431 375845 493461 375879
rect 493461 375845 493465 375879
rect 493503 375845 493529 375879
rect 493529 375845 493537 375879
rect 493575 375845 493597 375879
rect 493597 375845 493609 375879
rect 493647 375845 493665 375879
rect 493665 375845 493681 375879
rect 493719 375845 493733 375879
rect 493733 375845 493753 375879
rect 493791 375845 493801 375879
rect 493801 375845 493825 375879
rect 493863 375845 493869 375879
rect 493869 375845 493897 375879
rect 493935 375845 493937 375879
rect 493937 375845 493969 375879
rect 494007 375845 494039 375879
rect 494039 375845 494041 375879
rect 494079 375845 494107 375879
rect 494107 375845 494113 375879
rect 494151 375845 494175 375879
rect 494175 375845 494185 375879
rect 494223 375845 494243 375879
rect 494243 375845 494257 375879
rect 494295 375845 494311 375879
rect 494311 375845 494329 375879
rect 494367 375845 494379 375879
rect 494379 375845 494401 375879
rect 494439 375845 494447 375879
rect 494447 375845 494473 375879
rect 494511 375845 494515 375879
rect 494515 375845 494545 375879
rect 494583 375845 494617 375879
rect 493359 375387 493393 375421
rect 493431 375387 493461 375421
rect 493461 375387 493465 375421
rect 493503 375387 493529 375421
rect 493529 375387 493537 375421
rect 493575 375387 493597 375421
rect 493597 375387 493609 375421
rect 493647 375387 493665 375421
rect 493665 375387 493681 375421
rect 493719 375387 493733 375421
rect 493733 375387 493753 375421
rect 493791 375387 493801 375421
rect 493801 375387 493825 375421
rect 493863 375387 493869 375421
rect 493869 375387 493897 375421
rect 493935 375387 493937 375421
rect 493937 375387 493969 375421
rect 494007 375387 494039 375421
rect 494039 375387 494041 375421
rect 494079 375387 494107 375421
rect 494107 375387 494113 375421
rect 494151 375387 494175 375421
rect 494175 375387 494185 375421
rect 494223 375387 494243 375421
rect 494243 375387 494257 375421
rect 494295 375387 494311 375421
rect 494311 375387 494329 375421
rect 494367 375387 494379 375421
rect 494379 375387 494401 375421
rect 494439 375387 494447 375421
rect 494447 375387 494473 375421
rect 494511 375387 494515 375421
rect 494515 375387 494545 375421
rect 494583 375387 494617 375421
rect 493359 374929 493393 374963
rect 493431 374929 493461 374963
rect 493461 374929 493465 374963
rect 493503 374929 493529 374963
rect 493529 374929 493537 374963
rect 493575 374929 493597 374963
rect 493597 374929 493609 374963
rect 493647 374929 493665 374963
rect 493665 374929 493681 374963
rect 493719 374929 493733 374963
rect 493733 374929 493753 374963
rect 493791 374929 493801 374963
rect 493801 374929 493825 374963
rect 493863 374929 493869 374963
rect 493869 374929 493897 374963
rect 493935 374929 493937 374963
rect 493937 374929 493969 374963
rect 494007 374929 494039 374963
rect 494039 374929 494041 374963
rect 494079 374929 494107 374963
rect 494107 374929 494113 374963
rect 494151 374929 494175 374963
rect 494175 374929 494185 374963
rect 494223 374929 494243 374963
rect 494243 374929 494257 374963
rect 494295 374929 494311 374963
rect 494311 374929 494329 374963
rect 494367 374929 494379 374963
rect 494379 374929 494401 374963
rect 494439 374929 494447 374963
rect 494447 374929 494473 374963
rect 494511 374929 494515 374963
rect 494515 374929 494545 374963
rect 494583 374929 494617 374963
rect 493091 374707 493125 374741
rect 493091 374307 493125 374341
rect 493091 373907 493125 373941
rect 493359 374471 493393 374505
rect 493431 374471 493461 374505
rect 493461 374471 493465 374505
rect 493503 374471 493529 374505
rect 493529 374471 493537 374505
rect 493575 374471 493597 374505
rect 493597 374471 493609 374505
rect 493647 374471 493665 374505
rect 493665 374471 493681 374505
rect 493719 374471 493733 374505
rect 493733 374471 493753 374505
rect 493791 374471 493801 374505
rect 493801 374471 493825 374505
rect 493863 374471 493869 374505
rect 493869 374471 493897 374505
rect 493935 374471 493937 374505
rect 493937 374471 493969 374505
rect 494007 374471 494039 374505
rect 494039 374471 494041 374505
rect 494079 374471 494107 374505
rect 494107 374471 494113 374505
rect 494151 374471 494175 374505
rect 494175 374471 494185 374505
rect 494223 374471 494243 374505
rect 494243 374471 494257 374505
rect 494295 374471 494311 374505
rect 494311 374471 494329 374505
rect 494367 374471 494379 374505
rect 494379 374471 494401 374505
rect 494439 374471 494447 374505
rect 494447 374471 494473 374505
rect 494511 374471 494515 374505
rect 494515 374471 494545 374505
rect 494583 374471 494617 374505
rect 493359 374013 493393 374047
rect 493431 374013 493461 374047
rect 493461 374013 493465 374047
rect 493503 374013 493529 374047
rect 493529 374013 493537 374047
rect 493575 374013 493597 374047
rect 493597 374013 493609 374047
rect 493647 374013 493665 374047
rect 493665 374013 493681 374047
rect 493719 374013 493733 374047
rect 493733 374013 493753 374047
rect 493791 374013 493801 374047
rect 493801 374013 493825 374047
rect 493863 374013 493869 374047
rect 493869 374013 493897 374047
rect 493935 374013 493937 374047
rect 493937 374013 493969 374047
rect 494007 374013 494039 374047
rect 494039 374013 494041 374047
rect 494079 374013 494107 374047
rect 494107 374013 494113 374047
rect 494151 374013 494175 374047
rect 494175 374013 494185 374047
rect 494223 374013 494243 374047
rect 494243 374013 494257 374047
rect 494295 374013 494311 374047
rect 494311 374013 494329 374047
rect 494367 374013 494379 374047
rect 494379 374013 494401 374047
rect 494439 374013 494447 374047
rect 494447 374013 494473 374047
rect 494511 374013 494515 374047
rect 494515 374013 494545 374047
rect 494583 374013 494617 374047
rect 493091 373507 493125 373541
rect 493091 373107 493125 373141
rect 493091 372707 493125 372741
rect 493091 372307 493125 372341
rect 493359 373555 493393 373589
rect 493431 373555 493461 373589
rect 493461 373555 493465 373589
rect 493503 373555 493529 373589
rect 493529 373555 493537 373589
rect 493575 373555 493597 373589
rect 493597 373555 493609 373589
rect 493647 373555 493665 373589
rect 493665 373555 493681 373589
rect 493719 373555 493733 373589
rect 493733 373555 493753 373589
rect 493791 373555 493801 373589
rect 493801 373555 493825 373589
rect 493863 373555 493869 373589
rect 493869 373555 493897 373589
rect 493935 373555 493937 373589
rect 493937 373555 493969 373589
rect 494007 373555 494039 373589
rect 494039 373555 494041 373589
rect 494079 373555 494107 373589
rect 494107 373555 494113 373589
rect 494151 373555 494175 373589
rect 494175 373555 494185 373589
rect 494223 373555 494243 373589
rect 494243 373555 494257 373589
rect 494295 373555 494311 373589
rect 494311 373555 494329 373589
rect 494367 373555 494379 373589
rect 494379 373555 494401 373589
rect 494439 373555 494447 373589
rect 494447 373555 494473 373589
rect 494511 373555 494515 373589
rect 494515 373555 494545 373589
rect 494583 373555 494617 373589
rect 493359 373097 493393 373131
rect 493431 373097 493461 373131
rect 493461 373097 493465 373131
rect 493503 373097 493529 373131
rect 493529 373097 493537 373131
rect 493575 373097 493597 373131
rect 493597 373097 493609 373131
rect 493647 373097 493665 373131
rect 493665 373097 493681 373131
rect 493719 373097 493733 373131
rect 493733 373097 493753 373131
rect 493791 373097 493801 373131
rect 493801 373097 493825 373131
rect 493863 373097 493869 373131
rect 493869 373097 493897 373131
rect 493935 373097 493937 373131
rect 493937 373097 493969 373131
rect 494007 373097 494039 373131
rect 494039 373097 494041 373131
rect 494079 373097 494107 373131
rect 494107 373097 494113 373131
rect 494151 373097 494175 373131
rect 494175 373097 494185 373131
rect 494223 373097 494243 373131
rect 494243 373097 494257 373131
rect 494295 373097 494311 373131
rect 494311 373097 494329 373131
rect 494367 373097 494379 373131
rect 494379 373097 494401 373131
rect 494439 373097 494447 373131
rect 494447 373097 494473 373131
rect 494511 373097 494515 373131
rect 494515 373097 494545 373131
rect 494583 373097 494617 373131
rect 493359 372639 493393 372673
rect 493431 372639 493461 372673
rect 493461 372639 493465 372673
rect 493503 372639 493529 372673
rect 493529 372639 493537 372673
rect 493575 372639 493597 372673
rect 493597 372639 493609 372673
rect 493647 372639 493665 372673
rect 493665 372639 493681 372673
rect 493719 372639 493733 372673
rect 493733 372639 493753 372673
rect 493791 372639 493801 372673
rect 493801 372639 493825 372673
rect 493863 372639 493869 372673
rect 493869 372639 493897 372673
rect 493935 372639 493937 372673
rect 493937 372639 493969 372673
rect 494007 372639 494039 372673
rect 494039 372639 494041 372673
rect 494079 372639 494107 372673
rect 494107 372639 494113 372673
rect 494151 372639 494175 372673
rect 494175 372639 494185 372673
rect 494223 372639 494243 372673
rect 494243 372639 494257 372673
rect 494295 372639 494311 372673
rect 494311 372639 494329 372673
rect 494367 372639 494379 372673
rect 494379 372639 494401 372673
rect 494439 372639 494447 372673
rect 494447 372639 494473 372673
rect 494511 372639 494515 372673
rect 494515 372639 494545 372673
rect 494583 372639 494617 372673
rect 493359 372181 493393 372215
rect 493431 372181 493461 372215
rect 493461 372181 493465 372215
rect 493503 372181 493529 372215
rect 493529 372181 493537 372215
rect 493575 372181 493597 372215
rect 493597 372181 493609 372215
rect 493647 372181 493665 372215
rect 493665 372181 493681 372215
rect 493719 372181 493733 372215
rect 493733 372181 493753 372215
rect 493791 372181 493801 372215
rect 493801 372181 493825 372215
rect 493863 372181 493869 372215
rect 493869 372181 493897 372215
rect 493935 372181 493937 372215
rect 493937 372181 493969 372215
rect 494007 372181 494039 372215
rect 494039 372181 494041 372215
rect 494079 372181 494107 372215
rect 494107 372181 494113 372215
rect 494151 372181 494175 372215
rect 494175 372181 494185 372215
rect 494223 372181 494243 372215
rect 494243 372181 494257 372215
rect 494295 372181 494311 372215
rect 494311 372181 494329 372215
rect 494367 372181 494379 372215
rect 494379 372181 494401 372215
rect 494439 372181 494447 372215
rect 494447 372181 494473 372215
rect 494511 372181 494515 372215
rect 494515 372181 494545 372215
rect 494583 372181 494617 372215
rect 493091 371907 493125 371941
rect 493091 371507 493125 371541
rect 493091 371107 493125 371141
rect 493359 371723 493393 371757
rect 493431 371723 493461 371757
rect 493461 371723 493465 371757
rect 493503 371723 493529 371757
rect 493529 371723 493537 371757
rect 493575 371723 493597 371757
rect 493597 371723 493609 371757
rect 493647 371723 493665 371757
rect 493665 371723 493681 371757
rect 493719 371723 493733 371757
rect 493733 371723 493753 371757
rect 493791 371723 493801 371757
rect 493801 371723 493825 371757
rect 493863 371723 493869 371757
rect 493869 371723 493897 371757
rect 493935 371723 493937 371757
rect 493937 371723 493969 371757
rect 494007 371723 494039 371757
rect 494039 371723 494041 371757
rect 494079 371723 494107 371757
rect 494107 371723 494113 371757
rect 494151 371723 494175 371757
rect 494175 371723 494185 371757
rect 494223 371723 494243 371757
rect 494243 371723 494257 371757
rect 494295 371723 494311 371757
rect 494311 371723 494329 371757
rect 494367 371723 494379 371757
rect 494379 371723 494401 371757
rect 494439 371723 494447 371757
rect 494447 371723 494473 371757
rect 494511 371723 494515 371757
rect 494515 371723 494545 371757
rect 494583 371723 494617 371757
rect 493359 371265 493393 371299
rect 493431 371265 493461 371299
rect 493461 371265 493465 371299
rect 493503 371265 493529 371299
rect 493529 371265 493537 371299
rect 493575 371265 493597 371299
rect 493597 371265 493609 371299
rect 493647 371265 493665 371299
rect 493665 371265 493681 371299
rect 493719 371265 493733 371299
rect 493733 371265 493753 371299
rect 493791 371265 493801 371299
rect 493801 371265 493825 371299
rect 493863 371265 493869 371299
rect 493869 371265 493897 371299
rect 493935 371265 493937 371299
rect 493937 371265 493969 371299
rect 494007 371265 494039 371299
rect 494039 371265 494041 371299
rect 494079 371265 494107 371299
rect 494107 371265 494113 371299
rect 494151 371265 494175 371299
rect 494175 371265 494185 371299
rect 494223 371265 494243 371299
rect 494243 371265 494257 371299
rect 494295 371265 494311 371299
rect 494311 371265 494329 371299
rect 494367 371265 494379 371299
rect 494379 371265 494401 371299
rect 494439 371265 494447 371299
rect 494447 371265 494473 371299
rect 494511 371265 494515 371299
rect 494515 371265 494545 371299
rect 494583 371265 494617 371299
rect 493091 370707 493125 370741
rect 493091 370307 493125 370341
rect 493091 369907 493125 369941
rect 493359 370807 493393 370841
rect 493431 370807 493461 370841
rect 493461 370807 493465 370841
rect 493503 370807 493529 370841
rect 493529 370807 493537 370841
rect 493575 370807 493597 370841
rect 493597 370807 493609 370841
rect 493647 370807 493665 370841
rect 493665 370807 493681 370841
rect 493719 370807 493733 370841
rect 493733 370807 493753 370841
rect 493791 370807 493801 370841
rect 493801 370807 493825 370841
rect 493863 370807 493869 370841
rect 493869 370807 493897 370841
rect 493935 370807 493937 370841
rect 493937 370807 493969 370841
rect 494007 370807 494039 370841
rect 494039 370807 494041 370841
rect 494079 370807 494107 370841
rect 494107 370807 494113 370841
rect 494151 370807 494175 370841
rect 494175 370807 494185 370841
rect 494223 370807 494243 370841
rect 494243 370807 494257 370841
rect 494295 370807 494311 370841
rect 494311 370807 494329 370841
rect 494367 370807 494379 370841
rect 494379 370807 494401 370841
rect 494439 370807 494447 370841
rect 494447 370807 494473 370841
rect 494511 370807 494515 370841
rect 494515 370807 494545 370841
rect 494583 370807 494617 370841
rect 493359 370349 493393 370383
rect 493431 370349 493461 370383
rect 493461 370349 493465 370383
rect 493503 370349 493529 370383
rect 493529 370349 493537 370383
rect 493575 370349 493597 370383
rect 493597 370349 493609 370383
rect 493647 370349 493665 370383
rect 493665 370349 493681 370383
rect 493719 370349 493733 370383
rect 493733 370349 493753 370383
rect 493791 370349 493801 370383
rect 493801 370349 493825 370383
rect 493863 370349 493869 370383
rect 493869 370349 493897 370383
rect 493935 370349 493937 370383
rect 493937 370349 493969 370383
rect 494007 370349 494039 370383
rect 494039 370349 494041 370383
rect 494079 370349 494107 370383
rect 494107 370349 494113 370383
rect 494151 370349 494175 370383
rect 494175 370349 494185 370383
rect 494223 370349 494243 370383
rect 494243 370349 494257 370383
rect 494295 370349 494311 370383
rect 494311 370349 494329 370383
rect 494367 370349 494379 370383
rect 494379 370349 494401 370383
rect 494439 370349 494447 370383
rect 494447 370349 494473 370383
rect 494511 370349 494515 370383
rect 494515 370349 494545 370383
rect 494583 370349 494617 370383
rect 493091 369507 493125 369541
rect 493091 369107 493125 369141
rect 493091 368707 493125 368741
rect 493359 369891 493393 369925
rect 493431 369891 493461 369925
rect 493461 369891 493465 369925
rect 493503 369891 493529 369925
rect 493529 369891 493537 369925
rect 493575 369891 493597 369925
rect 493597 369891 493609 369925
rect 493647 369891 493665 369925
rect 493665 369891 493681 369925
rect 493719 369891 493733 369925
rect 493733 369891 493753 369925
rect 493791 369891 493801 369925
rect 493801 369891 493825 369925
rect 493863 369891 493869 369925
rect 493869 369891 493897 369925
rect 493935 369891 493937 369925
rect 493937 369891 493969 369925
rect 494007 369891 494039 369925
rect 494039 369891 494041 369925
rect 494079 369891 494107 369925
rect 494107 369891 494113 369925
rect 494151 369891 494175 369925
rect 494175 369891 494185 369925
rect 494223 369891 494243 369925
rect 494243 369891 494257 369925
rect 494295 369891 494311 369925
rect 494311 369891 494329 369925
rect 494367 369891 494379 369925
rect 494379 369891 494401 369925
rect 494439 369891 494447 369925
rect 494447 369891 494473 369925
rect 494511 369891 494515 369925
rect 494515 369891 494545 369925
rect 494583 369891 494617 369925
rect 493359 369433 493393 369467
rect 493431 369433 493461 369467
rect 493461 369433 493465 369467
rect 493503 369433 493529 369467
rect 493529 369433 493537 369467
rect 493575 369433 493597 369467
rect 493597 369433 493609 369467
rect 493647 369433 493665 369467
rect 493665 369433 493681 369467
rect 493719 369433 493733 369467
rect 493733 369433 493753 369467
rect 493791 369433 493801 369467
rect 493801 369433 493825 369467
rect 493863 369433 493869 369467
rect 493869 369433 493897 369467
rect 493935 369433 493937 369467
rect 493937 369433 493969 369467
rect 494007 369433 494039 369467
rect 494039 369433 494041 369467
rect 494079 369433 494107 369467
rect 494107 369433 494113 369467
rect 494151 369433 494175 369467
rect 494175 369433 494185 369467
rect 494223 369433 494243 369467
rect 494243 369433 494257 369467
rect 494295 369433 494311 369467
rect 494311 369433 494329 369467
rect 494367 369433 494379 369467
rect 494379 369433 494401 369467
rect 494439 369433 494447 369467
rect 494447 369433 494473 369467
rect 494511 369433 494515 369467
rect 494515 369433 494545 369467
rect 494583 369433 494617 369467
rect 493359 368975 493393 369009
rect 493431 368975 493461 369009
rect 493461 368975 493465 369009
rect 493503 368975 493529 369009
rect 493529 368975 493537 369009
rect 493575 368975 493597 369009
rect 493597 368975 493609 369009
rect 493647 368975 493665 369009
rect 493665 368975 493681 369009
rect 493719 368975 493733 369009
rect 493733 368975 493753 369009
rect 493791 368975 493801 369009
rect 493801 368975 493825 369009
rect 493863 368975 493869 369009
rect 493869 368975 493897 369009
rect 493935 368975 493937 369009
rect 493937 368975 493969 369009
rect 494007 368975 494039 369009
rect 494039 368975 494041 369009
rect 494079 368975 494107 369009
rect 494107 368975 494113 369009
rect 494151 368975 494175 369009
rect 494175 368975 494185 369009
rect 494223 368975 494243 369009
rect 494243 368975 494257 369009
rect 494295 368975 494311 369009
rect 494311 368975 494329 369009
rect 494367 368975 494379 369009
rect 494379 368975 494401 369009
rect 494439 368975 494447 369009
rect 494447 368975 494473 369009
rect 494511 368975 494515 369009
rect 494515 368975 494545 369009
rect 494583 368975 494617 369009
rect 493359 368517 493393 368551
rect 493431 368517 493461 368551
rect 493461 368517 493465 368551
rect 493503 368517 493529 368551
rect 493529 368517 493537 368551
rect 493575 368517 493597 368551
rect 493597 368517 493609 368551
rect 493647 368517 493665 368551
rect 493665 368517 493681 368551
rect 493719 368517 493733 368551
rect 493733 368517 493753 368551
rect 493791 368517 493801 368551
rect 493801 368517 493825 368551
rect 493863 368517 493869 368551
rect 493869 368517 493897 368551
rect 493935 368517 493937 368551
rect 493937 368517 493969 368551
rect 494007 368517 494039 368551
rect 494039 368517 494041 368551
rect 494079 368517 494107 368551
rect 494107 368517 494113 368551
rect 494151 368517 494175 368551
rect 494175 368517 494185 368551
rect 494223 368517 494243 368551
rect 494243 368517 494257 368551
rect 494295 368517 494311 368551
rect 494311 368517 494329 368551
rect 494367 368517 494379 368551
rect 494379 368517 494401 368551
rect 494439 368517 494447 368551
rect 494447 368517 494473 368551
rect 494511 368517 494515 368551
rect 494515 368517 494545 368551
rect 494583 368517 494617 368551
rect 493091 368307 493125 368341
rect 493091 367907 493125 367941
rect 493091 367507 493125 367541
rect 493091 367107 493125 367141
rect 493359 368059 493393 368093
rect 493431 368059 493461 368093
rect 493461 368059 493465 368093
rect 493503 368059 493529 368093
rect 493529 368059 493537 368093
rect 493575 368059 493597 368093
rect 493597 368059 493609 368093
rect 493647 368059 493665 368093
rect 493665 368059 493681 368093
rect 493719 368059 493733 368093
rect 493733 368059 493753 368093
rect 493791 368059 493801 368093
rect 493801 368059 493825 368093
rect 493863 368059 493869 368093
rect 493869 368059 493897 368093
rect 493935 368059 493937 368093
rect 493937 368059 493969 368093
rect 494007 368059 494039 368093
rect 494039 368059 494041 368093
rect 494079 368059 494107 368093
rect 494107 368059 494113 368093
rect 494151 368059 494175 368093
rect 494175 368059 494185 368093
rect 494223 368059 494243 368093
rect 494243 368059 494257 368093
rect 494295 368059 494311 368093
rect 494311 368059 494329 368093
rect 494367 368059 494379 368093
rect 494379 368059 494401 368093
rect 494439 368059 494447 368093
rect 494447 368059 494473 368093
rect 494511 368059 494515 368093
rect 494515 368059 494545 368093
rect 494583 368059 494617 368093
rect 493359 367601 493393 367635
rect 493431 367601 493461 367635
rect 493461 367601 493465 367635
rect 493503 367601 493529 367635
rect 493529 367601 493537 367635
rect 493575 367601 493597 367635
rect 493597 367601 493609 367635
rect 493647 367601 493665 367635
rect 493665 367601 493681 367635
rect 493719 367601 493733 367635
rect 493733 367601 493753 367635
rect 493791 367601 493801 367635
rect 493801 367601 493825 367635
rect 493863 367601 493869 367635
rect 493869 367601 493897 367635
rect 493935 367601 493937 367635
rect 493937 367601 493969 367635
rect 494007 367601 494039 367635
rect 494039 367601 494041 367635
rect 494079 367601 494107 367635
rect 494107 367601 494113 367635
rect 494151 367601 494175 367635
rect 494175 367601 494185 367635
rect 494223 367601 494243 367635
rect 494243 367601 494257 367635
rect 494295 367601 494311 367635
rect 494311 367601 494329 367635
rect 494367 367601 494379 367635
rect 494379 367601 494401 367635
rect 494439 367601 494447 367635
rect 494447 367601 494473 367635
rect 494511 367601 494515 367635
rect 494515 367601 494545 367635
rect 494583 367601 494617 367635
rect 493091 366707 493125 366741
rect 493091 366307 493125 366341
rect 493091 365907 493125 365941
rect 493359 367143 493393 367177
rect 493431 367143 493461 367177
rect 493461 367143 493465 367177
rect 493503 367143 493529 367177
rect 493529 367143 493537 367177
rect 493575 367143 493597 367177
rect 493597 367143 493609 367177
rect 493647 367143 493665 367177
rect 493665 367143 493681 367177
rect 493719 367143 493733 367177
rect 493733 367143 493753 367177
rect 493791 367143 493801 367177
rect 493801 367143 493825 367177
rect 493863 367143 493869 367177
rect 493869 367143 493897 367177
rect 493935 367143 493937 367177
rect 493937 367143 493969 367177
rect 494007 367143 494039 367177
rect 494039 367143 494041 367177
rect 494079 367143 494107 367177
rect 494107 367143 494113 367177
rect 494151 367143 494175 367177
rect 494175 367143 494185 367177
rect 494223 367143 494243 367177
rect 494243 367143 494257 367177
rect 494295 367143 494311 367177
rect 494311 367143 494329 367177
rect 494367 367143 494379 367177
rect 494379 367143 494401 367177
rect 494439 367143 494447 367177
rect 494447 367143 494473 367177
rect 494511 367143 494515 367177
rect 494515 367143 494545 367177
rect 494583 367143 494617 367177
rect 493359 366685 493393 366719
rect 493431 366685 493461 366719
rect 493461 366685 493465 366719
rect 493503 366685 493529 366719
rect 493529 366685 493537 366719
rect 493575 366685 493597 366719
rect 493597 366685 493609 366719
rect 493647 366685 493665 366719
rect 493665 366685 493681 366719
rect 493719 366685 493733 366719
rect 493733 366685 493753 366719
rect 493791 366685 493801 366719
rect 493801 366685 493825 366719
rect 493863 366685 493869 366719
rect 493869 366685 493897 366719
rect 493935 366685 493937 366719
rect 493937 366685 493969 366719
rect 494007 366685 494039 366719
rect 494039 366685 494041 366719
rect 494079 366685 494107 366719
rect 494107 366685 494113 366719
rect 494151 366685 494175 366719
rect 494175 366685 494185 366719
rect 494223 366685 494243 366719
rect 494243 366685 494257 366719
rect 494295 366685 494311 366719
rect 494311 366685 494329 366719
rect 494367 366685 494379 366719
rect 494379 366685 494401 366719
rect 494439 366685 494447 366719
rect 494447 366685 494473 366719
rect 494511 366685 494515 366719
rect 494515 366685 494545 366719
rect 494583 366685 494617 366719
rect 493359 366227 493393 366261
rect 493431 366227 493461 366261
rect 493461 366227 493465 366261
rect 493503 366227 493529 366261
rect 493529 366227 493537 366261
rect 493575 366227 493597 366261
rect 493597 366227 493609 366261
rect 493647 366227 493665 366261
rect 493665 366227 493681 366261
rect 493719 366227 493733 366261
rect 493733 366227 493753 366261
rect 493791 366227 493801 366261
rect 493801 366227 493825 366261
rect 493863 366227 493869 366261
rect 493869 366227 493897 366261
rect 493935 366227 493937 366261
rect 493937 366227 493969 366261
rect 494007 366227 494039 366261
rect 494039 366227 494041 366261
rect 494079 366227 494107 366261
rect 494107 366227 494113 366261
rect 494151 366227 494175 366261
rect 494175 366227 494185 366261
rect 494223 366227 494243 366261
rect 494243 366227 494257 366261
rect 494295 366227 494311 366261
rect 494311 366227 494329 366261
rect 494367 366227 494379 366261
rect 494379 366227 494401 366261
rect 494439 366227 494447 366261
rect 494447 366227 494473 366261
rect 494511 366227 494515 366261
rect 494515 366227 494545 366261
rect 494583 366227 494617 366261
rect 493359 365769 493393 365803
rect 493431 365769 493461 365803
rect 493461 365769 493465 365803
rect 493503 365769 493529 365803
rect 493529 365769 493537 365803
rect 493575 365769 493597 365803
rect 493597 365769 493609 365803
rect 493647 365769 493665 365803
rect 493665 365769 493681 365803
rect 493719 365769 493733 365803
rect 493733 365769 493753 365803
rect 493791 365769 493801 365803
rect 493801 365769 493825 365803
rect 493863 365769 493869 365803
rect 493869 365769 493897 365803
rect 493935 365769 493937 365803
rect 493937 365769 493969 365803
rect 494007 365769 494039 365803
rect 494039 365769 494041 365803
rect 494079 365769 494107 365803
rect 494107 365769 494113 365803
rect 494151 365769 494175 365803
rect 494175 365769 494185 365803
rect 494223 365769 494243 365803
rect 494243 365769 494257 365803
rect 494295 365769 494311 365803
rect 494311 365769 494329 365803
rect 494367 365769 494379 365803
rect 494379 365769 494401 365803
rect 494439 365769 494447 365803
rect 494447 365769 494473 365803
rect 494511 365769 494515 365803
rect 494515 365769 494545 365803
rect 494583 365769 494617 365803
rect 493091 365507 493125 365541
rect 493091 365107 493125 365141
rect 493091 364707 493125 364741
rect 493359 365311 493393 365345
rect 493431 365311 493461 365345
rect 493461 365311 493465 365345
rect 493503 365311 493529 365345
rect 493529 365311 493537 365345
rect 493575 365311 493597 365345
rect 493597 365311 493609 365345
rect 493647 365311 493665 365345
rect 493665 365311 493681 365345
rect 493719 365311 493733 365345
rect 493733 365311 493753 365345
rect 493791 365311 493801 365345
rect 493801 365311 493825 365345
rect 493863 365311 493869 365345
rect 493869 365311 493897 365345
rect 493935 365311 493937 365345
rect 493937 365311 493969 365345
rect 494007 365311 494039 365345
rect 494039 365311 494041 365345
rect 494079 365311 494107 365345
rect 494107 365311 494113 365345
rect 494151 365311 494175 365345
rect 494175 365311 494185 365345
rect 494223 365311 494243 365345
rect 494243 365311 494257 365345
rect 494295 365311 494311 365345
rect 494311 365311 494329 365345
rect 494367 365311 494379 365345
rect 494379 365311 494401 365345
rect 494439 365311 494447 365345
rect 494447 365311 494473 365345
rect 494511 365311 494515 365345
rect 494515 365311 494545 365345
rect 494583 365311 494617 365345
rect 493359 364853 493393 364887
rect 493431 364853 493461 364887
rect 493461 364853 493465 364887
rect 493503 364853 493529 364887
rect 493529 364853 493537 364887
rect 493575 364853 493597 364887
rect 493597 364853 493609 364887
rect 493647 364853 493665 364887
rect 493665 364853 493681 364887
rect 493719 364853 493733 364887
rect 493733 364853 493753 364887
rect 493791 364853 493801 364887
rect 493801 364853 493825 364887
rect 493863 364853 493869 364887
rect 493869 364853 493897 364887
rect 493935 364853 493937 364887
rect 493937 364853 493969 364887
rect 494007 364853 494039 364887
rect 494039 364853 494041 364887
rect 494079 364853 494107 364887
rect 494107 364853 494113 364887
rect 494151 364853 494175 364887
rect 494175 364853 494185 364887
rect 494223 364853 494243 364887
rect 494243 364853 494257 364887
rect 494295 364853 494311 364887
rect 494311 364853 494329 364887
rect 494367 364853 494379 364887
rect 494379 364853 494401 364887
rect 494439 364853 494447 364887
rect 494447 364853 494473 364887
rect 494511 364853 494515 364887
rect 494515 364853 494545 364887
rect 494583 364853 494617 364887
rect 493091 364307 493125 364341
rect 493091 363907 493125 363941
rect 493091 363507 493125 363541
rect 493091 363107 493125 363141
rect 493091 362707 493125 362741
rect 493359 364395 493393 364429
rect 493431 364395 493461 364429
rect 493461 364395 493465 364429
rect 493503 364395 493529 364429
rect 493529 364395 493537 364429
rect 493575 364395 493597 364429
rect 493597 364395 493609 364429
rect 493647 364395 493665 364429
rect 493665 364395 493681 364429
rect 493719 364395 493733 364429
rect 493733 364395 493753 364429
rect 493791 364395 493801 364429
rect 493801 364395 493825 364429
rect 493863 364395 493869 364429
rect 493869 364395 493897 364429
rect 493935 364395 493937 364429
rect 493937 364395 493969 364429
rect 494007 364395 494039 364429
rect 494039 364395 494041 364429
rect 494079 364395 494107 364429
rect 494107 364395 494113 364429
rect 494151 364395 494175 364429
rect 494175 364395 494185 364429
rect 494223 364395 494243 364429
rect 494243 364395 494257 364429
rect 494295 364395 494311 364429
rect 494311 364395 494329 364429
rect 494367 364395 494379 364429
rect 494379 364395 494401 364429
rect 494439 364395 494447 364429
rect 494447 364395 494473 364429
rect 494511 364395 494515 364429
rect 494515 364395 494545 364429
rect 494583 364395 494617 364429
rect 493359 363937 493393 363971
rect 493431 363937 493461 363971
rect 493461 363937 493465 363971
rect 493503 363937 493529 363971
rect 493529 363937 493537 363971
rect 493575 363937 493597 363971
rect 493597 363937 493609 363971
rect 493647 363937 493665 363971
rect 493665 363937 493681 363971
rect 493719 363937 493733 363971
rect 493733 363937 493753 363971
rect 493791 363937 493801 363971
rect 493801 363937 493825 363971
rect 493863 363937 493869 363971
rect 493869 363937 493897 363971
rect 493935 363937 493937 363971
rect 493937 363937 493969 363971
rect 494007 363937 494039 363971
rect 494039 363937 494041 363971
rect 494079 363937 494107 363971
rect 494107 363937 494113 363971
rect 494151 363937 494175 363971
rect 494175 363937 494185 363971
rect 494223 363937 494243 363971
rect 494243 363937 494257 363971
rect 494295 363937 494311 363971
rect 494311 363937 494329 363971
rect 494367 363937 494379 363971
rect 494379 363937 494401 363971
rect 494439 363937 494447 363971
rect 494447 363937 494473 363971
rect 494511 363937 494515 363971
rect 494515 363937 494545 363971
rect 494583 363937 494617 363971
rect 493359 363479 493393 363513
rect 493431 363479 493461 363513
rect 493461 363479 493465 363513
rect 493503 363479 493529 363513
rect 493529 363479 493537 363513
rect 493575 363479 493597 363513
rect 493597 363479 493609 363513
rect 493647 363479 493665 363513
rect 493665 363479 493681 363513
rect 493719 363479 493733 363513
rect 493733 363479 493753 363513
rect 493791 363479 493801 363513
rect 493801 363479 493825 363513
rect 493863 363479 493869 363513
rect 493869 363479 493897 363513
rect 493935 363479 493937 363513
rect 493937 363479 493969 363513
rect 494007 363479 494039 363513
rect 494039 363479 494041 363513
rect 494079 363479 494107 363513
rect 494107 363479 494113 363513
rect 494151 363479 494175 363513
rect 494175 363479 494185 363513
rect 494223 363479 494243 363513
rect 494243 363479 494257 363513
rect 494295 363479 494311 363513
rect 494311 363479 494329 363513
rect 494367 363479 494379 363513
rect 494379 363479 494401 363513
rect 494439 363479 494447 363513
rect 494447 363479 494473 363513
rect 494511 363479 494515 363513
rect 494515 363479 494545 363513
rect 494583 363479 494617 363513
rect 493359 363021 493393 363055
rect 493431 363021 493461 363055
rect 493461 363021 493465 363055
rect 493503 363021 493529 363055
rect 493529 363021 493537 363055
rect 493575 363021 493597 363055
rect 493597 363021 493609 363055
rect 493647 363021 493665 363055
rect 493665 363021 493681 363055
rect 493719 363021 493733 363055
rect 493733 363021 493753 363055
rect 493791 363021 493801 363055
rect 493801 363021 493825 363055
rect 493863 363021 493869 363055
rect 493869 363021 493897 363055
rect 493935 363021 493937 363055
rect 493937 363021 493969 363055
rect 494007 363021 494039 363055
rect 494039 363021 494041 363055
rect 494079 363021 494107 363055
rect 494107 363021 494113 363055
rect 494151 363021 494175 363055
rect 494175 363021 494185 363055
rect 494223 363021 494243 363055
rect 494243 363021 494257 363055
rect 494295 363021 494311 363055
rect 494311 363021 494329 363055
rect 494367 363021 494379 363055
rect 494379 363021 494401 363055
rect 494439 363021 494447 363055
rect 494447 363021 494473 363055
rect 494511 363021 494515 363055
rect 494515 363021 494545 363055
rect 494583 363021 494617 363055
rect 493359 362563 493393 362597
rect 493431 362563 493461 362597
rect 493461 362563 493465 362597
rect 493503 362563 493529 362597
rect 493529 362563 493537 362597
rect 493575 362563 493597 362597
rect 493597 362563 493609 362597
rect 493647 362563 493665 362597
rect 493665 362563 493681 362597
rect 493719 362563 493733 362597
rect 493733 362563 493753 362597
rect 493791 362563 493801 362597
rect 493801 362563 493825 362597
rect 493863 362563 493869 362597
rect 493869 362563 493897 362597
rect 493935 362563 493937 362597
rect 493937 362563 493969 362597
rect 494007 362563 494039 362597
rect 494039 362563 494041 362597
rect 494079 362563 494107 362597
rect 494107 362563 494113 362597
rect 494151 362563 494175 362597
rect 494175 362563 494185 362597
rect 494223 362563 494243 362597
rect 494243 362563 494257 362597
rect 494295 362563 494311 362597
rect 494311 362563 494329 362597
rect 494367 362563 494379 362597
rect 494379 362563 494401 362597
rect 494439 362563 494447 362597
rect 494447 362563 494473 362597
rect 494511 362563 494515 362597
rect 494515 362563 494545 362597
rect 494583 362563 494617 362597
rect 494971 389907 495005 389941
rect 494971 389507 495005 389541
rect 494971 389107 495005 389141
rect 494971 388707 495005 388741
rect 494971 388307 495005 388341
rect 494971 387907 495005 387941
rect 494971 387507 495005 387541
rect 494971 387107 495005 387141
rect 494971 386707 495005 386741
rect 494971 386307 495005 386341
rect 494971 385907 495005 385941
rect 494971 385507 495005 385541
rect 494971 385107 495005 385141
rect 494971 384707 495005 384741
rect 494971 384307 495005 384341
rect 494971 383907 495005 383941
rect 494971 383507 495005 383541
rect 494971 383107 495005 383141
rect 494971 382707 495005 382741
rect 494971 382307 495005 382341
rect 494971 381907 495005 381941
rect 494971 381507 495005 381541
rect 494971 381107 495005 381141
rect 494971 380707 495005 380741
rect 494971 380307 495005 380341
rect 494971 379907 495005 379941
rect 494971 379507 495005 379541
rect 494971 379107 495005 379141
rect 494971 378707 495005 378741
rect 494971 378307 495005 378341
rect 494971 377907 495005 377941
rect 494971 377507 495005 377541
rect 494971 377107 495005 377141
rect 494971 376707 495005 376741
rect 494971 376307 495005 376341
rect 494971 375907 495005 375941
rect 494971 375507 495005 375541
rect 494971 375107 495005 375141
rect 494971 374707 495005 374741
rect 494971 374307 495005 374341
rect 494971 373907 495005 373941
rect 494971 373507 495005 373541
rect 494971 373107 495005 373141
rect 494971 372707 495005 372741
rect 494971 372307 495005 372341
rect 496851 390107 496885 390141
rect 497119 390683 497153 390717
rect 497191 390683 497221 390717
rect 497221 390683 497225 390717
rect 497263 390683 497289 390717
rect 497289 390683 497297 390717
rect 497335 390683 497357 390717
rect 497357 390683 497369 390717
rect 497407 390683 497425 390717
rect 497425 390683 497441 390717
rect 497479 390683 497493 390717
rect 497493 390683 497513 390717
rect 497551 390683 497561 390717
rect 497561 390683 497585 390717
rect 497623 390683 497629 390717
rect 497629 390683 497657 390717
rect 497695 390683 497697 390717
rect 497697 390683 497729 390717
rect 497767 390683 497799 390717
rect 497799 390683 497801 390717
rect 497839 390683 497867 390717
rect 497867 390683 497873 390717
rect 497911 390683 497935 390717
rect 497935 390683 497945 390717
rect 497983 390683 498003 390717
rect 498003 390683 498017 390717
rect 498055 390683 498071 390717
rect 498071 390683 498089 390717
rect 498127 390683 498139 390717
rect 498139 390683 498161 390717
rect 498199 390683 498207 390717
rect 498207 390683 498233 390717
rect 498271 390683 498275 390717
rect 498275 390683 498305 390717
rect 498343 390683 498377 390717
rect 497119 390225 497153 390259
rect 497191 390225 497221 390259
rect 497221 390225 497225 390259
rect 497263 390225 497289 390259
rect 497289 390225 497297 390259
rect 497335 390225 497357 390259
rect 497357 390225 497369 390259
rect 497407 390225 497425 390259
rect 497425 390225 497441 390259
rect 497479 390225 497493 390259
rect 497493 390225 497513 390259
rect 497551 390225 497561 390259
rect 497561 390225 497585 390259
rect 497623 390225 497629 390259
rect 497629 390225 497657 390259
rect 497695 390225 497697 390259
rect 497697 390225 497729 390259
rect 497767 390225 497799 390259
rect 497799 390225 497801 390259
rect 497839 390225 497867 390259
rect 497867 390225 497873 390259
rect 497911 390225 497935 390259
rect 497935 390225 497945 390259
rect 497983 390225 498003 390259
rect 498003 390225 498017 390259
rect 498055 390225 498071 390259
rect 498071 390225 498089 390259
rect 498127 390225 498139 390259
rect 498139 390225 498161 390259
rect 498199 390225 498207 390259
rect 498207 390225 498233 390259
rect 498271 390225 498275 390259
rect 498275 390225 498305 390259
rect 498343 390225 498377 390259
rect 496851 389707 496885 389741
rect 496851 389307 496885 389341
rect 496851 388907 496885 388941
rect 497119 389767 497153 389801
rect 497191 389767 497221 389801
rect 497221 389767 497225 389801
rect 497263 389767 497289 389801
rect 497289 389767 497297 389801
rect 497335 389767 497357 389801
rect 497357 389767 497369 389801
rect 497407 389767 497425 389801
rect 497425 389767 497441 389801
rect 497479 389767 497493 389801
rect 497493 389767 497513 389801
rect 497551 389767 497561 389801
rect 497561 389767 497585 389801
rect 497623 389767 497629 389801
rect 497629 389767 497657 389801
rect 497695 389767 497697 389801
rect 497697 389767 497729 389801
rect 497767 389767 497799 389801
rect 497799 389767 497801 389801
rect 497839 389767 497867 389801
rect 497867 389767 497873 389801
rect 497911 389767 497935 389801
rect 497935 389767 497945 389801
rect 497983 389767 498003 389801
rect 498003 389767 498017 389801
rect 498055 389767 498071 389801
rect 498071 389767 498089 389801
rect 498127 389767 498139 389801
rect 498139 389767 498161 389801
rect 498199 389767 498207 389801
rect 498207 389767 498233 389801
rect 498271 389767 498275 389801
rect 498275 389767 498305 389801
rect 498343 389767 498377 389801
rect 497119 389309 497153 389343
rect 497191 389309 497221 389343
rect 497221 389309 497225 389343
rect 497263 389309 497289 389343
rect 497289 389309 497297 389343
rect 497335 389309 497357 389343
rect 497357 389309 497369 389343
rect 497407 389309 497425 389343
rect 497425 389309 497441 389343
rect 497479 389309 497493 389343
rect 497493 389309 497513 389343
rect 497551 389309 497561 389343
rect 497561 389309 497585 389343
rect 497623 389309 497629 389343
rect 497629 389309 497657 389343
rect 497695 389309 497697 389343
rect 497697 389309 497729 389343
rect 497767 389309 497799 389343
rect 497799 389309 497801 389343
rect 497839 389309 497867 389343
rect 497867 389309 497873 389343
rect 497911 389309 497935 389343
rect 497935 389309 497945 389343
rect 497983 389309 498003 389343
rect 498003 389309 498017 389343
rect 498055 389309 498071 389343
rect 498071 389309 498089 389343
rect 498127 389309 498139 389343
rect 498139 389309 498161 389343
rect 498199 389309 498207 389343
rect 498207 389309 498233 389343
rect 498271 389309 498275 389343
rect 498275 389309 498305 389343
rect 498343 389309 498377 389343
rect 496851 388507 496885 388541
rect 497119 388851 497153 388885
rect 497191 388851 497221 388885
rect 497221 388851 497225 388885
rect 497263 388851 497289 388885
rect 497289 388851 497297 388885
rect 497335 388851 497357 388885
rect 497357 388851 497369 388885
rect 497407 388851 497425 388885
rect 497425 388851 497441 388885
rect 497479 388851 497493 388885
rect 497493 388851 497513 388885
rect 497551 388851 497561 388885
rect 497561 388851 497585 388885
rect 497623 388851 497629 388885
rect 497629 388851 497657 388885
rect 497695 388851 497697 388885
rect 497697 388851 497729 388885
rect 497767 388851 497799 388885
rect 497799 388851 497801 388885
rect 497839 388851 497867 388885
rect 497867 388851 497873 388885
rect 497911 388851 497935 388885
rect 497935 388851 497945 388885
rect 497983 388851 498003 388885
rect 498003 388851 498017 388885
rect 498055 388851 498071 388885
rect 498071 388851 498089 388885
rect 498127 388851 498139 388885
rect 498139 388851 498161 388885
rect 498199 388851 498207 388885
rect 498207 388851 498233 388885
rect 498271 388851 498275 388885
rect 498275 388851 498305 388885
rect 498343 388851 498377 388885
rect 497119 388393 497153 388427
rect 497191 388393 497221 388427
rect 497221 388393 497225 388427
rect 497263 388393 497289 388427
rect 497289 388393 497297 388427
rect 497335 388393 497357 388427
rect 497357 388393 497369 388427
rect 497407 388393 497425 388427
rect 497425 388393 497441 388427
rect 497479 388393 497493 388427
rect 497493 388393 497513 388427
rect 497551 388393 497561 388427
rect 497561 388393 497585 388427
rect 497623 388393 497629 388427
rect 497629 388393 497657 388427
rect 497695 388393 497697 388427
rect 497697 388393 497729 388427
rect 497767 388393 497799 388427
rect 497799 388393 497801 388427
rect 497839 388393 497867 388427
rect 497867 388393 497873 388427
rect 497911 388393 497935 388427
rect 497935 388393 497945 388427
rect 497983 388393 498003 388427
rect 498003 388393 498017 388427
rect 498055 388393 498071 388427
rect 498071 388393 498089 388427
rect 498127 388393 498139 388427
rect 498139 388393 498161 388427
rect 498199 388393 498207 388427
rect 498207 388393 498233 388427
rect 498271 388393 498275 388427
rect 498275 388393 498305 388427
rect 498343 388393 498377 388427
rect 496851 388107 496885 388141
rect 496851 387707 496885 387741
rect 496851 387307 496885 387341
rect 497119 387935 497153 387969
rect 497191 387935 497221 387969
rect 497221 387935 497225 387969
rect 497263 387935 497289 387969
rect 497289 387935 497297 387969
rect 497335 387935 497357 387969
rect 497357 387935 497369 387969
rect 497407 387935 497425 387969
rect 497425 387935 497441 387969
rect 497479 387935 497493 387969
rect 497493 387935 497513 387969
rect 497551 387935 497561 387969
rect 497561 387935 497585 387969
rect 497623 387935 497629 387969
rect 497629 387935 497657 387969
rect 497695 387935 497697 387969
rect 497697 387935 497729 387969
rect 497767 387935 497799 387969
rect 497799 387935 497801 387969
rect 497839 387935 497867 387969
rect 497867 387935 497873 387969
rect 497911 387935 497935 387969
rect 497935 387935 497945 387969
rect 497983 387935 498003 387969
rect 498003 387935 498017 387969
rect 498055 387935 498071 387969
rect 498071 387935 498089 387969
rect 498127 387935 498139 387969
rect 498139 387935 498161 387969
rect 498199 387935 498207 387969
rect 498207 387935 498233 387969
rect 498271 387935 498275 387969
rect 498275 387935 498305 387969
rect 498343 387935 498377 387969
rect 497119 387477 497153 387511
rect 497191 387477 497221 387511
rect 497221 387477 497225 387511
rect 497263 387477 497289 387511
rect 497289 387477 497297 387511
rect 497335 387477 497357 387511
rect 497357 387477 497369 387511
rect 497407 387477 497425 387511
rect 497425 387477 497441 387511
rect 497479 387477 497493 387511
rect 497493 387477 497513 387511
rect 497551 387477 497561 387511
rect 497561 387477 497585 387511
rect 497623 387477 497629 387511
rect 497629 387477 497657 387511
rect 497695 387477 497697 387511
rect 497697 387477 497729 387511
rect 497767 387477 497799 387511
rect 497799 387477 497801 387511
rect 497839 387477 497867 387511
rect 497867 387477 497873 387511
rect 497911 387477 497935 387511
rect 497935 387477 497945 387511
rect 497983 387477 498003 387511
rect 498003 387477 498017 387511
rect 498055 387477 498071 387511
rect 498071 387477 498089 387511
rect 498127 387477 498139 387511
rect 498139 387477 498161 387511
rect 498199 387477 498207 387511
rect 498207 387477 498233 387511
rect 498271 387477 498275 387511
rect 498275 387477 498305 387511
rect 498343 387477 498377 387511
rect 496851 386907 496885 386941
rect 496851 386507 496885 386541
rect 496851 386107 496885 386141
rect 497119 387019 497153 387053
rect 497191 387019 497221 387053
rect 497221 387019 497225 387053
rect 497263 387019 497289 387053
rect 497289 387019 497297 387053
rect 497335 387019 497357 387053
rect 497357 387019 497369 387053
rect 497407 387019 497425 387053
rect 497425 387019 497441 387053
rect 497479 387019 497493 387053
rect 497493 387019 497513 387053
rect 497551 387019 497561 387053
rect 497561 387019 497585 387053
rect 497623 387019 497629 387053
rect 497629 387019 497657 387053
rect 497695 387019 497697 387053
rect 497697 387019 497729 387053
rect 497767 387019 497799 387053
rect 497799 387019 497801 387053
rect 497839 387019 497867 387053
rect 497867 387019 497873 387053
rect 497911 387019 497935 387053
rect 497935 387019 497945 387053
rect 497983 387019 498003 387053
rect 498003 387019 498017 387053
rect 498055 387019 498071 387053
rect 498071 387019 498089 387053
rect 498127 387019 498139 387053
rect 498139 387019 498161 387053
rect 498199 387019 498207 387053
rect 498207 387019 498233 387053
rect 498271 387019 498275 387053
rect 498275 387019 498305 387053
rect 498343 387019 498377 387053
rect 497119 386561 497153 386595
rect 497191 386561 497221 386595
rect 497221 386561 497225 386595
rect 497263 386561 497289 386595
rect 497289 386561 497297 386595
rect 497335 386561 497357 386595
rect 497357 386561 497369 386595
rect 497407 386561 497425 386595
rect 497425 386561 497441 386595
rect 497479 386561 497493 386595
rect 497493 386561 497513 386595
rect 497551 386561 497561 386595
rect 497561 386561 497585 386595
rect 497623 386561 497629 386595
rect 497629 386561 497657 386595
rect 497695 386561 497697 386595
rect 497697 386561 497729 386595
rect 497767 386561 497799 386595
rect 497799 386561 497801 386595
rect 497839 386561 497867 386595
rect 497867 386561 497873 386595
rect 497911 386561 497935 386595
rect 497935 386561 497945 386595
rect 497983 386561 498003 386595
rect 498003 386561 498017 386595
rect 498055 386561 498071 386595
rect 498071 386561 498089 386595
rect 498127 386561 498139 386595
rect 498139 386561 498161 386595
rect 498199 386561 498207 386595
rect 498207 386561 498233 386595
rect 498271 386561 498275 386595
rect 498275 386561 498305 386595
rect 498343 386561 498377 386595
rect 496851 385707 496885 385741
rect 496851 385307 496885 385341
rect 496851 384907 496885 384941
rect 497119 386103 497153 386137
rect 497191 386103 497221 386137
rect 497221 386103 497225 386137
rect 497263 386103 497289 386137
rect 497289 386103 497297 386137
rect 497335 386103 497357 386137
rect 497357 386103 497369 386137
rect 497407 386103 497425 386137
rect 497425 386103 497441 386137
rect 497479 386103 497493 386137
rect 497493 386103 497513 386137
rect 497551 386103 497561 386137
rect 497561 386103 497585 386137
rect 497623 386103 497629 386137
rect 497629 386103 497657 386137
rect 497695 386103 497697 386137
rect 497697 386103 497729 386137
rect 497767 386103 497799 386137
rect 497799 386103 497801 386137
rect 497839 386103 497867 386137
rect 497867 386103 497873 386137
rect 497911 386103 497935 386137
rect 497935 386103 497945 386137
rect 497983 386103 498003 386137
rect 498003 386103 498017 386137
rect 498055 386103 498071 386137
rect 498071 386103 498089 386137
rect 498127 386103 498139 386137
rect 498139 386103 498161 386137
rect 498199 386103 498207 386137
rect 498207 386103 498233 386137
rect 498271 386103 498275 386137
rect 498275 386103 498305 386137
rect 498343 386103 498377 386137
rect 497119 385645 497153 385679
rect 497191 385645 497221 385679
rect 497221 385645 497225 385679
rect 497263 385645 497289 385679
rect 497289 385645 497297 385679
rect 497335 385645 497357 385679
rect 497357 385645 497369 385679
rect 497407 385645 497425 385679
rect 497425 385645 497441 385679
rect 497479 385645 497493 385679
rect 497493 385645 497513 385679
rect 497551 385645 497561 385679
rect 497561 385645 497585 385679
rect 497623 385645 497629 385679
rect 497629 385645 497657 385679
rect 497695 385645 497697 385679
rect 497697 385645 497729 385679
rect 497767 385645 497799 385679
rect 497799 385645 497801 385679
rect 497839 385645 497867 385679
rect 497867 385645 497873 385679
rect 497911 385645 497935 385679
rect 497935 385645 497945 385679
rect 497983 385645 498003 385679
rect 498003 385645 498017 385679
rect 498055 385645 498071 385679
rect 498071 385645 498089 385679
rect 498127 385645 498139 385679
rect 498139 385645 498161 385679
rect 498199 385645 498207 385679
rect 498207 385645 498233 385679
rect 498271 385645 498275 385679
rect 498275 385645 498305 385679
rect 498343 385645 498377 385679
rect 497119 385187 497153 385221
rect 497191 385187 497221 385221
rect 497221 385187 497225 385221
rect 497263 385187 497289 385221
rect 497289 385187 497297 385221
rect 497335 385187 497357 385221
rect 497357 385187 497369 385221
rect 497407 385187 497425 385221
rect 497425 385187 497441 385221
rect 497479 385187 497493 385221
rect 497493 385187 497513 385221
rect 497551 385187 497561 385221
rect 497561 385187 497585 385221
rect 497623 385187 497629 385221
rect 497629 385187 497657 385221
rect 497695 385187 497697 385221
rect 497697 385187 497729 385221
rect 497767 385187 497799 385221
rect 497799 385187 497801 385221
rect 497839 385187 497867 385221
rect 497867 385187 497873 385221
rect 497911 385187 497935 385221
rect 497935 385187 497945 385221
rect 497983 385187 498003 385221
rect 498003 385187 498017 385221
rect 498055 385187 498071 385221
rect 498071 385187 498089 385221
rect 498127 385187 498139 385221
rect 498139 385187 498161 385221
rect 498199 385187 498207 385221
rect 498207 385187 498233 385221
rect 498271 385187 498275 385221
rect 498275 385187 498305 385221
rect 498343 385187 498377 385221
rect 497119 384729 497153 384763
rect 497191 384729 497221 384763
rect 497221 384729 497225 384763
rect 497263 384729 497289 384763
rect 497289 384729 497297 384763
rect 497335 384729 497357 384763
rect 497357 384729 497369 384763
rect 497407 384729 497425 384763
rect 497425 384729 497441 384763
rect 497479 384729 497493 384763
rect 497493 384729 497513 384763
rect 497551 384729 497561 384763
rect 497561 384729 497585 384763
rect 497623 384729 497629 384763
rect 497629 384729 497657 384763
rect 497695 384729 497697 384763
rect 497697 384729 497729 384763
rect 497767 384729 497799 384763
rect 497799 384729 497801 384763
rect 497839 384729 497867 384763
rect 497867 384729 497873 384763
rect 497911 384729 497935 384763
rect 497935 384729 497945 384763
rect 497983 384729 498003 384763
rect 498003 384729 498017 384763
rect 498055 384729 498071 384763
rect 498071 384729 498089 384763
rect 498127 384729 498139 384763
rect 498139 384729 498161 384763
rect 498199 384729 498207 384763
rect 498207 384729 498233 384763
rect 498271 384729 498275 384763
rect 498275 384729 498305 384763
rect 498343 384729 498377 384763
rect 496851 384507 496885 384541
rect 496851 384107 496885 384141
rect 496851 383707 496885 383741
rect 497119 384271 497153 384305
rect 497191 384271 497221 384305
rect 497221 384271 497225 384305
rect 497263 384271 497289 384305
rect 497289 384271 497297 384305
rect 497335 384271 497357 384305
rect 497357 384271 497369 384305
rect 497407 384271 497425 384305
rect 497425 384271 497441 384305
rect 497479 384271 497493 384305
rect 497493 384271 497513 384305
rect 497551 384271 497561 384305
rect 497561 384271 497585 384305
rect 497623 384271 497629 384305
rect 497629 384271 497657 384305
rect 497695 384271 497697 384305
rect 497697 384271 497729 384305
rect 497767 384271 497799 384305
rect 497799 384271 497801 384305
rect 497839 384271 497867 384305
rect 497867 384271 497873 384305
rect 497911 384271 497935 384305
rect 497935 384271 497945 384305
rect 497983 384271 498003 384305
rect 498003 384271 498017 384305
rect 498055 384271 498071 384305
rect 498071 384271 498089 384305
rect 498127 384271 498139 384305
rect 498139 384271 498161 384305
rect 498199 384271 498207 384305
rect 498207 384271 498233 384305
rect 498271 384271 498275 384305
rect 498275 384271 498305 384305
rect 498343 384271 498377 384305
rect 497119 383813 497153 383847
rect 497191 383813 497221 383847
rect 497221 383813 497225 383847
rect 497263 383813 497289 383847
rect 497289 383813 497297 383847
rect 497335 383813 497357 383847
rect 497357 383813 497369 383847
rect 497407 383813 497425 383847
rect 497425 383813 497441 383847
rect 497479 383813 497493 383847
rect 497493 383813 497513 383847
rect 497551 383813 497561 383847
rect 497561 383813 497585 383847
rect 497623 383813 497629 383847
rect 497629 383813 497657 383847
rect 497695 383813 497697 383847
rect 497697 383813 497729 383847
rect 497767 383813 497799 383847
rect 497799 383813 497801 383847
rect 497839 383813 497867 383847
rect 497867 383813 497873 383847
rect 497911 383813 497935 383847
rect 497935 383813 497945 383847
rect 497983 383813 498003 383847
rect 498003 383813 498017 383847
rect 498055 383813 498071 383847
rect 498071 383813 498089 383847
rect 498127 383813 498139 383847
rect 498139 383813 498161 383847
rect 498199 383813 498207 383847
rect 498207 383813 498233 383847
rect 498271 383813 498275 383847
rect 498275 383813 498305 383847
rect 498343 383813 498377 383847
rect 496851 383307 496885 383341
rect 496851 382907 496885 382941
rect 496851 382507 496885 382541
rect 496851 382107 496885 382141
rect 497119 383355 497153 383389
rect 497191 383355 497221 383389
rect 497221 383355 497225 383389
rect 497263 383355 497289 383389
rect 497289 383355 497297 383389
rect 497335 383355 497357 383389
rect 497357 383355 497369 383389
rect 497407 383355 497425 383389
rect 497425 383355 497441 383389
rect 497479 383355 497493 383389
rect 497493 383355 497513 383389
rect 497551 383355 497561 383389
rect 497561 383355 497585 383389
rect 497623 383355 497629 383389
rect 497629 383355 497657 383389
rect 497695 383355 497697 383389
rect 497697 383355 497729 383389
rect 497767 383355 497799 383389
rect 497799 383355 497801 383389
rect 497839 383355 497867 383389
rect 497867 383355 497873 383389
rect 497911 383355 497935 383389
rect 497935 383355 497945 383389
rect 497983 383355 498003 383389
rect 498003 383355 498017 383389
rect 498055 383355 498071 383389
rect 498071 383355 498089 383389
rect 498127 383355 498139 383389
rect 498139 383355 498161 383389
rect 498199 383355 498207 383389
rect 498207 383355 498233 383389
rect 498271 383355 498275 383389
rect 498275 383355 498305 383389
rect 498343 383355 498377 383389
rect 497119 382897 497153 382931
rect 497191 382897 497221 382931
rect 497221 382897 497225 382931
rect 497263 382897 497289 382931
rect 497289 382897 497297 382931
rect 497335 382897 497357 382931
rect 497357 382897 497369 382931
rect 497407 382897 497425 382931
rect 497425 382897 497441 382931
rect 497479 382897 497493 382931
rect 497493 382897 497513 382931
rect 497551 382897 497561 382931
rect 497561 382897 497585 382931
rect 497623 382897 497629 382931
rect 497629 382897 497657 382931
rect 497695 382897 497697 382931
rect 497697 382897 497729 382931
rect 497767 382897 497799 382931
rect 497799 382897 497801 382931
rect 497839 382897 497867 382931
rect 497867 382897 497873 382931
rect 497911 382897 497935 382931
rect 497935 382897 497945 382931
rect 497983 382897 498003 382931
rect 498003 382897 498017 382931
rect 498055 382897 498071 382931
rect 498071 382897 498089 382931
rect 498127 382897 498139 382931
rect 498139 382897 498161 382931
rect 498199 382897 498207 382931
rect 498207 382897 498233 382931
rect 498271 382897 498275 382931
rect 498275 382897 498305 382931
rect 498343 382897 498377 382931
rect 497119 382439 497153 382473
rect 497191 382439 497221 382473
rect 497221 382439 497225 382473
rect 497263 382439 497289 382473
rect 497289 382439 497297 382473
rect 497335 382439 497357 382473
rect 497357 382439 497369 382473
rect 497407 382439 497425 382473
rect 497425 382439 497441 382473
rect 497479 382439 497493 382473
rect 497493 382439 497513 382473
rect 497551 382439 497561 382473
rect 497561 382439 497585 382473
rect 497623 382439 497629 382473
rect 497629 382439 497657 382473
rect 497695 382439 497697 382473
rect 497697 382439 497729 382473
rect 497767 382439 497799 382473
rect 497799 382439 497801 382473
rect 497839 382439 497867 382473
rect 497867 382439 497873 382473
rect 497911 382439 497935 382473
rect 497935 382439 497945 382473
rect 497983 382439 498003 382473
rect 498003 382439 498017 382473
rect 498055 382439 498071 382473
rect 498071 382439 498089 382473
rect 498127 382439 498139 382473
rect 498139 382439 498161 382473
rect 498199 382439 498207 382473
rect 498207 382439 498233 382473
rect 498271 382439 498275 382473
rect 498275 382439 498305 382473
rect 498343 382439 498377 382473
rect 497119 381981 497153 382015
rect 497191 381981 497221 382015
rect 497221 381981 497225 382015
rect 497263 381981 497289 382015
rect 497289 381981 497297 382015
rect 497335 381981 497357 382015
rect 497357 381981 497369 382015
rect 497407 381981 497425 382015
rect 497425 381981 497441 382015
rect 497479 381981 497493 382015
rect 497493 381981 497513 382015
rect 497551 381981 497561 382015
rect 497561 381981 497585 382015
rect 497623 381981 497629 382015
rect 497629 381981 497657 382015
rect 497695 381981 497697 382015
rect 497697 381981 497729 382015
rect 497767 381981 497799 382015
rect 497799 381981 497801 382015
rect 497839 381981 497867 382015
rect 497867 381981 497873 382015
rect 497911 381981 497935 382015
rect 497935 381981 497945 382015
rect 497983 381981 498003 382015
rect 498003 381981 498017 382015
rect 498055 381981 498071 382015
rect 498071 381981 498089 382015
rect 498127 381981 498139 382015
rect 498139 381981 498161 382015
rect 498199 381981 498207 382015
rect 498207 381981 498233 382015
rect 498271 381981 498275 382015
rect 498275 381981 498305 382015
rect 498343 381981 498377 382015
rect 496851 381707 496885 381741
rect 496851 381307 496885 381341
rect 496851 380907 496885 380941
rect 497119 381523 497153 381557
rect 497191 381523 497221 381557
rect 497221 381523 497225 381557
rect 497263 381523 497289 381557
rect 497289 381523 497297 381557
rect 497335 381523 497357 381557
rect 497357 381523 497369 381557
rect 497407 381523 497425 381557
rect 497425 381523 497441 381557
rect 497479 381523 497493 381557
rect 497493 381523 497513 381557
rect 497551 381523 497561 381557
rect 497561 381523 497585 381557
rect 497623 381523 497629 381557
rect 497629 381523 497657 381557
rect 497695 381523 497697 381557
rect 497697 381523 497729 381557
rect 497767 381523 497799 381557
rect 497799 381523 497801 381557
rect 497839 381523 497867 381557
rect 497867 381523 497873 381557
rect 497911 381523 497935 381557
rect 497935 381523 497945 381557
rect 497983 381523 498003 381557
rect 498003 381523 498017 381557
rect 498055 381523 498071 381557
rect 498071 381523 498089 381557
rect 498127 381523 498139 381557
rect 498139 381523 498161 381557
rect 498199 381523 498207 381557
rect 498207 381523 498233 381557
rect 498271 381523 498275 381557
rect 498275 381523 498305 381557
rect 498343 381523 498377 381557
rect 497119 381065 497153 381099
rect 497191 381065 497221 381099
rect 497221 381065 497225 381099
rect 497263 381065 497289 381099
rect 497289 381065 497297 381099
rect 497335 381065 497357 381099
rect 497357 381065 497369 381099
rect 497407 381065 497425 381099
rect 497425 381065 497441 381099
rect 497479 381065 497493 381099
rect 497493 381065 497513 381099
rect 497551 381065 497561 381099
rect 497561 381065 497585 381099
rect 497623 381065 497629 381099
rect 497629 381065 497657 381099
rect 497695 381065 497697 381099
rect 497697 381065 497729 381099
rect 497767 381065 497799 381099
rect 497799 381065 497801 381099
rect 497839 381065 497867 381099
rect 497867 381065 497873 381099
rect 497911 381065 497935 381099
rect 497935 381065 497945 381099
rect 497983 381065 498003 381099
rect 498003 381065 498017 381099
rect 498055 381065 498071 381099
rect 498071 381065 498089 381099
rect 498127 381065 498139 381099
rect 498139 381065 498161 381099
rect 498199 381065 498207 381099
rect 498207 381065 498233 381099
rect 498271 381065 498275 381099
rect 498275 381065 498305 381099
rect 498343 381065 498377 381099
rect 496851 380507 496885 380541
rect 496851 380107 496885 380141
rect 496851 379707 496885 379741
rect 497119 380607 497153 380641
rect 497191 380607 497221 380641
rect 497221 380607 497225 380641
rect 497263 380607 497289 380641
rect 497289 380607 497297 380641
rect 497335 380607 497357 380641
rect 497357 380607 497369 380641
rect 497407 380607 497425 380641
rect 497425 380607 497441 380641
rect 497479 380607 497493 380641
rect 497493 380607 497513 380641
rect 497551 380607 497561 380641
rect 497561 380607 497585 380641
rect 497623 380607 497629 380641
rect 497629 380607 497657 380641
rect 497695 380607 497697 380641
rect 497697 380607 497729 380641
rect 497767 380607 497799 380641
rect 497799 380607 497801 380641
rect 497839 380607 497867 380641
rect 497867 380607 497873 380641
rect 497911 380607 497935 380641
rect 497935 380607 497945 380641
rect 497983 380607 498003 380641
rect 498003 380607 498017 380641
rect 498055 380607 498071 380641
rect 498071 380607 498089 380641
rect 498127 380607 498139 380641
rect 498139 380607 498161 380641
rect 498199 380607 498207 380641
rect 498207 380607 498233 380641
rect 498271 380607 498275 380641
rect 498275 380607 498305 380641
rect 498343 380607 498377 380641
rect 497119 380149 497153 380183
rect 497191 380149 497221 380183
rect 497221 380149 497225 380183
rect 497263 380149 497289 380183
rect 497289 380149 497297 380183
rect 497335 380149 497357 380183
rect 497357 380149 497369 380183
rect 497407 380149 497425 380183
rect 497425 380149 497441 380183
rect 497479 380149 497493 380183
rect 497493 380149 497513 380183
rect 497551 380149 497561 380183
rect 497561 380149 497585 380183
rect 497623 380149 497629 380183
rect 497629 380149 497657 380183
rect 497695 380149 497697 380183
rect 497697 380149 497729 380183
rect 497767 380149 497799 380183
rect 497799 380149 497801 380183
rect 497839 380149 497867 380183
rect 497867 380149 497873 380183
rect 497911 380149 497935 380183
rect 497935 380149 497945 380183
rect 497983 380149 498003 380183
rect 498003 380149 498017 380183
rect 498055 380149 498071 380183
rect 498071 380149 498089 380183
rect 498127 380149 498139 380183
rect 498139 380149 498161 380183
rect 498199 380149 498207 380183
rect 498207 380149 498233 380183
rect 498271 380149 498275 380183
rect 498275 380149 498305 380183
rect 498343 380149 498377 380183
rect 496851 379307 496885 379341
rect 496851 378907 496885 378941
rect 496851 378507 496885 378541
rect 497119 379691 497153 379725
rect 497191 379691 497221 379725
rect 497221 379691 497225 379725
rect 497263 379691 497289 379725
rect 497289 379691 497297 379725
rect 497335 379691 497357 379725
rect 497357 379691 497369 379725
rect 497407 379691 497425 379725
rect 497425 379691 497441 379725
rect 497479 379691 497493 379725
rect 497493 379691 497513 379725
rect 497551 379691 497561 379725
rect 497561 379691 497585 379725
rect 497623 379691 497629 379725
rect 497629 379691 497657 379725
rect 497695 379691 497697 379725
rect 497697 379691 497729 379725
rect 497767 379691 497799 379725
rect 497799 379691 497801 379725
rect 497839 379691 497867 379725
rect 497867 379691 497873 379725
rect 497911 379691 497935 379725
rect 497935 379691 497945 379725
rect 497983 379691 498003 379725
rect 498003 379691 498017 379725
rect 498055 379691 498071 379725
rect 498071 379691 498089 379725
rect 498127 379691 498139 379725
rect 498139 379691 498161 379725
rect 498199 379691 498207 379725
rect 498207 379691 498233 379725
rect 498271 379691 498275 379725
rect 498275 379691 498305 379725
rect 498343 379691 498377 379725
rect 497119 379233 497153 379267
rect 497191 379233 497221 379267
rect 497221 379233 497225 379267
rect 497263 379233 497289 379267
rect 497289 379233 497297 379267
rect 497335 379233 497357 379267
rect 497357 379233 497369 379267
rect 497407 379233 497425 379267
rect 497425 379233 497441 379267
rect 497479 379233 497493 379267
rect 497493 379233 497513 379267
rect 497551 379233 497561 379267
rect 497561 379233 497585 379267
rect 497623 379233 497629 379267
rect 497629 379233 497657 379267
rect 497695 379233 497697 379267
rect 497697 379233 497729 379267
rect 497767 379233 497799 379267
rect 497799 379233 497801 379267
rect 497839 379233 497867 379267
rect 497867 379233 497873 379267
rect 497911 379233 497935 379267
rect 497935 379233 497945 379267
rect 497983 379233 498003 379267
rect 498003 379233 498017 379267
rect 498055 379233 498071 379267
rect 498071 379233 498089 379267
rect 498127 379233 498139 379267
rect 498139 379233 498161 379267
rect 498199 379233 498207 379267
rect 498207 379233 498233 379267
rect 498271 379233 498275 379267
rect 498275 379233 498305 379267
rect 498343 379233 498377 379267
rect 497119 378775 497153 378809
rect 497191 378775 497221 378809
rect 497221 378775 497225 378809
rect 497263 378775 497289 378809
rect 497289 378775 497297 378809
rect 497335 378775 497357 378809
rect 497357 378775 497369 378809
rect 497407 378775 497425 378809
rect 497425 378775 497441 378809
rect 497479 378775 497493 378809
rect 497493 378775 497513 378809
rect 497551 378775 497561 378809
rect 497561 378775 497585 378809
rect 497623 378775 497629 378809
rect 497629 378775 497657 378809
rect 497695 378775 497697 378809
rect 497697 378775 497729 378809
rect 497767 378775 497799 378809
rect 497799 378775 497801 378809
rect 497839 378775 497867 378809
rect 497867 378775 497873 378809
rect 497911 378775 497935 378809
rect 497935 378775 497945 378809
rect 497983 378775 498003 378809
rect 498003 378775 498017 378809
rect 498055 378775 498071 378809
rect 498071 378775 498089 378809
rect 498127 378775 498139 378809
rect 498139 378775 498161 378809
rect 498199 378775 498207 378809
rect 498207 378775 498233 378809
rect 498271 378775 498275 378809
rect 498275 378775 498305 378809
rect 498343 378775 498377 378809
rect 497119 378317 497153 378351
rect 497191 378317 497221 378351
rect 497221 378317 497225 378351
rect 497263 378317 497289 378351
rect 497289 378317 497297 378351
rect 497335 378317 497357 378351
rect 497357 378317 497369 378351
rect 497407 378317 497425 378351
rect 497425 378317 497441 378351
rect 497479 378317 497493 378351
rect 497493 378317 497513 378351
rect 497551 378317 497561 378351
rect 497561 378317 497585 378351
rect 497623 378317 497629 378351
rect 497629 378317 497657 378351
rect 497695 378317 497697 378351
rect 497697 378317 497729 378351
rect 497767 378317 497799 378351
rect 497799 378317 497801 378351
rect 497839 378317 497867 378351
rect 497867 378317 497873 378351
rect 497911 378317 497935 378351
rect 497935 378317 497945 378351
rect 497983 378317 498003 378351
rect 498003 378317 498017 378351
rect 498055 378317 498071 378351
rect 498071 378317 498089 378351
rect 498127 378317 498139 378351
rect 498139 378317 498161 378351
rect 498199 378317 498207 378351
rect 498207 378317 498233 378351
rect 498271 378317 498275 378351
rect 498275 378317 498305 378351
rect 498343 378317 498377 378351
rect 496851 378107 496885 378141
rect 496851 377707 496885 377741
rect 496851 377307 496885 377341
rect 496851 376907 496885 376941
rect 497119 377859 497153 377893
rect 497191 377859 497221 377893
rect 497221 377859 497225 377893
rect 497263 377859 497289 377893
rect 497289 377859 497297 377893
rect 497335 377859 497357 377893
rect 497357 377859 497369 377893
rect 497407 377859 497425 377893
rect 497425 377859 497441 377893
rect 497479 377859 497493 377893
rect 497493 377859 497513 377893
rect 497551 377859 497561 377893
rect 497561 377859 497585 377893
rect 497623 377859 497629 377893
rect 497629 377859 497657 377893
rect 497695 377859 497697 377893
rect 497697 377859 497729 377893
rect 497767 377859 497799 377893
rect 497799 377859 497801 377893
rect 497839 377859 497867 377893
rect 497867 377859 497873 377893
rect 497911 377859 497935 377893
rect 497935 377859 497945 377893
rect 497983 377859 498003 377893
rect 498003 377859 498017 377893
rect 498055 377859 498071 377893
rect 498071 377859 498089 377893
rect 498127 377859 498139 377893
rect 498139 377859 498161 377893
rect 498199 377859 498207 377893
rect 498207 377859 498233 377893
rect 498271 377859 498275 377893
rect 498275 377859 498305 377893
rect 498343 377859 498377 377893
rect 497119 377401 497153 377435
rect 497191 377401 497221 377435
rect 497221 377401 497225 377435
rect 497263 377401 497289 377435
rect 497289 377401 497297 377435
rect 497335 377401 497357 377435
rect 497357 377401 497369 377435
rect 497407 377401 497425 377435
rect 497425 377401 497441 377435
rect 497479 377401 497493 377435
rect 497493 377401 497513 377435
rect 497551 377401 497561 377435
rect 497561 377401 497585 377435
rect 497623 377401 497629 377435
rect 497629 377401 497657 377435
rect 497695 377401 497697 377435
rect 497697 377401 497729 377435
rect 497767 377401 497799 377435
rect 497799 377401 497801 377435
rect 497839 377401 497867 377435
rect 497867 377401 497873 377435
rect 497911 377401 497935 377435
rect 497935 377401 497945 377435
rect 497983 377401 498003 377435
rect 498003 377401 498017 377435
rect 498055 377401 498071 377435
rect 498071 377401 498089 377435
rect 498127 377401 498139 377435
rect 498139 377401 498161 377435
rect 498199 377401 498207 377435
rect 498207 377401 498233 377435
rect 498271 377401 498275 377435
rect 498275 377401 498305 377435
rect 498343 377401 498377 377435
rect 496851 376507 496885 376541
rect 496851 376107 496885 376141
rect 496851 375707 496885 375741
rect 497119 376943 497153 376977
rect 497191 376943 497221 376977
rect 497221 376943 497225 376977
rect 497263 376943 497289 376977
rect 497289 376943 497297 376977
rect 497335 376943 497357 376977
rect 497357 376943 497369 376977
rect 497407 376943 497425 376977
rect 497425 376943 497441 376977
rect 497479 376943 497493 376977
rect 497493 376943 497513 376977
rect 497551 376943 497561 376977
rect 497561 376943 497585 376977
rect 497623 376943 497629 376977
rect 497629 376943 497657 376977
rect 497695 376943 497697 376977
rect 497697 376943 497729 376977
rect 497767 376943 497799 376977
rect 497799 376943 497801 376977
rect 497839 376943 497867 376977
rect 497867 376943 497873 376977
rect 497911 376943 497935 376977
rect 497935 376943 497945 376977
rect 497983 376943 498003 376977
rect 498003 376943 498017 376977
rect 498055 376943 498071 376977
rect 498071 376943 498089 376977
rect 498127 376943 498139 376977
rect 498139 376943 498161 376977
rect 498199 376943 498207 376977
rect 498207 376943 498233 376977
rect 498271 376943 498275 376977
rect 498275 376943 498305 376977
rect 498343 376943 498377 376977
rect 497119 376485 497153 376519
rect 497191 376485 497221 376519
rect 497221 376485 497225 376519
rect 497263 376485 497289 376519
rect 497289 376485 497297 376519
rect 497335 376485 497357 376519
rect 497357 376485 497369 376519
rect 497407 376485 497425 376519
rect 497425 376485 497441 376519
rect 497479 376485 497493 376519
rect 497493 376485 497513 376519
rect 497551 376485 497561 376519
rect 497561 376485 497585 376519
rect 497623 376485 497629 376519
rect 497629 376485 497657 376519
rect 497695 376485 497697 376519
rect 497697 376485 497729 376519
rect 497767 376485 497799 376519
rect 497799 376485 497801 376519
rect 497839 376485 497867 376519
rect 497867 376485 497873 376519
rect 497911 376485 497935 376519
rect 497935 376485 497945 376519
rect 497983 376485 498003 376519
rect 498003 376485 498017 376519
rect 498055 376485 498071 376519
rect 498071 376485 498089 376519
rect 498127 376485 498139 376519
rect 498139 376485 498161 376519
rect 498199 376485 498207 376519
rect 498207 376485 498233 376519
rect 498271 376485 498275 376519
rect 498275 376485 498305 376519
rect 498343 376485 498377 376519
rect 497119 376027 497153 376061
rect 497191 376027 497221 376061
rect 497221 376027 497225 376061
rect 497263 376027 497289 376061
rect 497289 376027 497297 376061
rect 497335 376027 497357 376061
rect 497357 376027 497369 376061
rect 497407 376027 497425 376061
rect 497425 376027 497441 376061
rect 497479 376027 497493 376061
rect 497493 376027 497513 376061
rect 497551 376027 497561 376061
rect 497561 376027 497585 376061
rect 497623 376027 497629 376061
rect 497629 376027 497657 376061
rect 497695 376027 497697 376061
rect 497697 376027 497729 376061
rect 497767 376027 497799 376061
rect 497799 376027 497801 376061
rect 497839 376027 497867 376061
rect 497867 376027 497873 376061
rect 497911 376027 497935 376061
rect 497935 376027 497945 376061
rect 497983 376027 498003 376061
rect 498003 376027 498017 376061
rect 498055 376027 498071 376061
rect 498071 376027 498089 376061
rect 498127 376027 498139 376061
rect 498139 376027 498161 376061
rect 498199 376027 498207 376061
rect 498207 376027 498233 376061
rect 498271 376027 498275 376061
rect 498275 376027 498305 376061
rect 498343 376027 498377 376061
rect 497119 375569 497153 375603
rect 497191 375569 497221 375603
rect 497221 375569 497225 375603
rect 497263 375569 497289 375603
rect 497289 375569 497297 375603
rect 497335 375569 497357 375603
rect 497357 375569 497369 375603
rect 497407 375569 497425 375603
rect 497425 375569 497441 375603
rect 497479 375569 497493 375603
rect 497493 375569 497513 375603
rect 497551 375569 497561 375603
rect 497561 375569 497585 375603
rect 497623 375569 497629 375603
rect 497629 375569 497657 375603
rect 497695 375569 497697 375603
rect 497697 375569 497729 375603
rect 497767 375569 497799 375603
rect 497799 375569 497801 375603
rect 497839 375569 497867 375603
rect 497867 375569 497873 375603
rect 497911 375569 497935 375603
rect 497935 375569 497945 375603
rect 497983 375569 498003 375603
rect 498003 375569 498017 375603
rect 498055 375569 498071 375603
rect 498071 375569 498089 375603
rect 498127 375569 498139 375603
rect 498139 375569 498161 375603
rect 498199 375569 498207 375603
rect 498207 375569 498233 375603
rect 498271 375569 498275 375603
rect 498275 375569 498305 375603
rect 498343 375569 498377 375603
rect 496851 375307 496885 375341
rect 496851 374907 496885 374941
rect 496851 374507 496885 374541
rect 497119 375111 497153 375145
rect 497191 375111 497221 375145
rect 497221 375111 497225 375145
rect 497263 375111 497289 375145
rect 497289 375111 497297 375145
rect 497335 375111 497357 375145
rect 497357 375111 497369 375145
rect 497407 375111 497425 375145
rect 497425 375111 497441 375145
rect 497479 375111 497493 375145
rect 497493 375111 497513 375145
rect 497551 375111 497561 375145
rect 497561 375111 497585 375145
rect 497623 375111 497629 375145
rect 497629 375111 497657 375145
rect 497695 375111 497697 375145
rect 497697 375111 497729 375145
rect 497767 375111 497799 375145
rect 497799 375111 497801 375145
rect 497839 375111 497867 375145
rect 497867 375111 497873 375145
rect 497911 375111 497935 375145
rect 497935 375111 497945 375145
rect 497983 375111 498003 375145
rect 498003 375111 498017 375145
rect 498055 375111 498071 375145
rect 498071 375111 498089 375145
rect 498127 375111 498139 375145
rect 498139 375111 498161 375145
rect 498199 375111 498207 375145
rect 498207 375111 498233 375145
rect 498271 375111 498275 375145
rect 498275 375111 498305 375145
rect 498343 375111 498377 375145
rect 497119 374653 497153 374687
rect 497191 374653 497221 374687
rect 497221 374653 497225 374687
rect 497263 374653 497289 374687
rect 497289 374653 497297 374687
rect 497335 374653 497357 374687
rect 497357 374653 497369 374687
rect 497407 374653 497425 374687
rect 497425 374653 497441 374687
rect 497479 374653 497493 374687
rect 497493 374653 497513 374687
rect 497551 374653 497561 374687
rect 497561 374653 497585 374687
rect 497623 374653 497629 374687
rect 497629 374653 497657 374687
rect 497695 374653 497697 374687
rect 497697 374653 497729 374687
rect 497767 374653 497799 374687
rect 497799 374653 497801 374687
rect 497839 374653 497867 374687
rect 497867 374653 497873 374687
rect 497911 374653 497935 374687
rect 497935 374653 497945 374687
rect 497983 374653 498003 374687
rect 498003 374653 498017 374687
rect 498055 374653 498071 374687
rect 498071 374653 498089 374687
rect 498127 374653 498139 374687
rect 498139 374653 498161 374687
rect 498199 374653 498207 374687
rect 498207 374653 498233 374687
rect 498271 374653 498275 374687
rect 498275 374653 498305 374687
rect 498343 374653 498377 374687
rect 496851 374107 496885 374141
rect 496851 373707 496885 373741
rect 496851 373307 496885 373341
rect 496851 372907 496885 372941
rect 496851 372507 496885 372541
rect 497119 374195 497153 374229
rect 497191 374195 497221 374229
rect 497221 374195 497225 374229
rect 497263 374195 497289 374229
rect 497289 374195 497297 374229
rect 497335 374195 497357 374229
rect 497357 374195 497369 374229
rect 497407 374195 497425 374229
rect 497425 374195 497441 374229
rect 497479 374195 497493 374229
rect 497493 374195 497513 374229
rect 497551 374195 497561 374229
rect 497561 374195 497585 374229
rect 497623 374195 497629 374229
rect 497629 374195 497657 374229
rect 497695 374195 497697 374229
rect 497697 374195 497729 374229
rect 497767 374195 497799 374229
rect 497799 374195 497801 374229
rect 497839 374195 497867 374229
rect 497867 374195 497873 374229
rect 497911 374195 497935 374229
rect 497935 374195 497945 374229
rect 497983 374195 498003 374229
rect 498003 374195 498017 374229
rect 498055 374195 498071 374229
rect 498071 374195 498089 374229
rect 498127 374195 498139 374229
rect 498139 374195 498161 374229
rect 498199 374195 498207 374229
rect 498207 374195 498233 374229
rect 498271 374195 498275 374229
rect 498275 374195 498305 374229
rect 498343 374195 498377 374229
rect 497119 373737 497153 373771
rect 497191 373737 497221 373771
rect 497221 373737 497225 373771
rect 497263 373737 497289 373771
rect 497289 373737 497297 373771
rect 497335 373737 497357 373771
rect 497357 373737 497369 373771
rect 497407 373737 497425 373771
rect 497425 373737 497441 373771
rect 497479 373737 497493 373771
rect 497493 373737 497513 373771
rect 497551 373737 497561 373771
rect 497561 373737 497585 373771
rect 497623 373737 497629 373771
rect 497629 373737 497657 373771
rect 497695 373737 497697 373771
rect 497697 373737 497729 373771
rect 497767 373737 497799 373771
rect 497799 373737 497801 373771
rect 497839 373737 497867 373771
rect 497867 373737 497873 373771
rect 497911 373737 497935 373771
rect 497935 373737 497945 373771
rect 497983 373737 498003 373771
rect 498003 373737 498017 373771
rect 498055 373737 498071 373771
rect 498071 373737 498089 373771
rect 498127 373737 498139 373771
rect 498139 373737 498161 373771
rect 498199 373737 498207 373771
rect 498207 373737 498233 373771
rect 498271 373737 498275 373771
rect 498275 373737 498305 373771
rect 498343 373737 498377 373771
rect 497119 373279 497153 373313
rect 497191 373279 497221 373313
rect 497221 373279 497225 373313
rect 497263 373279 497289 373313
rect 497289 373279 497297 373313
rect 497335 373279 497357 373313
rect 497357 373279 497369 373313
rect 497407 373279 497425 373313
rect 497425 373279 497441 373313
rect 497479 373279 497493 373313
rect 497493 373279 497513 373313
rect 497551 373279 497561 373313
rect 497561 373279 497585 373313
rect 497623 373279 497629 373313
rect 497629 373279 497657 373313
rect 497695 373279 497697 373313
rect 497697 373279 497729 373313
rect 497767 373279 497799 373313
rect 497799 373279 497801 373313
rect 497839 373279 497867 373313
rect 497867 373279 497873 373313
rect 497911 373279 497935 373313
rect 497935 373279 497945 373313
rect 497983 373279 498003 373313
rect 498003 373279 498017 373313
rect 498055 373279 498071 373313
rect 498071 373279 498089 373313
rect 498127 373279 498139 373313
rect 498139 373279 498161 373313
rect 498199 373279 498207 373313
rect 498207 373279 498233 373313
rect 498271 373279 498275 373313
rect 498275 373279 498305 373313
rect 498343 373279 498377 373313
rect 497119 372821 497153 372855
rect 497191 372821 497221 372855
rect 497221 372821 497225 372855
rect 497263 372821 497289 372855
rect 497289 372821 497297 372855
rect 497335 372821 497357 372855
rect 497357 372821 497369 372855
rect 497407 372821 497425 372855
rect 497425 372821 497441 372855
rect 497479 372821 497493 372855
rect 497493 372821 497513 372855
rect 497551 372821 497561 372855
rect 497561 372821 497585 372855
rect 497623 372821 497629 372855
rect 497629 372821 497657 372855
rect 497695 372821 497697 372855
rect 497697 372821 497729 372855
rect 497767 372821 497799 372855
rect 497799 372821 497801 372855
rect 497839 372821 497867 372855
rect 497867 372821 497873 372855
rect 497911 372821 497935 372855
rect 497935 372821 497945 372855
rect 497983 372821 498003 372855
rect 498003 372821 498017 372855
rect 498055 372821 498071 372855
rect 498071 372821 498089 372855
rect 498127 372821 498139 372855
rect 498139 372821 498161 372855
rect 498199 372821 498207 372855
rect 498207 372821 498233 372855
rect 498271 372821 498275 372855
rect 498275 372821 498305 372855
rect 498343 372821 498377 372855
rect 497119 372363 497153 372397
rect 497191 372363 497221 372397
rect 497221 372363 497225 372397
rect 497263 372363 497289 372397
rect 497289 372363 497297 372397
rect 497335 372363 497357 372397
rect 497357 372363 497369 372397
rect 497407 372363 497425 372397
rect 497425 372363 497441 372397
rect 497479 372363 497493 372397
rect 497493 372363 497513 372397
rect 497551 372363 497561 372397
rect 497561 372363 497585 372397
rect 497623 372363 497629 372397
rect 497629 372363 497657 372397
rect 497695 372363 497697 372397
rect 497697 372363 497729 372397
rect 497767 372363 497799 372397
rect 497799 372363 497801 372397
rect 497839 372363 497867 372397
rect 497867 372363 497873 372397
rect 497911 372363 497935 372397
rect 497935 372363 497945 372397
rect 497983 372363 498003 372397
rect 498003 372363 498017 372397
rect 498055 372363 498071 372397
rect 498071 372363 498089 372397
rect 498127 372363 498139 372397
rect 498139 372363 498161 372397
rect 498199 372363 498207 372397
rect 498207 372363 498233 372397
rect 498271 372363 498275 372397
rect 498275 372363 498305 372397
rect 498343 372363 498377 372397
rect 498591 385451 498625 385485
rect 504371 399859 504405 399893
rect 498731 399707 498765 399741
rect 498731 399307 498765 399341
rect 498731 398907 498765 398941
rect 498731 398507 498765 398541
rect 498731 398107 498765 398141
rect 498731 397707 498765 397741
rect 498731 397307 498765 397341
rect 498731 396907 498765 396941
rect 498731 396507 498765 396541
rect 498731 396107 498765 396141
rect 498731 395707 498765 395741
rect 498731 395307 498765 395341
rect 498731 394907 498765 394941
rect 498731 394507 498765 394541
rect 498731 394107 498765 394141
rect 498731 393707 498765 393741
rect 498731 393307 498765 393341
rect 498731 392907 498765 392941
rect 500611 399607 500645 399641
rect 500611 399207 500645 399241
rect 500611 398807 500645 398841
rect 500611 398407 500645 398441
rect 500611 398007 500645 398041
rect 500611 397607 500645 397641
rect 500611 397207 500645 397241
rect 500611 396807 500645 396841
rect 500611 396407 500645 396441
rect 500611 396007 500645 396041
rect 500611 395607 500645 395641
rect 500611 395207 500645 395241
rect 500611 394807 500645 394841
rect 500611 394407 500645 394441
rect 500611 394007 500645 394041
rect 500611 393607 500645 393641
rect 500611 393207 500645 393241
rect 500611 392807 500645 392841
rect 502491 399607 502525 399641
rect 502491 399207 502525 399241
rect 502491 398807 502525 398841
rect 506251 400259 506285 400293
rect 506251 400059 506285 400093
rect 506251 399859 506285 399893
rect 504371 399659 504405 399693
rect 504371 399459 504405 399493
rect 504371 399259 504405 399293
rect 506251 399659 506285 399693
rect 506251 399459 506285 399493
rect 504371 399059 504405 399093
rect 504639 398856 505177 399250
rect 505599 398856 506137 399250
rect 506251 399259 506285 399293
rect 506251 399059 506285 399093
rect 502491 398407 502525 398441
rect 502491 398007 502525 398041
rect 502491 397607 502525 397641
rect 502491 397207 502525 397241
rect 502491 396807 502525 396841
rect 502491 396407 502525 396441
rect 504371 398315 504405 398349
rect 504371 398115 504405 398149
rect 504639 398119 505177 398513
rect 505599 398119 506137 398513
rect 506251 398315 506285 398349
rect 506251 398115 506285 398149
rect 504371 397915 504405 397949
rect 504371 397715 504405 397749
rect 506251 397915 506285 397949
rect 506251 397715 506285 397749
rect 504371 397515 504405 397549
rect 504371 397315 504405 397349
rect 504371 397115 504405 397149
rect 506251 397515 506285 397549
rect 506251 397315 506285 397349
rect 506251 397115 506285 397149
rect 504371 396915 504405 396949
rect 504371 396715 504405 396749
rect 504371 396515 504405 396549
rect 506251 396915 506285 396949
rect 506251 396715 506285 396749
rect 504371 396315 504405 396349
rect 504639 396112 505177 396506
rect 505599 396112 506137 396506
rect 506251 396515 506285 396549
rect 506251 396315 506285 396349
rect 511891 398217 511925 398251
rect 511891 398017 511925 398051
rect 512159 398021 512697 398415
rect 513119 398021 513657 398415
rect 513771 398217 513805 398251
rect 513771 398017 513805 398051
rect 511891 397817 511925 397851
rect 511891 397617 511925 397651
rect 513771 397817 513805 397851
rect 513771 397617 513805 397651
rect 511891 397417 511925 397451
rect 511891 397217 511925 397251
rect 511891 397017 511925 397051
rect 513771 397417 513805 397451
rect 513771 397217 513805 397251
rect 513771 397017 513805 397051
rect 511891 396817 511925 396851
rect 511891 396617 511925 396651
rect 511891 396417 511925 396451
rect 513771 396817 513805 396851
rect 513771 396617 513805 396651
rect 511891 396217 511925 396251
rect 502491 396007 502525 396041
rect 512159 396014 512697 396408
rect 513119 396014 513657 396408
rect 513771 396417 513805 396451
rect 513771 396217 513805 396251
rect 502491 395607 502525 395641
rect 502491 395207 502525 395241
rect 502491 394807 502525 394841
rect 502491 394407 502525 394441
rect 502491 394007 502525 394041
rect 502491 393607 502525 393641
rect 502491 393207 502525 393241
rect 502491 392807 502525 392841
rect 504371 395569 504405 395603
rect 504371 395369 504405 395403
rect 504639 395374 505177 395768
rect 505599 395374 506137 395768
rect 506251 395569 506285 395603
rect 506251 395369 506285 395403
rect 504371 395169 504405 395203
rect 504371 394969 504405 395003
rect 504371 394769 504405 394803
rect 504371 394569 504405 394603
rect 506251 395169 506285 395203
rect 506251 394969 506285 395003
rect 506251 394769 506285 394803
rect 504371 394369 504405 394403
rect 504371 394169 504405 394203
rect 504371 393969 504405 394003
rect 506251 394569 506285 394603
rect 506251 394369 506285 394403
rect 506251 394169 506285 394203
rect 504371 393769 504405 393803
rect 504371 393569 504405 393603
rect 504371 393369 504405 393403
rect 506251 393969 506285 394003
rect 506251 393769 506285 393803
rect 506251 393569 506285 393603
rect 506251 393369 506285 393403
rect 504371 393169 504405 393203
rect 504371 392969 504405 393003
rect 504639 392793 505177 393187
rect 505599 392793 506137 393187
rect 508131 395473 508165 395507
rect 508131 395273 508165 395307
rect 508399 395277 508937 395671
rect 509359 395277 509897 395671
rect 510011 395473 510045 395507
rect 510011 395273 510045 395307
rect 508131 395073 508165 395107
rect 508131 394873 508165 394907
rect 510011 395073 510045 395107
rect 510011 394873 510045 394907
rect 508131 394673 508165 394707
rect 508131 394473 508165 394507
rect 508131 394273 508165 394307
rect 510011 394673 510045 394707
rect 510011 394473 510045 394507
rect 510011 394273 510045 394307
rect 508131 394073 508165 394107
rect 508131 393873 508165 393907
rect 508131 393673 508165 393707
rect 510011 394073 510045 394107
rect 510011 393873 510045 393907
rect 508131 393473 508165 393507
rect 508399 393270 508937 393664
rect 509359 393270 509897 393664
rect 510011 393673 510045 393707
rect 510011 393473 510045 393507
rect 511891 395473 511925 395507
rect 511891 395273 511925 395307
rect 512159 395277 512697 395671
rect 513119 395277 513657 395671
rect 513771 395473 513805 395507
rect 513771 395273 513805 395307
rect 511891 395073 511925 395107
rect 511891 394873 511925 394907
rect 513771 395073 513805 395107
rect 513771 394873 513805 394907
rect 511891 394673 511925 394707
rect 511891 394473 511925 394507
rect 511891 394273 511925 394307
rect 513771 394673 513805 394707
rect 513771 394473 513805 394507
rect 513771 394273 513805 394307
rect 511891 394073 511925 394107
rect 511891 393873 511925 393907
rect 511891 393673 511925 393707
rect 513771 394073 513805 394107
rect 513771 393873 513805 393907
rect 511891 393473 511925 393507
rect 512159 393270 512697 393664
rect 513119 393270 513657 393664
rect 513771 393673 513805 393707
rect 513771 393473 513805 393507
rect 506251 393169 506285 393203
rect 506251 392969 506285 393003
rect 508131 392727 508165 392761
rect 498731 392507 498765 392541
rect 508131 392527 508165 392561
rect 498731 392107 498765 392141
rect 498731 391707 498765 391741
rect 498731 391307 498765 391341
rect 498731 390907 498765 390941
rect 498731 390507 498765 390541
rect 498731 390107 498765 390141
rect 498731 389707 498765 389741
rect 498731 389307 498765 389341
rect 498731 388907 498765 388941
rect 498731 388507 498765 388541
rect 498731 388107 498765 388141
rect 498731 387707 498765 387741
rect 498731 387307 498765 387341
rect 498731 386907 498765 386941
rect 500611 392063 500645 392097
rect 500611 391663 500645 391697
rect 500879 392199 500913 392233
rect 500951 392199 500981 392233
rect 500981 392199 500985 392233
rect 501023 392199 501049 392233
rect 501049 392199 501057 392233
rect 501095 392199 501117 392233
rect 501117 392199 501129 392233
rect 501167 392199 501185 392233
rect 501185 392199 501201 392233
rect 501239 392199 501253 392233
rect 501253 392199 501273 392233
rect 501311 392199 501321 392233
rect 501321 392199 501345 392233
rect 501383 392199 501389 392233
rect 501389 392199 501417 392233
rect 501455 392199 501457 392233
rect 501457 392199 501489 392233
rect 501527 392199 501559 392233
rect 501559 392199 501561 392233
rect 501599 392199 501627 392233
rect 501627 392199 501633 392233
rect 501671 392199 501695 392233
rect 501695 392199 501705 392233
rect 501743 392199 501763 392233
rect 501763 392199 501777 392233
rect 501815 392199 501831 392233
rect 501831 392199 501849 392233
rect 501887 392199 501899 392233
rect 501899 392199 501921 392233
rect 501959 392199 501967 392233
rect 501967 392199 501993 392233
rect 502031 392199 502035 392233
rect 502035 392199 502065 392233
rect 502103 392199 502137 392233
rect 502229 392167 502263 392201
rect 500879 391741 500913 391775
rect 500951 391741 500981 391775
rect 500981 391741 500985 391775
rect 501023 391741 501049 391775
rect 501049 391741 501057 391775
rect 501095 391741 501117 391775
rect 501117 391741 501129 391775
rect 501167 391741 501185 391775
rect 501185 391741 501201 391775
rect 501239 391741 501253 391775
rect 501253 391741 501273 391775
rect 501311 391741 501321 391775
rect 501321 391741 501345 391775
rect 501383 391741 501389 391775
rect 501389 391741 501417 391775
rect 501455 391741 501457 391775
rect 501457 391741 501489 391775
rect 501527 391741 501559 391775
rect 501559 391741 501561 391775
rect 501599 391741 501627 391775
rect 501627 391741 501633 391775
rect 501671 391741 501695 391775
rect 501695 391741 501705 391775
rect 501743 391741 501763 391775
rect 501763 391741 501777 391775
rect 501815 391741 501831 391775
rect 501831 391741 501849 391775
rect 501887 391741 501899 391775
rect 501899 391741 501921 391775
rect 501959 391741 501967 391775
rect 501967 391741 501993 391775
rect 502031 391741 502035 391775
rect 502035 391741 502065 391775
rect 502103 391741 502137 391775
rect 500611 391263 500645 391297
rect 500611 390863 500645 390897
rect 500611 390463 500645 390497
rect 500611 390063 500645 390097
rect 500879 391283 500913 391317
rect 500951 391283 500981 391317
rect 500981 391283 500985 391317
rect 501023 391283 501049 391317
rect 501049 391283 501057 391317
rect 501095 391283 501117 391317
rect 501117 391283 501129 391317
rect 501167 391283 501185 391317
rect 501185 391283 501201 391317
rect 501239 391283 501253 391317
rect 501253 391283 501273 391317
rect 501311 391283 501321 391317
rect 501321 391283 501345 391317
rect 501383 391283 501389 391317
rect 501389 391283 501417 391317
rect 501455 391283 501457 391317
rect 501457 391283 501489 391317
rect 501527 391283 501559 391317
rect 501559 391283 501561 391317
rect 501599 391283 501627 391317
rect 501627 391283 501633 391317
rect 501671 391283 501695 391317
rect 501695 391283 501705 391317
rect 501743 391283 501763 391317
rect 501763 391283 501777 391317
rect 501815 391283 501831 391317
rect 501831 391283 501849 391317
rect 501887 391283 501899 391317
rect 501899 391283 501921 391317
rect 501959 391283 501967 391317
rect 501967 391283 501993 391317
rect 502031 391283 502035 391317
rect 502035 391283 502065 391317
rect 502103 391283 502137 391317
rect 500879 390825 500913 390859
rect 500951 390825 500981 390859
rect 500981 390825 500985 390859
rect 501023 390825 501049 390859
rect 501049 390825 501057 390859
rect 501095 390825 501117 390859
rect 501117 390825 501129 390859
rect 501167 390825 501185 390859
rect 501185 390825 501201 390859
rect 501239 390825 501253 390859
rect 501253 390825 501273 390859
rect 501311 390825 501321 390859
rect 501321 390825 501345 390859
rect 501383 390825 501389 390859
rect 501389 390825 501417 390859
rect 501455 390825 501457 390859
rect 501457 390825 501489 390859
rect 501527 390825 501559 390859
rect 501559 390825 501561 390859
rect 501599 390825 501627 390859
rect 501627 390825 501633 390859
rect 501671 390825 501695 390859
rect 501695 390825 501705 390859
rect 501743 390825 501763 390859
rect 501763 390825 501777 390859
rect 501815 390825 501831 390859
rect 501831 390825 501849 390859
rect 501887 390825 501899 390859
rect 501899 390825 501921 390859
rect 501959 390825 501967 390859
rect 501967 390825 501993 390859
rect 502031 390825 502035 390859
rect 502035 390825 502065 390859
rect 502103 390825 502137 390859
rect 500879 390367 500913 390401
rect 500951 390367 500981 390401
rect 500981 390367 500985 390401
rect 501023 390367 501049 390401
rect 501049 390367 501057 390401
rect 501095 390367 501117 390401
rect 501117 390367 501129 390401
rect 501167 390367 501185 390401
rect 501185 390367 501201 390401
rect 501239 390367 501253 390401
rect 501253 390367 501273 390401
rect 501311 390367 501321 390401
rect 501321 390367 501345 390401
rect 501383 390367 501389 390401
rect 501389 390367 501417 390401
rect 501455 390367 501457 390401
rect 501457 390367 501489 390401
rect 501527 390367 501559 390401
rect 501559 390367 501561 390401
rect 501599 390367 501627 390401
rect 501627 390367 501633 390401
rect 501671 390367 501695 390401
rect 501695 390367 501705 390401
rect 501743 390367 501763 390401
rect 501763 390367 501777 390401
rect 501815 390367 501831 390401
rect 501831 390367 501849 390401
rect 501887 390367 501899 390401
rect 501899 390367 501921 390401
rect 501959 390367 501967 390401
rect 501967 390367 501993 390401
rect 502031 390367 502035 390401
rect 502035 390367 502065 390401
rect 502103 390367 502137 390401
rect 500801 390051 500835 390085
rect 500879 389909 500913 389943
rect 500951 389909 500981 389943
rect 500981 389909 500985 389943
rect 501023 389909 501049 389943
rect 501049 389909 501057 389943
rect 501095 389909 501117 389943
rect 501117 389909 501129 389943
rect 501167 389909 501185 389943
rect 501185 389909 501201 389943
rect 501239 389909 501253 389943
rect 501253 389909 501273 389943
rect 501311 389909 501321 389943
rect 501321 389909 501345 389943
rect 501383 389909 501389 389943
rect 501389 389909 501417 389943
rect 501455 389909 501457 389943
rect 501457 389909 501489 389943
rect 501527 389909 501559 389943
rect 501559 389909 501561 389943
rect 501599 389909 501627 389943
rect 501627 389909 501633 389943
rect 501671 389909 501695 389943
rect 501695 389909 501705 389943
rect 501743 389909 501763 389943
rect 501763 389909 501777 389943
rect 501815 389909 501831 389943
rect 501831 389909 501849 389943
rect 501887 389909 501899 389943
rect 501899 389909 501921 389943
rect 501959 389909 501967 389943
rect 501967 389909 501993 389943
rect 502031 389909 502035 389943
rect 502035 389909 502065 389943
rect 502103 389909 502137 389943
rect 500611 389663 500645 389697
rect 500611 389263 500645 389297
rect 500611 388863 500645 388897
rect 500879 389451 500913 389485
rect 500951 389451 500981 389485
rect 500981 389451 500985 389485
rect 501023 389451 501049 389485
rect 501049 389451 501057 389485
rect 501095 389451 501117 389485
rect 501117 389451 501129 389485
rect 501167 389451 501185 389485
rect 501185 389451 501201 389485
rect 501239 389451 501253 389485
rect 501253 389451 501273 389485
rect 501311 389451 501321 389485
rect 501321 389451 501345 389485
rect 501383 389451 501389 389485
rect 501389 389451 501417 389485
rect 501455 389451 501457 389485
rect 501457 389451 501489 389485
rect 501527 389451 501559 389485
rect 501559 389451 501561 389485
rect 501599 389451 501627 389485
rect 501627 389451 501633 389485
rect 501671 389451 501695 389485
rect 501695 389451 501705 389485
rect 501743 389451 501763 389485
rect 501763 389451 501777 389485
rect 501815 389451 501831 389485
rect 501831 389451 501849 389485
rect 501887 389451 501899 389485
rect 501899 389451 501921 389485
rect 501959 389451 501967 389485
rect 501967 389451 501993 389485
rect 502031 389451 502035 389485
rect 502035 389451 502065 389485
rect 502103 389451 502137 389485
rect 500879 388993 500913 389027
rect 500951 388993 500981 389027
rect 500981 388993 500985 389027
rect 501023 388993 501049 389027
rect 501049 388993 501057 389027
rect 501095 388993 501117 389027
rect 501117 388993 501129 389027
rect 501167 388993 501185 389027
rect 501185 388993 501201 389027
rect 501239 388993 501253 389027
rect 501253 388993 501273 389027
rect 501311 388993 501321 389027
rect 501321 388993 501345 389027
rect 501383 388993 501389 389027
rect 501389 388993 501417 389027
rect 501455 388993 501457 389027
rect 501457 388993 501489 389027
rect 501527 388993 501559 389027
rect 501559 388993 501561 389027
rect 501599 388993 501627 389027
rect 501627 388993 501633 389027
rect 501671 388993 501695 389027
rect 501695 388993 501705 389027
rect 501743 388993 501763 389027
rect 501763 388993 501777 389027
rect 501815 388993 501831 389027
rect 501831 388993 501849 389027
rect 501887 388993 501899 389027
rect 501899 388993 501921 389027
rect 501959 388993 501967 389027
rect 501967 388993 501993 389027
rect 502031 388993 502035 389027
rect 502035 388993 502065 389027
rect 502103 388993 502137 389027
rect 500611 388463 500645 388497
rect 500611 388063 500645 388097
rect 500611 387663 500645 387697
rect 500611 387263 500645 387297
rect 500611 386863 500645 386897
rect 500879 388535 500913 388569
rect 500951 388535 500981 388569
rect 500981 388535 500985 388569
rect 501023 388535 501049 388569
rect 501049 388535 501057 388569
rect 501095 388535 501117 388569
rect 501117 388535 501129 388569
rect 501167 388535 501185 388569
rect 501185 388535 501201 388569
rect 501239 388535 501253 388569
rect 501253 388535 501273 388569
rect 501311 388535 501321 388569
rect 501321 388535 501345 388569
rect 501383 388535 501389 388569
rect 501389 388535 501417 388569
rect 501455 388535 501457 388569
rect 501457 388535 501489 388569
rect 501527 388535 501559 388569
rect 501559 388535 501561 388569
rect 501599 388535 501627 388569
rect 501627 388535 501633 388569
rect 501671 388535 501695 388569
rect 501695 388535 501705 388569
rect 501743 388535 501763 388569
rect 501763 388535 501777 388569
rect 501815 388535 501831 388569
rect 501831 388535 501849 388569
rect 501887 388535 501899 388569
rect 501899 388535 501921 388569
rect 501959 388535 501967 388569
rect 501967 388535 501993 388569
rect 502031 388535 502035 388569
rect 502035 388535 502065 388569
rect 502103 388535 502137 388569
rect 500879 388077 500913 388111
rect 500951 388077 500981 388111
rect 500981 388077 500985 388111
rect 501023 388077 501049 388111
rect 501049 388077 501057 388111
rect 501095 388077 501117 388111
rect 501117 388077 501129 388111
rect 501167 388077 501185 388111
rect 501185 388077 501201 388111
rect 501239 388077 501253 388111
rect 501253 388077 501273 388111
rect 501311 388077 501321 388111
rect 501321 388077 501345 388111
rect 501383 388077 501389 388111
rect 501389 388077 501417 388111
rect 501455 388077 501457 388111
rect 501457 388077 501489 388111
rect 501527 388077 501559 388111
rect 501559 388077 501561 388111
rect 501599 388077 501627 388111
rect 501627 388077 501633 388111
rect 501671 388077 501695 388111
rect 501695 388077 501705 388111
rect 501743 388077 501763 388111
rect 501763 388077 501777 388111
rect 501815 388077 501831 388111
rect 501831 388077 501849 388111
rect 501887 388077 501899 388111
rect 501899 388077 501921 388111
rect 501959 388077 501967 388111
rect 501967 388077 501993 388111
rect 502031 388077 502035 388111
rect 502035 388077 502065 388111
rect 502103 388077 502137 388111
rect 500879 387619 500913 387653
rect 500951 387619 500981 387653
rect 500981 387619 500985 387653
rect 501023 387619 501049 387653
rect 501049 387619 501057 387653
rect 501095 387619 501117 387653
rect 501117 387619 501129 387653
rect 501167 387619 501185 387653
rect 501185 387619 501201 387653
rect 501239 387619 501253 387653
rect 501253 387619 501273 387653
rect 501311 387619 501321 387653
rect 501321 387619 501345 387653
rect 501383 387619 501389 387653
rect 501389 387619 501417 387653
rect 501455 387619 501457 387653
rect 501457 387619 501489 387653
rect 501527 387619 501559 387653
rect 501559 387619 501561 387653
rect 501599 387619 501627 387653
rect 501627 387619 501633 387653
rect 501671 387619 501695 387653
rect 501695 387619 501705 387653
rect 501743 387619 501763 387653
rect 501763 387619 501777 387653
rect 501815 387619 501831 387653
rect 501831 387619 501849 387653
rect 501887 387619 501899 387653
rect 501899 387619 501921 387653
rect 501959 387619 501967 387653
rect 501967 387619 501993 387653
rect 502031 387619 502035 387653
rect 502035 387619 502065 387653
rect 502103 387619 502137 387653
rect 500879 387161 500913 387195
rect 500951 387161 500981 387195
rect 500981 387161 500985 387195
rect 501023 387161 501049 387195
rect 501049 387161 501057 387195
rect 501095 387161 501117 387195
rect 501117 387161 501129 387195
rect 501167 387161 501185 387195
rect 501185 387161 501201 387195
rect 501239 387161 501253 387195
rect 501253 387161 501273 387195
rect 501311 387161 501321 387195
rect 501321 387161 501345 387195
rect 501383 387161 501389 387195
rect 501389 387161 501417 387195
rect 501455 387161 501457 387195
rect 501457 387161 501489 387195
rect 501527 387161 501559 387195
rect 501559 387161 501561 387195
rect 501599 387161 501627 387195
rect 501627 387161 501633 387195
rect 501671 387161 501695 387195
rect 501695 387161 501705 387195
rect 501743 387161 501763 387195
rect 501763 387161 501777 387195
rect 501815 387161 501831 387195
rect 501831 387161 501849 387195
rect 501887 387161 501899 387195
rect 501899 387161 501921 387195
rect 501959 387161 501967 387195
rect 501967 387161 501993 387195
rect 502031 387161 502035 387195
rect 502035 387161 502065 387195
rect 502103 387161 502137 387195
rect 502229 386831 502263 386865
rect 500879 386703 500913 386737
rect 500951 386703 500981 386737
rect 500981 386703 500985 386737
rect 501023 386703 501049 386737
rect 501049 386703 501057 386737
rect 501095 386703 501117 386737
rect 501117 386703 501129 386737
rect 501167 386703 501185 386737
rect 501185 386703 501201 386737
rect 501239 386703 501253 386737
rect 501253 386703 501273 386737
rect 501311 386703 501321 386737
rect 501321 386703 501345 386737
rect 501383 386703 501389 386737
rect 501389 386703 501417 386737
rect 501455 386703 501457 386737
rect 501457 386703 501489 386737
rect 501527 386703 501559 386737
rect 501559 386703 501561 386737
rect 501599 386703 501627 386737
rect 501627 386703 501633 386737
rect 501671 386703 501695 386737
rect 501695 386703 501705 386737
rect 501743 386703 501763 386737
rect 501763 386703 501777 386737
rect 501815 386703 501831 386737
rect 501831 386703 501849 386737
rect 501887 386703 501899 386737
rect 501899 386703 501921 386737
rect 501959 386703 501967 386737
rect 501967 386703 501993 386737
rect 502031 386703 502035 386737
rect 502035 386703 502065 386737
rect 502103 386703 502137 386737
rect 502365 386647 502399 386681
rect 502491 392063 502525 392097
rect 502491 391663 502525 391697
rect 502491 391263 502525 391297
rect 502491 390863 502525 390897
rect 502491 390463 502525 390497
rect 502491 390063 502525 390097
rect 504371 392239 504405 392273
rect 504371 392039 504405 392073
rect 504639 392043 505177 392437
rect 505599 392043 506137 392437
rect 506251 392239 506285 392273
rect 506251 392039 506285 392073
rect 504371 391839 504405 391873
rect 504371 391639 504405 391673
rect 506251 391839 506285 391873
rect 506251 391639 506285 391673
rect 504371 391439 504405 391473
rect 504371 391239 504405 391273
rect 504371 391039 504405 391073
rect 506251 391439 506285 391473
rect 506251 391239 506285 391273
rect 506251 391039 506285 391073
rect 504371 390839 504405 390873
rect 504371 390639 504405 390673
rect 504371 390439 504405 390473
rect 506251 390839 506285 390873
rect 506251 390639 506285 390673
rect 504371 390239 504405 390273
rect 504639 390036 505177 390430
rect 505599 390036 506137 390430
rect 506251 390439 506285 390473
rect 506251 390239 506285 390273
rect 508399 392532 508937 392926
rect 509359 392532 509897 392926
rect 510011 392727 510045 392761
rect 510011 392527 510045 392561
rect 508131 392327 508165 392361
rect 508131 392127 508165 392161
rect 508131 391927 508165 391961
rect 508131 391727 508165 391761
rect 510011 392327 510045 392361
rect 510011 392127 510045 392161
rect 510011 391927 510045 391961
rect 508131 391527 508165 391561
rect 508131 391327 508165 391361
rect 508131 391127 508165 391161
rect 510011 391727 510045 391761
rect 510011 391527 510045 391561
rect 510011 391327 510045 391361
rect 508131 390927 508165 390961
rect 508131 390727 508165 390761
rect 508131 390527 508165 390561
rect 510011 391127 510045 391161
rect 510011 390927 510045 390961
rect 510011 390727 510045 390761
rect 510011 390527 510045 390561
rect 508131 390327 508165 390361
rect 508131 390127 508165 390161
rect 508399 389951 508937 390345
rect 509359 389951 509897 390345
rect 511891 392729 511925 392763
rect 511891 392529 511925 392563
rect 512159 392533 512697 392927
rect 513119 392533 513657 392927
rect 513771 392729 513805 392763
rect 513771 392529 513805 392563
rect 511891 392329 511925 392363
rect 511891 392129 511925 392163
rect 513771 392329 513805 392363
rect 513771 392129 513805 392163
rect 511891 391929 511925 391963
rect 511891 391729 511925 391763
rect 511891 391529 511925 391563
rect 513771 391929 513805 391963
rect 513771 391729 513805 391763
rect 513771 391529 513805 391563
rect 511891 391329 511925 391363
rect 511891 391129 511925 391163
rect 511891 390929 511925 390963
rect 513771 391329 513805 391363
rect 513771 391129 513805 391163
rect 511891 390729 511925 390763
rect 512159 390526 512697 390920
rect 513119 390526 513657 390920
rect 513771 390929 513805 390963
rect 513771 390729 513805 390763
rect 515651 392337 515685 392371
rect 515651 392137 515685 392171
rect 515919 392141 516457 392535
rect 516879 392141 517417 392535
rect 517531 392337 517565 392371
rect 517531 392137 517565 392171
rect 515651 391937 515685 391971
rect 515651 391737 515685 391771
rect 517531 391937 517565 391971
rect 517531 391737 517565 391771
rect 515651 391537 515685 391571
rect 515651 391337 515685 391371
rect 515651 391137 515685 391171
rect 517531 391537 517565 391571
rect 517531 391337 517565 391371
rect 517531 391137 517565 391171
rect 515651 390937 515685 390971
rect 515651 390737 515685 390771
rect 515651 390537 515685 390571
rect 517531 390937 517565 390971
rect 517531 390737 517565 390771
rect 510011 390327 510045 390361
rect 510011 390127 510045 390161
rect 515651 390337 515685 390371
rect 515919 390134 516457 390528
rect 516879 390134 517417 390528
rect 517531 390537 517565 390571
rect 517531 390337 517565 390371
rect 519411 390867 519445 390901
rect 519411 390667 519445 390701
rect 519679 390671 520217 391065
rect 520639 390671 521177 391065
rect 521291 390867 521325 390901
rect 521291 390667 521325 390701
rect 519411 390467 519445 390501
rect 519411 390267 519445 390301
rect 521291 390467 521325 390501
rect 521291 390267 521325 390301
rect 519411 390067 519445 390101
rect 502491 389663 502525 389697
rect 519411 389867 519445 389901
rect 519411 389667 519445 389701
rect 502491 389263 502525 389297
rect 502491 388863 502525 388897
rect 502491 388463 502525 388497
rect 502491 388063 502525 388097
rect 502491 387663 502525 387697
rect 502491 387263 502525 387297
rect 502491 386863 502525 386897
rect 504371 389319 504405 389353
rect 504371 388919 504405 388953
rect 504371 388519 504405 388553
rect 504371 388119 504405 388153
rect 504371 387719 504405 387753
rect 504371 387319 504405 387353
rect 504371 386919 504405 386953
rect 498731 386507 498765 386541
rect 498731 386107 498765 386141
rect 498731 385707 498765 385741
rect 504371 386519 504405 386553
rect 504371 386119 504405 386153
rect 504371 385719 504405 385753
rect 498731 385307 498765 385341
rect 498731 384907 498765 384941
rect 498731 384507 498765 384541
rect 498731 384107 498765 384141
rect 498731 383707 498765 383741
rect 498731 383307 498765 383341
rect 498731 382907 498765 382941
rect 498731 382507 498765 382541
rect 498731 382107 498765 382141
rect 498731 381707 498765 381741
rect 498731 381307 498765 381341
rect 498731 380907 498765 380941
rect 498731 380507 498765 380541
rect 498731 380107 498765 380141
rect 500611 385399 500645 385433
rect 500611 384999 500645 385033
rect 500879 385535 500913 385569
rect 500951 385535 500981 385569
rect 500981 385535 500985 385569
rect 501023 385535 501049 385569
rect 501049 385535 501057 385569
rect 501095 385535 501117 385569
rect 501117 385535 501129 385569
rect 501167 385535 501185 385569
rect 501185 385535 501201 385569
rect 501239 385535 501253 385569
rect 501253 385535 501273 385569
rect 501311 385535 501321 385569
rect 501321 385535 501345 385569
rect 501383 385535 501389 385569
rect 501389 385535 501417 385569
rect 501455 385535 501457 385569
rect 501457 385535 501489 385569
rect 501527 385535 501559 385569
rect 501559 385535 501561 385569
rect 501599 385535 501627 385569
rect 501627 385535 501633 385569
rect 501671 385535 501695 385569
rect 501695 385535 501705 385569
rect 501743 385535 501763 385569
rect 501763 385535 501777 385569
rect 501815 385535 501831 385569
rect 501831 385535 501849 385569
rect 501887 385535 501899 385569
rect 501899 385535 501921 385569
rect 501959 385535 501967 385569
rect 501967 385535 501993 385569
rect 502031 385535 502035 385569
rect 502035 385535 502065 385569
rect 502103 385535 502137 385569
rect 500879 385077 500913 385111
rect 500951 385077 500981 385111
rect 500981 385077 500985 385111
rect 501023 385077 501049 385111
rect 501049 385077 501057 385111
rect 501095 385077 501117 385111
rect 501117 385077 501129 385111
rect 501167 385077 501185 385111
rect 501185 385077 501201 385111
rect 501239 385077 501253 385111
rect 501253 385077 501273 385111
rect 501311 385077 501321 385111
rect 501321 385077 501345 385111
rect 501383 385077 501389 385111
rect 501389 385077 501417 385111
rect 501455 385077 501457 385111
rect 501457 385077 501489 385111
rect 501527 385077 501559 385111
rect 501559 385077 501561 385111
rect 501599 385077 501627 385111
rect 501627 385077 501633 385111
rect 501671 385077 501695 385111
rect 501695 385077 501705 385111
rect 501743 385077 501763 385111
rect 501763 385077 501777 385111
rect 501815 385077 501831 385111
rect 501831 385077 501849 385111
rect 501887 385077 501899 385111
rect 501899 385077 501921 385111
rect 501959 385077 501967 385111
rect 501967 385077 501993 385111
rect 502031 385077 502035 385111
rect 502035 385077 502065 385111
rect 502103 385077 502137 385111
rect 500611 384599 500645 384633
rect 500611 384199 500645 384233
rect 500611 383799 500645 383833
rect 500611 383399 500645 383433
rect 500879 384619 500913 384653
rect 500951 384619 500981 384653
rect 500981 384619 500985 384653
rect 501023 384619 501049 384653
rect 501049 384619 501057 384653
rect 501095 384619 501117 384653
rect 501117 384619 501129 384653
rect 501167 384619 501185 384653
rect 501185 384619 501201 384653
rect 501239 384619 501253 384653
rect 501253 384619 501273 384653
rect 501311 384619 501321 384653
rect 501321 384619 501345 384653
rect 501383 384619 501389 384653
rect 501389 384619 501417 384653
rect 501455 384619 501457 384653
rect 501457 384619 501489 384653
rect 501527 384619 501559 384653
rect 501559 384619 501561 384653
rect 501599 384619 501627 384653
rect 501627 384619 501633 384653
rect 501671 384619 501695 384653
rect 501695 384619 501705 384653
rect 501743 384619 501763 384653
rect 501763 384619 501777 384653
rect 501815 384619 501831 384653
rect 501831 384619 501849 384653
rect 501887 384619 501899 384653
rect 501899 384619 501921 384653
rect 501959 384619 501967 384653
rect 501967 384619 501993 384653
rect 502031 384619 502035 384653
rect 502035 384619 502065 384653
rect 502103 384619 502137 384653
rect 500879 384161 500913 384195
rect 500951 384161 500981 384195
rect 500981 384161 500985 384195
rect 501023 384161 501049 384195
rect 501049 384161 501057 384195
rect 501095 384161 501117 384195
rect 501117 384161 501129 384195
rect 501167 384161 501185 384195
rect 501185 384161 501201 384195
rect 501239 384161 501253 384195
rect 501253 384161 501273 384195
rect 501311 384161 501321 384195
rect 501321 384161 501345 384195
rect 501383 384161 501389 384195
rect 501389 384161 501417 384195
rect 501455 384161 501457 384195
rect 501457 384161 501489 384195
rect 501527 384161 501559 384195
rect 501559 384161 501561 384195
rect 501599 384161 501627 384195
rect 501627 384161 501633 384195
rect 501671 384161 501695 384195
rect 501695 384161 501705 384195
rect 501743 384161 501763 384195
rect 501763 384161 501777 384195
rect 501815 384161 501831 384195
rect 501831 384161 501849 384195
rect 501887 384161 501899 384195
rect 501899 384161 501921 384195
rect 501959 384161 501967 384195
rect 501967 384161 501993 384195
rect 502031 384161 502035 384195
rect 502035 384161 502065 384195
rect 502103 384161 502137 384195
rect 500879 383703 500913 383737
rect 500951 383703 500981 383737
rect 500981 383703 500985 383737
rect 501023 383703 501049 383737
rect 501049 383703 501057 383737
rect 501095 383703 501117 383737
rect 501117 383703 501129 383737
rect 501167 383703 501185 383737
rect 501185 383703 501201 383737
rect 501239 383703 501253 383737
rect 501253 383703 501273 383737
rect 501311 383703 501321 383737
rect 501321 383703 501345 383737
rect 501383 383703 501389 383737
rect 501389 383703 501417 383737
rect 501455 383703 501457 383737
rect 501457 383703 501489 383737
rect 501527 383703 501559 383737
rect 501559 383703 501561 383737
rect 501599 383703 501627 383737
rect 501627 383703 501633 383737
rect 501671 383703 501695 383737
rect 501695 383703 501705 383737
rect 501743 383703 501763 383737
rect 501763 383703 501777 383737
rect 501815 383703 501831 383737
rect 501831 383703 501849 383737
rect 501887 383703 501899 383737
rect 501899 383703 501921 383737
rect 501959 383703 501967 383737
rect 501967 383703 501993 383737
rect 502031 383703 502035 383737
rect 502035 383703 502065 383737
rect 502103 383703 502137 383737
rect 500879 383245 500913 383279
rect 500951 383245 500981 383279
rect 500981 383245 500985 383279
rect 501023 383245 501049 383279
rect 501049 383245 501057 383279
rect 501095 383245 501117 383279
rect 501117 383245 501129 383279
rect 501167 383245 501185 383279
rect 501185 383245 501201 383279
rect 501239 383245 501253 383279
rect 501253 383245 501273 383279
rect 501311 383245 501321 383279
rect 501321 383245 501345 383279
rect 501383 383245 501389 383279
rect 501389 383245 501417 383279
rect 501455 383245 501457 383279
rect 501457 383245 501489 383279
rect 501527 383245 501559 383279
rect 501559 383245 501561 383279
rect 501599 383245 501627 383279
rect 501627 383245 501633 383279
rect 501671 383245 501695 383279
rect 501695 383245 501705 383279
rect 501743 383245 501763 383279
rect 501763 383245 501777 383279
rect 501815 383245 501831 383279
rect 501831 383245 501849 383279
rect 501887 383245 501899 383279
rect 501899 383245 501921 383279
rect 501959 383245 501967 383279
rect 501967 383245 501993 383279
rect 502031 383245 502035 383279
rect 502035 383245 502065 383279
rect 502103 383245 502137 383279
rect 500611 382999 500645 383033
rect 500611 382599 500645 382633
rect 500611 382199 500645 382233
rect 500879 382787 500913 382821
rect 500951 382787 500981 382821
rect 500981 382787 500985 382821
rect 501023 382787 501049 382821
rect 501049 382787 501057 382821
rect 501095 382787 501117 382821
rect 501117 382787 501129 382821
rect 501167 382787 501185 382821
rect 501185 382787 501201 382821
rect 501239 382787 501253 382821
rect 501253 382787 501273 382821
rect 501311 382787 501321 382821
rect 501321 382787 501345 382821
rect 501383 382787 501389 382821
rect 501389 382787 501417 382821
rect 501455 382787 501457 382821
rect 501457 382787 501489 382821
rect 501527 382787 501559 382821
rect 501559 382787 501561 382821
rect 501599 382787 501627 382821
rect 501627 382787 501633 382821
rect 501671 382787 501695 382821
rect 501695 382787 501705 382821
rect 501743 382787 501763 382821
rect 501763 382787 501777 382821
rect 501815 382787 501831 382821
rect 501831 382787 501849 382821
rect 501887 382787 501899 382821
rect 501899 382787 501921 382821
rect 501959 382787 501967 382821
rect 501967 382787 501993 382821
rect 502031 382787 502035 382821
rect 502035 382787 502065 382821
rect 502103 382787 502137 382821
rect 500879 382329 500913 382363
rect 500951 382329 500981 382363
rect 500981 382329 500985 382363
rect 501023 382329 501049 382363
rect 501049 382329 501057 382363
rect 501095 382329 501117 382363
rect 501117 382329 501129 382363
rect 501167 382329 501185 382363
rect 501185 382329 501201 382363
rect 501239 382329 501253 382363
rect 501253 382329 501273 382363
rect 501311 382329 501321 382363
rect 501321 382329 501345 382363
rect 501383 382329 501389 382363
rect 501389 382329 501417 382363
rect 501455 382329 501457 382363
rect 501457 382329 501489 382363
rect 501527 382329 501559 382363
rect 501559 382329 501561 382363
rect 501599 382329 501627 382363
rect 501627 382329 501633 382363
rect 501671 382329 501695 382363
rect 501695 382329 501705 382363
rect 501743 382329 501763 382363
rect 501763 382329 501777 382363
rect 501815 382329 501831 382363
rect 501831 382329 501849 382363
rect 501887 382329 501899 382363
rect 501899 382329 501921 382363
rect 501959 382329 501967 382363
rect 501967 382329 501993 382363
rect 502031 382329 502035 382363
rect 502035 382329 502065 382363
rect 502103 382329 502137 382363
rect 500611 381799 500645 381833
rect 500611 381399 500645 381433
rect 500611 380999 500645 381033
rect 500611 380599 500645 380633
rect 500611 380199 500645 380233
rect 500879 381871 500913 381905
rect 500951 381871 500981 381905
rect 500981 381871 500985 381905
rect 501023 381871 501049 381905
rect 501049 381871 501057 381905
rect 501095 381871 501117 381905
rect 501117 381871 501129 381905
rect 501167 381871 501185 381905
rect 501185 381871 501201 381905
rect 501239 381871 501253 381905
rect 501253 381871 501273 381905
rect 501311 381871 501321 381905
rect 501321 381871 501345 381905
rect 501383 381871 501389 381905
rect 501389 381871 501417 381905
rect 501455 381871 501457 381905
rect 501457 381871 501489 381905
rect 501527 381871 501559 381905
rect 501559 381871 501561 381905
rect 501599 381871 501627 381905
rect 501627 381871 501633 381905
rect 501671 381871 501695 381905
rect 501695 381871 501705 381905
rect 501743 381871 501763 381905
rect 501763 381871 501777 381905
rect 501815 381871 501831 381905
rect 501831 381871 501849 381905
rect 501887 381871 501899 381905
rect 501899 381871 501921 381905
rect 501959 381871 501967 381905
rect 501967 381871 501993 381905
rect 502031 381871 502035 381905
rect 502035 381871 502065 381905
rect 502103 381871 502137 381905
rect 500879 381413 500913 381447
rect 500951 381413 500981 381447
rect 500981 381413 500985 381447
rect 501023 381413 501049 381447
rect 501049 381413 501057 381447
rect 501095 381413 501117 381447
rect 501117 381413 501129 381447
rect 501167 381413 501185 381447
rect 501185 381413 501201 381447
rect 501239 381413 501253 381447
rect 501253 381413 501273 381447
rect 501311 381413 501321 381447
rect 501321 381413 501345 381447
rect 501383 381413 501389 381447
rect 501389 381413 501417 381447
rect 501455 381413 501457 381447
rect 501457 381413 501489 381447
rect 501527 381413 501559 381447
rect 501559 381413 501561 381447
rect 501599 381413 501627 381447
rect 501627 381413 501633 381447
rect 501671 381413 501695 381447
rect 501695 381413 501705 381447
rect 501743 381413 501763 381447
rect 501763 381413 501777 381447
rect 501815 381413 501831 381447
rect 501831 381413 501849 381447
rect 501887 381413 501899 381447
rect 501899 381413 501921 381447
rect 501959 381413 501967 381447
rect 501967 381413 501993 381447
rect 502031 381413 502035 381447
rect 502035 381413 502065 381447
rect 502103 381413 502137 381447
rect 500879 380955 500913 380989
rect 500951 380955 500981 380989
rect 500981 380955 500985 380989
rect 501023 380955 501049 380989
rect 501049 380955 501057 380989
rect 501095 380955 501117 380989
rect 501117 380955 501129 380989
rect 501167 380955 501185 380989
rect 501185 380955 501201 380989
rect 501239 380955 501253 380989
rect 501253 380955 501273 380989
rect 501311 380955 501321 380989
rect 501321 380955 501345 380989
rect 501383 380955 501389 380989
rect 501389 380955 501417 380989
rect 501455 380955 501457 380989
rect 501457 380955 501489 380989
rect 501527 380955 501559 380989
rect 501559 380955 501561 380989
rect 501599 380955 501627 380989
rect 501627 380955 501633 380989
rect 501671 380955 501695 380989
rect 501695 380955 501705 380989
rect 501743 380955 501763 380989
rect 501763 380955 501777 380989
rect 501815 380955 501831 380989
rect 501831 380955 501849 380989
rect 501887 380955 501899 380989
rect 501899 380955 501921 380989
rect 501959 380955 501967 380989
rect 501967 380955 501993 380989
rect 502031 380955 502035 380989
rect 502035 380955 502065 380989
rect 502103 380955 502137 380989
rect 500879 380497 500913 380531
rect 500951 380497 500981 380531
rect 500981 380497 500985 380531
rect 501023 380497 501049 380531
rect 501049 380497 501057 380531
rect 501095 380497 501117 380531
rect 501117 380497 501129 380531
rect 501167 380497 501185 380531
rect 501185 380497 501201 380531
rect 501239 380497 501253 380531
rect 501253 380497 501273 380531
rect 501311 380497 501321 380531
rect 501321 380497 501345 380531
rect 501383 380497 501389 380531
rect 501389 380497 501417 380531
rect 501455 380497 501457 380531
rect 501457 380497 501489 380531
rect 501527 380497 501559 380531
rect 501559 380497 501561 380531
rect 501599 380497 501627 380531
rect 501627 380497 501633 380531
rect 501671 380497 501695 380531
rect 501695 380497 501705 380531
rect 501743 380497 501763 380531
rect 501763 380497 501777 380531
rect 501815 380497 501831 380531
rect 501831 380497 501849 380531
rect 501887 380497 501899 380531
rect 501899 380497 501921 380531
rect 501959 380497 501967 380531
rect 501967 380497 501993 380531
rect 502031 380497 502035 380531
rect 502035 380497 502065 380531
rect 502103 380497 502137 380531
rect 500879 380039 500913 380073
rect 500951 380039 500981 380073
rect 500981 380039 500985 380073
rect 501023 380039 501049 380073
rect 501049 380039 501057 380073
rect 501095 380039 501117 380073
rect 501117 380039 501129 380073
rect 501167 380039 501185 380073
rect 501185 380039 501201 380073
rect 501239 380039 501253 380073
rect 501253 380039 501273 380073
rect 501311 380039 501321 380073
rect 501321 380039 501345 380073
rect 501383 380039 501389 380073
rect 501389 380039 501417 380073
rect 501455 380039 501457 380073
rect 501457 380039 501489 380073
rect 501527 380039 501559 380073
rect 501559 380039 501561 380073
rect 501599 380039 501627 380073
rect 501627 380039 501633 380073
rect 501671 380039 501695 380073
rect 501695 380039 501705 380073
rect 501743 380039 501763 380073
rect 501763 380039 501777 380073
rect 501815 380039 501831 380073
rect 501831 380039 501849 380073
rect 501887 380039 501899 380073
rect 501899 380039 501921 380073
rect 501959 380039 501967 380073
rect 501967 380039 501993 380073
rect 502031 380039 502035 380073
rect 502035 380039 502065 380073
rect 502103 380039 502137 380073
rect 502365 385451 502399 385485
rect 502491 385399 502525 385433
rect 504891 389490 504911 389524
rect 504911 389490 504925 389524
rect 504963 389490 504979 389524
rect 504979 389490 504997 389524
rect 505035 389490 505047 389524
rect 505047 389490 505069 389524
rect 505107 389490 505115 389524
rect 505115 389490 505141 389524
rect 505179 389490 505183 389524
rect 505183 389490 505213 389524
rect 505251 389490 505285 389524
rect 505323 389490 505353 389524
rect 505353 389490 505357 389524
rect 505395 389490 505421 389524
rect 505421 389490 505429 389524
rect 505467 389490 505489 389524
rect 505489 389490 505501 389524
rect 505539 389490 505557 389524
rect 505557 389490 505573 389524
rect 505611 389490 505625 389524
rect 505625 389490 505645 389524
rect 504891 389032 504911 389066
rect 504911 389032 504925 389066
rect 504963 389032 504979 389066
rect 504979 389032 504997 389066
rect 505035 389032 505047 389066
rect 505047 389032 505069 389066
rect 505107 389032 505115 389066
rect 505115 389032 505141 389066
rect 505179 389032 505183 389066
rect 505183 389032 505213 389066
rect 505251 389032 505285 389066
rect 505323 389032 505353 389066
rect 505353 389032 505357 389066
rect 505395 389032 505421 389066
rect 505421 389032 505429 389066
rect 505467 389032 505489 389066
rect 505489 389032 505501 389066
rect 505539 389032 505557 389066
rect 505557 389032 505573 389066
rect 505611 389032 505625 389066
rect 505625 389032 505645 389066
rect 504891 388574 504911 388608
rect 504911 388574 504925 388608
rect 504963 388574 504979 388608
rect 504979 388574 504997 388608
rect 505035 388574 505047 388608
rect 505047 388574 505069 388608
rect 505107 388574 505115 388608
rect 505115 388574 505141 388608
rect 505179 388574 505183 388608
rect 505183 388574 505213 388608
rect 505251 388574 505285 388608
rect 505323 388574 505353 388608
rect 505353 388574 505357 388608
rect 505395 388574 505421 388608
rect 505421 388574 505429 388608
rect 505467 388574 505489 388608
rect 505489 388574 505501 388608
rect 505539 388574 505557 388608
rect 505557 388574 505573 388608
rect 505611 388574 505625 388608
rect 505625 388574 505645 388608
rect 504891 388116 504911 388150
rect 504911 388116 504925 388150
rect 504963 388116 504979 388150
rect 504979 388116 504997 388150
rect 505035 388116 505047 388150
rect 505047 388116 505069 388150
rect 505107 388116 505115 388150
rect 505115 388116 505141 388150
rect 505179 388116 505183 388150
rect 505183 388116 505213 388150
rect 505251 388116 505285 388150
rect 505323 388116 505353 388150
rect 505353 388116 505357 388150
rect 505395 388116 505421 388150
rect 505421 388116 505429 388150
rect 505467 388116 505489 388150
rect 505489 388116 505501 388150
rect 505539 388116 505557 388150
rect 505557 388116 505573 388150
rect 505611 388116 505625 388150
rect 505625 388116 505645 388150
rect 504891 387658 504911 387692
rect 504911 387658 504925 387692
rect 504963 387658 504979 387692
rect 504979 387658 504997 387692
rect 505035 387658 505047 387692
rect 505047 387658 505069 387692
rect 505107 387658 505115 387692
rect 505115 387658 505141 387692
rect 505179 387658 505183 387692
rect 505183 387658 505213 387692
rect 505251 387658 505285 387692
rect 505323 387658 505353 387692
rect 505353 387658 505357 387692
rect 505395 387658 505421 387692
rect 505421 387658 505429 387692
rect 505467 387658 505489 387692
rect 505489 387658 505501 387692
rect 505539 387658 505557 387692
rect 505557 387658 505573 387692
rect 505611 387658 505625 387692
rect 505625 387658 505645 387692
rect 504891 387200 504911 387234
rect 504911 387200 504925 387234
rect 504963 387200 504979 387234
rect 504979 387200 504997 387234
rect 505035 387200 505047 387234
rect 505047 387200 505069 387234
rect 505107 387200 505115 387234
rect 505115 387200 505141 387234
rect 505179 387200 505183 387234
rect 505183 387200 505213 387234
rect 505251 387200 505285 387234
rect 505323 387200 505353 387234
rect 505353 387200 505357 387234
rect 505395 387200 505421 387234
rect 505421 387200 505429 387234
rect 505467 387200 505489 387234
rect 505489 387200 505501 387234
rect 505539 387200 505557 387234
rect 505557 387200 505573 387234
rect 505611 387200 505625 387234
rect 505625 387200 505645 387234
rect 506251 389319 506285 389353
rect 506251 388919 506285 388953
rect 515651 389319 515685 389353
rect 515651 388919 515685 388953
rect 506251 388519 506285 388553
rect 506251 388119 506285 388153
rect 506251 387719 506285 387753
rect 506251 387319 506285 387353
rect 505901 386831 505935 386865
rect 504891 386742 504911 386776
rect 504911 386742 504925 386776
rect 504963 386742 504979 386776
rect 504979 386742 504997 386776
rect 505035 386742 505047 386776
rect 505047 386742 505069 386776
rect 505107 386742 505115 386776
rect 505115 386742 505141 386776
rect 505179 386742 505183 386776
rect 505183 386742 505213 386776
rect 505251 386742 505285 386776
rect 505323 386742 505353 386776
rect 505353 386742 505357 386776
rect 505395 386742 505421 386776
rect 505421 386742 505429 386776
rect 505467 386742 505489 386776
rect 505489 386742 505501 386776
rect 505539 386742 505557 386776
rect 505557 386742 505573 386776
rect 505611 386742 505625 386776
rect 505625 386742 505645 386776
rect 504891 386284 504911 386318
rect 504911 386284 504925 386318
rect 504963 386284 504979 386318
rect 504979 386284 504997 386318
rect 505035 386284 505047 386318
rect 505047 386284 505069 386318
rect 505107 386284 505115 386318
rect 505115 386284 505141 386318
rect 505179 386284 505183 386318
rect 505183 386284 505213 386318
rect 505251 386284 505285 386318
rect 505323 386284 505353 386318
rect 505353 386284 505357 386318
rect 505395 386284 505421 386318
rect 505421 386284 505429 386318
rect 505467 386284 505489 386318
rect 505489 386284 505501 386318
rect 505539 386284 505557 386318
rect 505557 386284 505573 386318
rect 505611 386284 505625 386318
rect 505625 386284 505645 386318
rect 504891 385826 504911 385860
rect 504911 385826 504925 385860
rect 504963 385826 504979 385860
rect 504979 385826 504997 385860
rect 505035 385826 505047 385860
rect 505047 385826 505069 385860
rect 505107 385826 505115 385860
rect 505115 385826 505141 385860
rect 505179 385826 505183 385860
rect 505183 385826 505213 385860
rect 505251 385826 505285 385860
rect 505323 385826 505353 385860
rect 505353 385826 505357 385860
rect 505395 385826 505421 385860
rect 505421 385826 505429 385860
rect 505467 385826 505489 385860
rect 505489 385826 505501 385860
rect 505539 385826 505557 385860
rect 505557 385826 505573 385860
rect 505611 385826 505625 385860
rect 505625 385826 505645 385860
rect 504891 385368 504911 385402
rect 504911 385368 504925 385402
rect 504963 385368 504979 385402
rect 504979 385368 504997 385402
rect 505035 385368 505047 385402
rect 505047 385368 505069 385402
rect 505107 385368 505115 385402
rect 505115 385368 505141 385402
rect 505179 385368 505183 385402
rect 505183 385368 505213 385402
rect 505251 385368 505285 385402
rect 505323 385368 505353 385402
rect 505353 385368 505357 385402
rect 505395 385368 505421 385402
rect 505421 385368 505429 385402
rect 505467 385368 505489 385402
rect 505489 385368 505501 385402
rect 505539 385368 505557 385402
rect 505557 385368 505573 385402
rect 505611 385368 505625 385402
rect 505625 385368 505645 385402
rect 506251 386919 506285 386953
rect 506251 386519 506285 386553
rect 506251 386119 506285 386153
rect 506251 385719 506285 385753
rect 508131 388533 508165 388567
rect 508131 388133 508165 388167
rect 508131 387733 508165 387767
rect 508131 387333 508165 387367
rect 508131 386933 508165 386967
rect 508131 386533 508165 386567
rect 508131 386133 508165 386167
rect 508131 385733 508165 385767
rect 502491 384999 502525 385033
rect 508131 385333 508165 385367
rect 502491 384599 502525 384633
rect 502491 384199 502525 384233
rect 502491 383799 502525 383833
rect 502491 383399 502525 383433
rect 502491 382999 502525 383033
rect 502491 382599 502525 382633
rect 502491 382199 502525 382233
rect 502491 381799 502525 381833
rect 502491 381399 502525 381433
rect 502491 380999 502525 381033
rect 502491 380599 502525 380633
rect 502491 380199 502525 380233
rect 504371 384809 504405 384843
rect 504371 384409 504405 384443
rect 504371 384009 504405 384043
rect 504371 383609 504405 383643
rect 504371 383209 504405 383243
rect 504371 382809 504405 382843
rect 504371 382409 504405 382443
rect 504371 382009 504405 382043
rect 504371 381609 504405 381643
rect 504371 381209 504405 381243
rect 504371 380809 504405 380843
rect 504371 380409 504405 380443
rect 504371 380009 504405 380043
rect 498731 379707 498765 379741
rect 498731 379307 498765 379341
rect 498731 378907 498765 378941
rect 498731 378507 498765 378541
rect 498731 378107 498765 378141
rect 504371 379609 504405 379643
rect 504371 379209 504405 379243
rect 504371 378809 504405 378843
rect 504371 378409 504405 378443
rect 504371 378009 504405 378043
rect 506251 384809 506285 384843
rect 506251 384409 506285 384443
rect 506251 384009 506285 384043
rect 506251 383609 506285 383643
rect 506251 383209 506285 383243
rect 506251 382809 506285 382843
rect 506251 382409 506285 382443
rect 506251 382009 506285 382043
rect 506251 381609 506285 381643
rect 508131 384933 508165 384967
rect 508131 384533 508165 384567
rect 508131 384133 508165 384167
rect 508131 383733 508165 383767
rect 508131 383333 508165 383367
rect 508131 382933 508165 382967
rect 508131 382533 508165 382567
rect 508131 382133 508165 382167
rect 508131 381733 508165 381767
rect 510011 388533 510045 388567
rect 510011 388133 510045 388167
rect 510011 387733 510045 387767
rect 515651 388519 515685 388553
rect 515651 388119 515685 388153
rect 510011 387333 510045 387367
rect 510011 386933 510045 386967
rect 510011 386533 510045 386567
rect 510011 386133 510045 386167
rect 510011 385733 510045 385767
rect 510011 385333 510045 385367
rect 511891 387535 511925 387569
rect 511891 387335 511925 387369
rect 512159 387339 512697 387733
rect 513119 387339 513657 387733
rect 513771 387535 513805 387569
rect 513771 387335 513805 387369
rect 511891 387135 511925 387169
rect 511891 386935 511925 386969
rect 513771 387135 513805 387169
rect 513771 386935 513805 386969
rect 511891 386735 511925 386769
rect 511891 386535 511925 386569
rect 511891 386335 511925 386369
rect 513771 386735 513805 386769
rect 513771 386535 513805 386569
rect 513771 386335 513805 386369
rect 511891 386135 511925 386169
rect 511891 385935 511925 385969
rect 511891 385735 511925 385769
rect 513771 386135 513805 386169
rect 513771 385935 513805 385969
rect 511891 385535 511925 385569
rect 512159 385332 512697 385726
rect 513119 385332 513657 385726
rect 513771 385735 513805 385769
rect 513771 385535 513805 385569
rect 515651 387719 515685 387753
rect 515651 387319 515685 387353
rect 515651 386919 515685 386953
rect 515651 386519 515685 386553
rect 515651 386119 515685 386153
rect 515651 385719 515685 385753
rect 516171 389490 516191 389524
rect 516191 389490 516205 389524
rect 516243 389490 516259 389524
rect 516259 389490 516277 389524
rect 516315 389490 516327 389524
rect 516327 389490 516349 389524
rect 516387 389490 516395 389524
rect 516395 389490 516421 389524
rect 516459 389490 516463 389524
rect 516463 389490 516493 389524
rect 516531 389490 516565 389524
rect 516603 389490 516633 389524
rect 516633 389490 516637 389524
rect 516675 389490 516701 389524
rect 516701 389490 516709 389524
rect 516747 389490 516769 389524
rect 516769 389490 516781 389524
rect 516819 389490 516837 389524
rect 516837 389490 516853 389524
rect 516891 389490 516905 389524
rect 516905 389490 516925 389524
rect 516171 389032 516191 389066
rect 516191 389032 516205 389066
rect 516243 389032 516259 389066
rect 516259 389032 516277 389066
rect 516315 389032 516327 389066
rect 516327 389032 516349 389066
rect 516387 389032 516395 389066
rect 516395 389032 516421 389066
rect 516459 389032 516463 389066
rect 516463 389032 516493 389066
rect 516531 389032 516565 389066
rect 516603 389032 516633 389066
rect 516633 389032 516637 389066
rect 516675 389032 516701 389066
rect 516701 389032 516709 389066
rect 516747 389032 516769 389066
rect 516769 389032 516781 389066
rect 516819 389032 516837 389066
rect 516837 389032 516853 389066
rect 516891 389032 516905 389066
rect 516905 389032 516925 389066
rect 516171 388574 516191 388608
rect 516191 388574 516205 388608
rect 516243 388574 516259 388608
rect 516259 388574 516277 388608
rect 516315 388574 516327 388608
rect 516327 388574 516349 388608
rect 516387 388574 516395 388608
rect 516395 388574 516421 388608
rect 516459 388574 516463 388608
rect 516463 388574 516493 388608
rect 516531 388574 516565 388608
rect 516603 388574 516633 388608
rect 516633 388574 516637 388608
rect 516675 388574 516701 388608
rect 516701 388574 516709 388608
rect 516747 388574 516769 388608
rect 516769 388574 516781 388608
rect 516819 388574 516837 388608
rect 516837 388574 516853 388608
rect 516891 388574 516905 388608
rect 516905 388574 516925 388608
rect 516171 388116 516191 388150
rect 516191 388116 516205 388150
rect 516243 388116 516259 388150
rect 516259 388116 516277 388150
rect 516315 388116 516327 388150
rect 516327 388116 516349 388150
rect 516387 388116 516395 388150
rect 516395 388116 516421 388150
rect 516459 388116 516463 388150
rect 516463 388116 516493 388150
rect 516531 388116 516565 388150
rect 516603 388116 516633 388150
rect 516633 388116 516637 388150
rect 516675 388116 516701 388150
rect 516701 388116 516709 388150
rect 516747 388116 516769 388150
rect 516769 388116 516781 388150
rect 516819 388116 516837 388150
rect 516837 388116 516853 388150
rect 516891 388116 516905 388150
rect 516905 388116 516925 388150
rect 516171 387658 516191 387692
rect 516191 387658 516205 387692
rect 516243 387658 516259 387692
rect 516259 387658 516277 387692
rect 516315 387658 516327 387692
rect 516327 387658 516349 387692
rect 516387 387658 516395 387692
rect 516395 387658 516421 387692
rect 516459 387658 516463 387692
rect 516463 387658 516493 387692
rect 516531 387658 516565 387692
rect 516603 387658 516633 387692
rect 516633 387658 516637 387692
rect 516675 387658 516701 387692
rect 516701 387658 516709 387692
rect 516747 387658 516769 387692
rect 516769 387658 516781 387692
rect 516819 387658 516837 387692
rect 516837 387658 516853 387692
rect 516891 387658 516905 387692
rect 516905 387658 516925 387692
rect 516171 387200 516191 387234
rect 516191 387200 516205 387234
rect 516243 387200 516259 387234
rect 516259 387200 516277 387234
rect 516315 387200 516327 387234
rect 516327 387200 516349 387234
rect 516387 387200 516395 387234
rect 516395 387200 516421 387234
rect 516459 387200 516463 387234
rect 516463 387200 516493 387234
rect 516531 387200 516565 387234
rect 516603 387200 516633 387234
rect 516633 387200 516637 387234
rect 516675 387200 516701 387234
rect 516701 387200 516709 387234
rect 516747 387200 516769 387234
rect 516769 387200 516781 387234
rect 516819 387200 516837 387234
rect 516837 387200 516853 387234
rect 516891 387200 516905 387234
rect 516905 387200 516925 387234
rect 516171 386742 516191 386776
rect 516191 386742 516205 386776
rect 516243 386742 516259 386776
rect 516259 386742 516277 386776
rect 516315 386742 516327 386776
rect 516327 386742 516349 386776
rect 516387 386742 516395 386776
rect 516395 386742 516421 386776
rect 516459 386742 516463 386776
rect 516463 386742 516493 386776
rect 516531 386742 516565 386776
rect 516603 386742 516633 386776
rect 516633 386742 516637 386776
rect 516675 386742 516701 386776
rect 516701 386742 516709 386776
rect 516747 386742 516769 386776
rect 516769 386742 516781 386776
rect 516819 386742 516837 386776
rect 516837 386742 516853 386776
rect 516891 386742 516905 386776
rect 516905 386742 516925 386776
rect 516171 386284 516191 386318
rect 516191 386284 516205 386318
rect 516243 386284 516259 386318
rect 516259 386284 516277 386318
rect 516315 386284 516327 386318
rect 516327 386284 516349 386318
rect 516387 386284 516395 386318
rect 516395 386284 516421 386318
rect 516459 386284 516463 386318
rect 516463 386284 516493 386318
rect 516531 386284 516565 386318
rect 516603 386284 516633 386318
rect 516633 386284 516637 386318
rect 516675 386284 516701 386318
rect 516701 386284 516709 386318
rect 516747 386284 516769 386318
rect 516769 386284 516781 386318
rect 516819 386284 516837 386318
rect 516837 386284 516853 386318
rect 516891 386284 516905 386318
rect 516905 386284 516925 386318
rect 516171 385826 516191 385860
rect 516191 385826 516205 385860
rect 516243 385826 516259 385860
rect 516259 385826 516277 385860
rect 516315 385826 516327 385860
rect 516327 385826 516349 385860
rect 516387 385826 516395 385860
rect 516395 385826 516421 385860
rect 516459 385826 516463 385860
rect 516463 385826 516493 385860
rect 516531 385826 516565 385860
rect 516603 385826 516633 385860
rect 516633 385826 516637 385860
rect 516675 385826 516701 385860
rect 516701 385826 516709 385860
rect 516747 385826 516769 385860
rect 516769 385826 516781 385860
rect 516819 385826 516837 385860
rect 516837 385826 516853 385860
rect 516891 385826 516905 385860
rect 516905 385826 516925 385860
rect 516171 385368 516191 385402
rect 516191 385368 516205 385402
rect 516243 385368 516259 385402
rect 516259 385368 516277 385402
rect 516315 385368 516327 385402
rect 516327 385368 516349 385402
rect 516387 385368 516395 385402
rect 516395 385368 516421 385402
rect 516459 385368 516463 385402
rect 516463 385368 516493 385402
rect 516531 385368 516565 385402
rect 516603 385368 516633 385402
rect 516633 385368 516637 385402
rect 516675 385368 516701 385402
rect 516701 385368 516709 385402
rect 516747 385368 516769 385402
rect 516769 385368 516781 385402
rect 516819 385368 516837 385402
rect 516837 385368 516853 385402
rect 516891 385368 516905 385402
rect 516905 385368 516925 385402
rect 517531 389319 517565 389353
rect 517531 388919 517565 388953
rect 521291 390067 521325 390101
rect 521291 389867 521325 389901
rect 521291 389667 521325 389701
rect 519411 389467 519445 389501
rect 519411 389267 519445 389301
rect 519411 389067 519445 389101
rect 521291 389467 521325 389501
rect 521291 389267 521325 389301
rect 519411 388867 519445 388901
rect 519679 388664 520217 389058
rect 520639 388664 521177 389058
rect 521291 389067 521325 389101
rect 521291 388867 521325 388901
rect 523171 389907 523205 389941
rect 523171 389507 523205 389541
rect 523439 390043 523473 390077
rect 523511 390043 523541 390077
rect 523541 390043 523545 390077
rect 523583 390043 523609 390077
rect 523609 390043 523617 390077
rect 523655 390043 523677 390077
rect 523677 390043 523689 390077
rect 523727 390043 523745 390077
rect 523745 390043 523761 390077
rect 523799 390043 523813 390077
rect 523813 390043 523833 390077
rect 523871 390043 523881 390077
rect 523881 390043 523905 390077
rect 523943 390043 523949 390077
rect 523949 390043 523977 390077
rect 524015 390043 524017 390077
rect 524017 390043 524049 390077
rect 524087 390043 524119 390077
rect 524119 390043 524121 390077
rect 524159 390043 524187 390077
rect 524187 390043 524193 390077
rect 524231 390043 524255 390077
rect 524255 390043 524265 390077
rect 524303 390043 524323 390077
rect 524323 390043 524337 390077
rect 524375 390043 524391 390077
rect 524391 390043 524409 390077
rect 524447 390043 524459 390077
rect 524459 390043 524481 390077
rect 524519 390043 524527 390077
rect 524527 390043 524553 390077
rect 524591 390043 524595 390077
rect 524595 390043 524625 390077
rect 524663 390043 524697 390077
rect 523439 389585 523473 389619
rect 523511 389585 523541 389619
rect 523541 389585 523545 389619
rect 523583 389585 523609 389619
rect 523609 389585 523617 389619
rect 523655 389585 523677 389619
rect 523677 389585 523689 389619
rect 523727 389585 523745 389619
rect 523745 389585 523761 389619
rect 523799 389585 523813 389619
rect 523813 389585 523833 389619
rect 523871 389585 523881 389619
rect 523881 389585 523905 389619
rect 523943 389585 523949 389619
rect 523949 389585 523977 389619
rect 524015 389585 524017 389619
rect 524017 389585 524049 389619
rect 524087 389585 524119 389619
rect 524119 389585 524121 389619
rect 524159 389585 524187 389619
rect 524187 389585 524193 389619
rect 524231 389585 524255 389619
rect 524255 389585 524265 389619
rect 524303 389585 524323 389619
rect 524323 389585 524337 389619
rect 524375 389585 524391 389619
rect 524391 389585 524409 389619
rect 524447 389585 524459 389619
rect 524459 389585 524481 389619
rect 524519 389585 524527 389619
rect 524527 389585 524553 389619
rect 524591 389585 524595 389619
rect 524595 389585 524625 389619
rect 524663 389585 524697 389619
rect 523171 389107 523205 389141
rect 523171 388707 523205 388741
rect 517531 388519 517565 388553
rect 517189 387383 517223 387417
rect 517531 388119 517565 388153
rect 517531 387719 517565 387753
rect 523171 388307 523205 388341
rect 523171 387907 523205 387941
rect 523439 389127 523473 389161
rect 523511 389127 523541 389161
rect 523541 389127 523545 389161
rect 523583 389127 523609 389161
rect 523609 389127 523617 389161
rect 523655 389127 523677 389161
rect 523677 389127 523689 389161
rect 523727 389127 523745 389161
rect 523745 389127 523761 389161
rect 523799 389127 523813 389161
rect 523813 389127 523833 389161
rect 523871 389127 523881 389161
rect 523881 389127 523905 389161
rect 523943 389127 523949 389161
rect 523949 389127 523977 389161
rect 524015 389127 524017 389161
rect 524017 389127 524049 389161
rect 524087 389127 524119 389161
rect 524119 389127 524121 389161
rect 524159 389127 524187 389161
rect 524187 389127 524193 389161
rect 524231 389127 524255 389161
rect 524255 389127 524265 389161
rect 524303 389127 524323 389161
rect 524323 389127 524337 389161
rect 524375 389127 524391 389161
rect 524391 389127 524409 389161
rect 524447 389127 524459 389161
rect 524459 389127 524481 389161
rect 524519 389127 524527 389161
rect 524527 389127 524553 389161
rect 524591 389127 524595 389161
rect 524595 389127 524625 389161
rect 524663 389127 524697 389161
rect 523439 388669 523473 388703
rect 523511 388669 523541 388703
rect 523541 388669 523545 388703
rect 523583 388669 523609 388703
rect 523609 388669 523617 388703
rect 523655 388669 523677 388703
rect 523677 388669 523689 388703
rect 523727 388669 523745 388703
rect 523745 388669 523761 388703
rect 523799 388669 523813 388703
rect 523813 388669 523833 388703
rect 523871 388669 523881 388703
rect 523881 388669 523905 388703
rect 523943 388669 523949 388703
rect 523949 388669 523977 388703
rect 524015 388669 524017 388703
rect 524017 388669 524049 388703
rect 524087 388669 524119 388703
rect 524119 388669 524121 388703
rect 524159 388669 524187 388703
rect 524187 388669 524193 388703
rect 524231 388669 524255 388703
rect 524255 388669 524265 388703
rect 524303 388669 524323 388703
rect 524323 388669 524337 388703
rect 524375 388669 524391 388703
rect 524391 388669 524409 388703
rect 524447 388669 524459 388703
rect 524459 388669 524481 388703
rect 524519 388669 524527 388703
rect 524527 388669 524553 388703
rect 524591 388669 524595 388703
rect 524595 388669 524625 388703
rect 524663 388669 524697 388703
rect 517531 387319 517565 387353
rect 517531 386919 517565 386953
rect 517531 386519 517565 386553
rect 517531 386119 517565 386153
rect 517531 385719 517565 385753
rect 519411 387535 519445 387569
rect 519411 387335 519445 387369
rect 519679 387339 520217 387733
rect 520639 387339 521177 387733
rect 521291 387535 521325 387569
rect 521291 387335 521325 387369
rect 519411 387135 519445 387169
rect 519411 386935 519445 386969
rect 521291 387135 521325 387169
rect 521291 386935 521325 386969
rect 519411 386735 519445 386769
rect 519411 386535 519445 386569
rect 519411 386335 519445 386369
rect 521291 386735 521325 386769
rect 521291 386535 521325 386569
rect 521291 386335 521325 386369
rect 519411 386135 519445 386169
rect 519411 385935 519445 385969
rect 519411 385735 519445 385769
rect 521291 386135 521325 386169
rect 521291 385935 521325 385969
rect 519411 385535 519445 385569
rect 519679 385332 520217 385726
rect 520639 385332 521177 385726
rect 521291 385735 521325 385769
rect 521291 385535 521325 385569
rect 523439 388211 523473 388245
rect 523511 388211 523541 388245
rect 523541 388211 523545 388245
rect 523583 388211 523609 388245
rect 523609 388211 523617 388245
rect 523655 388211 523677 388245
rect 523677 388211 523689 388245
rect 523727 388211 523745 388245
rect 523745 388211 523761 388245
rect 523799 388211 523813 388245
rect 523813 388211 523833 388245
rect 523871 388211 523881 388245
rect 523881 388211 523905 388245
rect 523943 388211 523949 388245
rect 523949 388211 523977 388245
rect 524015 388211 524017 388245
rect 524017 388211 524049 388245
rect 524087 388211 524119 388245
rect 524119 388211 524121 388245
rect 524159 388211 524187 388245
rect 524187 388211 524193 388245
rect 524231 388211 524255 388245
rect 524255 388211 524265 388245
rect 524303 388211 524323 388245
rect 524323 388211 524337 388245
rect 524375 388211 524391 388245
rect 524391 388211 524409 388245
rect 524447 388211 524459 388245
rect 524459 388211 524481 388245
rect 524519 388211 524527 388245
rect 524527 388211 524553 388245
rect 524591 388211 524595 388245
rect 524595 388211 524625 388245
rect 524663 388211 524697 388245
rect 523439 387753 523473 387787
rect 523511 387753 523541 387787
rect 523541 387753 523545 387787
rect 523583 387753 523609 387787
rect 523609 387753 523617 387787
rect 523655 387753 523677 387787
rect 523677 387753 523689 387787
rect 523727 387753 523745 387787
rect 523745 387753 523761 387787
rect 523799 387753 523813 387787
rect 523813 387753 523833 387787
rect 523871 387753 523881 387787
rect 523881 387753 523905 387787
rect 523943 387753 523949 387787
rect 523949 387753 523977 387787
rect 524015 387753 524017 387787
rect 524017 387753 524049 387787
rect 524087 387753 524119 387787
rect 524119 387753 524121 387787
rect 524159 387753 524187 387787
rect 524187 387753 524193 387787
rect 524231 387753 524255 387787
rect 524255 387753 524265 387787
rect 524303 387753 524323 387787
rect 524323 387753 524337 387787
rect 524375 387753 524391 387787
rect 524391 387753 524409 387787
rect 524447 387753 524459 387787
rect 524459 387753 524481 387787
rect 524519 387753 524527 387787
rect 524527 387753 524553 387787
rect 524591 387753 524595 387787
rect 524595 387753 524625 387787
rect 524663 387753 524697 387787
rect 523171 387507 523205 387541
rect 523171 387107 523205 387141
rect 523171 386707 523205 386741
rect 523439 387295 523473 387329
rect 523511 387295 523541 387329
rect 523541 387295 523545 387329
rect 523583 387295 523609 387329
rect 523609 387295 523617 387329
rect 523655 387295 523677 387329
rect 523677 387295 523689 387329
rect 523727 387295 523745 387329
rect 523745 387295 523761 387329
rect 523799 387295 523813 387329
rect 523813 387295 523833 387329
rect 523871 387295 523881 387329
rect 523881 387295 523905 387329
rect 523943 387295 523949 387329
rect 523949 387295 523977 387329
rect 524015 387295 524017 387329
rect 524017 387295 524049 387329
rect 524087 387295 524119 387329
rect 524119 387295 524121 387329
rect 524159 387295 524187 387329
rect 524187 387295 524193 387329
rect 524231 387295 524255 387329
rect 524255 387295 524265 387329
rect 524303 387295 524323 387329
rect 524323 387295 524337 387329
rect 524375 387295 524391 387329
rect 524391 387295 524409 387329
rect 524447 387295 524459 387329
rect 524459 387295 524481 387329
rect 524519 387295 524527 387329
rect 524527 387295 524553 387329
rect 524591 387295 524595 387329
rect 524595 387295 524625 387329
rect 524663 387295 524697 387329
rect 523439 386837 523473 386871
rect 523511 386837 523541 386871
rect 523541 386837 523545 386871
rect 523583 386837 523609 386871
rect 523609 386837 523617 386871
rect 523655 386837 523677 386871
rect 523677 386837 523689 386871
rect 523727 386837 523745 386871
rect 523745 386837 523761 386871
rect 523799 386837 523813 386871
rect 523813 386837 523833 386871
rect 523871 386837 523881 386871
rect 523881 386837 523905 386871
rect 523943 386837 523949 386871
rect 523949 386837 523977 386871
rect 524015 386837 524017 386871
rect 524017 386837 524049 386871
rect 524087 386837 524119 386871
rect 524119 386837 524121 386871
rect 524159 386837 524187 386871
rect 524187 386837 524193 386871
rect 524231 386837 524255 386871
rect 524255 386837 524265 386871
rect 524303 386837 524323 386871
rect 524323 386837 524337 386871
rect 524375 386837 524391 386871
rect 524391 386837 524409 386871
rect 524447 386837 524459 386871
rect 524459 386837 524481 386871
rect 524519 386837 524527 386871
rect 524527 386837 524553 386871
rect 524591 386837 524595 386871
rect 524595 386837 524625 386871
rect 524663 386837 524697 386871
rect 523171 386307 523205 386341
rect 523171 385907 523205 385941
rect 523171 385507 523205 385541
rect 523439 386379 523473 386413
rect 523511 386379 523541 386413
rect 523541 386379 523545 386413
rect 523583 386379 523609 386413
rect 523609 386379 523617 386413
rect 523655 386379 523677 386413
rect 523677 386379 523689 386413
rect 523727 386379 523745 386413
rect 523745 386379 523761 386413
rect 523799 386379 523813 386413
rect 523813 386379 523833 386413
rect 523871 386379 523881 386413
rect 523881 386379 523905 386413
rect 523943 386379 523949 386413
rect 523949 386379 523977 386413
rect 524015 386379 524017 386413
rect 524017 386379 524049 386413
rect 524087 386379 524119 386413
rect 524119 386379 524121 386413
rect 524159 386379 524187 386413
rect 524187 386379 524193 386413
rect 524231 386379 524255 386413
rect 524255 386379 524265 386413
rect 524303 386379 524323 386413
rect 524323 386379 524337 386413
rect 524375 386379 524391 386413
rect 524391 386379 524409 386413
rect 524447 386379 524459 386413
rect 524459 386379 524481 386413
rect 524519 386379 524527 386413
rect 524527 386379 524553 386413
rect 524591 386379 524595 386413
rect 524595 386379 524625 386413
rect 524663 386379 524697 386413
rect 523439 385921 523473 385955
rect 523511 385921 523541 385955
rect 523541 385921 523545 385955
rect 523583 385921 523609 385955
rect 523609 385921 523617 385955
rect 523655 385921 523677 385955
rect 523677 385921 523689 385955
rect 523727 385921 523745 385955
rect 523745 385921 523761 385955
rect 523799 385921 523813 385955
rect 523813 385921 523833 385955
rect 523871 385921 523881 385955
rect 523881 385921 523905 385955
rect 523943 385921 523949 385955
rect 523949 385921 523977 385955
rect 524015 385921 524017 385955
rect 524017 385921 524049 385955
rect 524087 385921 524119 385955
rect 524119 385921 524121 385955
rect 524159 385921 524187 385955
rect 524187 385921 524193 385955
rect 524231 385921 524255 385955
rect 524255 385921 524265 385955
rect 524303 385921 524323 385955
rect 524323 385921 524337 385955
rect 524375 385921 524391 385955
rect 524391 385921 524409 385955
rect 524447 385921 524459 385955
rect 524459 385921 524481 385955
rect 524519 385921 524527 385955
rect 524527 385921 524553 385955
rect 524591 385921 524595 385955
rect 524595 385921 524625 385955
rect 524663 385921 524697 385955
rect 523171 385107 523205 385141
rect 510011 384933 510045 384967
rect 510011 384533 510045 384567
rect 510011 384133 510045 384167
rect 510011 383733 510045 383767
rect 510011 383333 510045 383367
rect 510011 382933 510045 382967
rect 510011 382533 510045 382567
rect 510011 382133 510045 382167
rect 510011 381733 510045 381767
rect 511891 384809 511925 384843
rect 511891 384409 511925 384443
rect 511891 384009 511925 384043
rect 511891 383609 511925 383643
rect 511891 383209 511925 383243
rect 511891 382809 511925 382843
rect 511891 382409 511925 382443
rect 511891 382009 511925 382043
rect 511891 381609 511925 381643
rect 506251 381209 506285 381243
rect 506251 380809 506285 380843
rect 506251 380409 506285 380443
rect 506251 380009 506285 380043
rect 506251 379609 506285 379643
rect 506251 379209 506285 379243
rect 506251 378809 506285 378843
rect 506251 378409 506285 378443
rect 506251 378009 506285 378043
rect 508131 381085 508165 381119
rect 508131 380685 508165 380719
rect 508131 380285 508165 380319
rect 508131 379885 508165 379919
rect 508131 379485 508165 379519
rect 508131 379085 508165 379119
rect 508131 378685 508165 378719
rect 508131 378285 508165 378319
rect 508131 377885 508165 377919
rect 498731 377707 498765 377741
rect 498731 377307 498765 377341
rect 498731 376907 498765 376941
rect 498731 376507 498765 376541
rect 498731 376107 498765 376141
rect 498731 375707 498765 375741
rect 498731 375307 498765 375341
rect 498731 374907 498765 374941
rect 498731 374507 498765 374541
rect 498731 374107 498765 374141
rect 498731 373707 498765 373741
rect 500611 377461 500645 377495
rect 500611 377061 500645 377095
rect 500611 376661 500645 376695
rect 500611 376261 500645 376295
rect 500611 375861 500645 375895
rect 500611 375461 500645 375495
rect 500611 375061 500645 375095
rect 500611 374661 500645 374695
rect 500611 374261 500645 374295
rect 500611 373861 500645 373895
rect 501131 377632 501151 377666
rect 501151 377632 501165 377666
rect 501203 377632 501219 377666
rect 501219 377632 501237 377666
rect 501275 377632 501287 377666
rect 501287 377632 501309 377666
rect 501347 377632 501355 377666
rect 501355 377632 501381 377666
rect 501419 377632 501423 377666
rect 501423 377632 501453 377666
rect 501491 377632 501525 377666
rect 501563 377632 501593 377666
rect 501593 377632 501597 377666
rect 501635 377632 501661 377666
rect 501661 377632 501669 377666
rect 501707 377632 501729 377666
rect 501729 377632 501741 377666
rect 501779 377632 501797 377666
rect 501797 377632 501813 377666
rect 501851 377632 501865 377666
rect 501865 377632 501885 377666
rect 501131 377174 501151 377208
rect 501151 377174 501165 377208
rect 501203 377174 501219 377208
rect 501219 377174 501237 377208
rect 501275 377174 501287 377208
rect 501287 377174 501309 377208
rect 501347 377174 501355 377208
rect 501355 377174 501381 377208
rect 501419 377174 501423 377208
rect 501423 377174 501453 377208
rect 501491 377174 501525 377208
rect 501563 377174 501593 377208
rect 501593 377174 501597 377208
rect 501635 377174 501661 377208
rect 501661 377174 501669 377208
rect 501707 377174 501729 377208
rect 501729 377174 501741 377208
rect 501779 377174 501797 377208
rect 501797 377174 501813 377208
rect 501851 377174 501865 377208
rect 501865 377174 501885 377208
rect 501131 376716 501151 376750
rect 501151 376716 501165 376750
rect 501203 376716 501219 376750
rect 501219 376716 501237 376750
rect 501275 376716 501287 376750
rect 501287 376716 501309 376750
rect 501347 376716 501355 376750
rect 501355 376716 501381 376750
rect 501419 376716 501423 376750
rect 501423 376716 501453 376750
rect 501491 376716 501525 376750
rect 501563 376716 501593 376750
rect 501593 376716 501597 376750
rect 501635 376716 501661 376750
rect 501661 376716 501669 376750
rect 501707 376716 501729 376750
rect 501729 376716 501741 376750
rect 501779 376716 501797 376750
rect 501797 376716 501813 376750
rect 501851 376716 501865 376750
rect 501865 376716 501885 376750
rect 501131 376258 501151 376292
rect 501151 376258 501165 376292
rect 501203 376258 501219 376292
rect 501219 376258 501237 376292
rect 501275 376258 501287 376292
rect 501287 376258 501309 376292
rect 501347 376258 501355 376292
rect 501355 376258 501381 376292
rect 501419 376258 501423 376292
rect 501423 376258 501453 376292
rect 501491 376258 501525 376292
rect 501563 376258 501593 376292
rect 501593 376258 501597 376292
rect 501635 376258 501661 376292
rect 501661 376258 501669 376292
rect 501707 376258 501729 376292
rect 501729 376258 501741 376292
rect 501779 376258 501797 376292
rect 501797 376258 501813 376292
rect 501851 376258 501865 376292
rect 501865 376258 501885 376292
rect 501131 375800 501151 375834
rect 501151 375800 501165 375834
rect 501203 375800 501219 375834
rect 501219 375800 501237 375834
rect 501275 375800 501287 375834
rect 501287 375800 501309 375834
rect 501347 375800 501355 375834
rect 501355 375800 501381 375834
rect 501419 375800 501423 375834
rect 501423 375800 501453 375834
rect 501491 375800 501525 375834
rect 501563 375800 501593 375834
rect 501593 375800 501597 375834
rect 501635 375800 501661 375834
rect 501661 375800 501669 375834
rect 501707 375800 501729 375834
rect 501729 375800 501741 375834
rect 501779 375800 501797 375834
rect 501797 375800 501813 375834
rect 501851 375800 501865 375834
rect 501865 375800 501885 375834
rect 501131 375342 501151 375376
rect 501151 375342 501165 375376
rect 501203 375342 501219 375376
rect 501219 375342 501237 375376
rect 501275 375342 501287 375376
rect 501287 375342 501309 375376
rect 501347 375342 501355 375376
rect 501355 375342 501381 375376
rect 501419 375342 501423 375376
rect 501423 375342 501453 375376
rect 501491 375342 501525 375376
rect 501563 375342 501593 375376
rect 501593 375342 501597 375376
rect 501635 375342 501661 375376
rect 501661 375342 501669 375376
rect 501707 375342 501729 375376
rect 501729 375342 501741 375376
rect 501779 375342 501797 375376
rect 501797 375342 501813 375376
rect 501851 375342 501865 375376
rect 501865 375342 501885 375376
rect 501131 374884 501151 374918
rect 501151 374884 501165 374918
rect 501203 374884 501219 374918
rect 501219 374884 501237 374918
rect 501275 374884 501287 374918
rect 501287 374884 501309 374918
rect 501347 374884 501355 374918
rect 501355 374884 501381 374918
rect 501419 374884 501423 374918
rect 501423 374884 501453 374918
rect 501491 374884 501525 374918
rect 501563 374884 501593 374918
rect 501593 374884 501597 374918
rect 501635 374884 501661 374918
rect 501661 374884 501669 374918
rect 501707 374884 501729 374918
rect 501729 374884 501741 374918
rect 501779 374884 501797 374918
rect 501797 374884 501813 374918
rect 501851 374884 501865 374918
rect 501865 374884 501885 374918
rect 501131 374426 501151 374460
rect 501151 374426 501165 374460
rect 501203 374426 501219 374460
rect 501219 374426 501237 374460
rect 501275 374426 501287 374460
rect 501287 374426 501309 374460
rect 501347 374426 501355 374460
rect 501355 374426 501381 374460
rect 501419 374426 501423 374460
rect 501423 374426 501453 374460
rect 501491 374426 501525 374460
rect 501563 374426 501593 374460
rect 501593 374426 501597 374460
rect 501635 374426 501661 374460
rect 501661 374426 501669 374460
rect 501707 374426 501729 374460
rect 501729 374426 501741 374460
rect 501779 374426 501797 374460
rect 501797 374426 501813 374460
rect 501851 374426 501865 374460
rect 501865 374426 501885 374460
rect 501131 373968 501151 374002
rect 501151 373968 501165 374002
rect 501203 373968 501219 374002
rect 501219 373968 501237 374002
rect 501275 373968 501287 374002
rect 501287 373968 501309 374002
rect 501347 373968 501355 374002
rect 501355 373968 501381 374002
rect 501419 373968 501423 374002
rect 501423 373968 501453 374002
rect 501491 373968 501525 374002
rect 501563 373968 501593 374002
rect 501593 373968 501597 374002
rect 501635 373968 501661 374002
rect 501661 373968 501669 374002
rect 501707 373968 501729 374002
rect 501729 373968 501741 374002
rect 501779 373968 501797 374002
rect 501797 373968 501813 374002
rect 501851 373968 501865 374002
rect 501865 373968 501885 374002
rect 501131 373510 501151 373544
rect 501151 373510 501165 373544
rect 501203 373510 501219 373544
rect 501219 373510 501237 373544
rect 501275 373510 501287 373544
rect 501287 373510 501309 373544
rect 501347 373510 501355 373544
rect 501355 373510 501381 373544
rect 501419 373510 501423 373544
rect 501423 373510 501453 373544
rect 501491 373510 501525 373544
rect 501563 373510 501593 373544
rect 501593 373510 501597 373544
rect 501635 373510 501661 373544
rect 501661 373510 501669 373544
rect 501707 373510 501729 373544
rect 501729 373510 501741 373544
rect 501779 373510 501797 373544
rect 501797 373510 501813 373544
rect 501851 373510 501865 373544
rect 501865 373510 501885 373544
rect 502491 377461 502525 377495
rect 502491 377061 502525 377095
rect 502491 376661 502525 376695
rect 502491 376261 502525 376295
rect 502491 375861 502525 375895
rect 502491 375461 502525 375495
rect 502161 373491 502195 373525
rect 502491 375061 502525 375095
rect 502491 374661 502525 374695
rect 504371 377265 504405 377299
rect 504371 376865 504405 376899
rect 504639 377401 504673 377435
rect 504711 377401 504741 377435
rect 504741 377401 504745 377435
rect 504783 377401 504809 377435
rect 504809 377401 504817 377435
rect 504855 377401 504877 377435
rect 504877 377401 504889 377435
rect 504927 377401 504945 377435
rect 504945 377401 504961 377435
rect 504999 377401 505013 377435
rect 505013 377401 505033 377435
rect 505071 377401 505081 377435
rect 505081 377401 505105 377435
rect 505143 377401 505149 377435
rect 505149 377401 505177 377435
rect 505215 377401 505217 377435
rect 505217 377401 505249 377435
rect 505287 377401 505319 377435
rect 505319 377401 505321 377435
rect 505359 377401 505387 377435
rect 505387 377401 505393 377435
rect 505431 377401 505455 377435
rect 505455 377401 505465 377435
rect 505503 377401 505523 377435
rect 505523 377401 505537 377435
rect 505575 377401 505591 377435
rect 505591 377401 505609 377435
rect 505647 377401 505659 377435
rect 505659 377401 505681 377435
rect 505719 377401 505727 377435
rect 505727 377401 505753 377435
rect 505791 377401 505795 377435
rect 505795 377401 505825 377435
rect 505863 377401 505897 377435
rect 504541 377355 504575 377389
rect 506003 377355 506037 377389
rect 504639 376943 504673 376977
rect 504711 376943 504741 376977
rect 504741 376943 504745 376977
rect 504783 376943 504809 376977
rect 504809 376943 504817 376977
rect 504855 376943 504877 376977
rect 504877 376943 504889 376977
rect 504927 376943 504945 376977
rect 504945 376943 504961 376977
rect 504999 376943 505013 376977
rect 505013 376943 505033 376977
rect 505071 376943 505081 376977
rect 505081 376943 505105 376977
rect 505143 376943 505149 376977
rect 505149 376943 505177 376977
rect 505215 376943 505217 376977
rect 505217 376943 505249 376977
rect 505287 376943 505319 376977
rect 505319 376943 505321 376977
rect 505359 376943 505387 376977
rect 505387 376943 505393 376977
rect 505431 376943 505455 376977
rect 505455 376943 505465 376977
rect 505503 376943 505523 376977
rect 505523 376943 505537 376977
rect 505575 376943 505591 376977
rect 505591 376943 505609 376977
rect 505647 376943 505659 376977
rect 505659 376943 505681 376977
rect 505719 376943 505727 376977
rect 505727 376943 505753 376977
rect 505791 376943 505795 376977
rect 505795 376943 505825 376977
rect 505863 376943 505897 376977
rect 504371 376465 504405 376499
rect 504371 376065 504405 376099
rect 504371 375665 504405 375699
rect 504371 375265 504405 375299
rect 504371 374865 504405 374899
rect 504639 376485 504673 376519
rect 504711 376485 504741 376519
rect 504741 376485 504745 376519
rect 504783 376485 504809 376519
rect 504809 376485 504817 376519
rect 504855 376485 504877 376519
rect 504877 376485 504889 376519
rect 504927 376485 504945 376519
rect 504945 376485 504961 376519
rect 504999 376485 505013 376519
rect 505013 376485 505033 376519
rect 505071 376485 505081 376519
rect 505081 376485 505105 376519
rect 505143 376485 505149 376519
rect 505149 376485 505177 376519
rect 505215 376485 505217 376519
rect 505217 376485 505249 376519
rect 505287 376485 505319 376519
rect 505319 376485 505321 376519
rect 505359 376485 505387 376519
rect 505387 376485 505393 376519
rect 505431 376485 505455 376519
rect 505455 376485 505465 376519
rect 505503 376485 505523 376519
rect 505523 376485 505537 376519
rect 505575 376485 505591 376519
rect 505591 376485 505609 376519
rect 505647 376485 505659 376519
rect 505659 376485 505681 376519
rect 505719 376485 505727 376519
rect 505727 376485 505753 376519
rect 505791 376485 505795 376519
rect 505795 376485 505825 376519
rect 505863 376485 505897 376519
rect 504639 376027 504673 376061
rect 504711 376027 504741 376061
rect 504741 376027 504745 376061
rect 504783 376027 504809 376061
rect 504809 376027 504817 376061
rect 504855 376027 504877 376061
rect 504877 376027 504889 376061
rect 504927 376027 504945 376061
rect 504945 376027 504961 376061
rect 504999 376027 505013 376061
rect 505013 376027 505033 376061
rect 505071 376027 505081 376061
rect 505081 376027 505105 376061
rect 505143 376027 505149 376061
rect 505149 376027 505177 376061
rect 505215 376027 505217 376061
rect 505217 376027 505249 376061
rect 505287 376027 505319 376061
rect 505319 376027 505321 376061
rect 505359 376027 505387 376061
rect 505387 376027 505393 376061
rect 505431 376027 505455 376061
rect 505455 376027 505465 376061
rect 505503 376027 505523 376061
rect 505523 376027 505537 376061
rect 505575 376027 505591 376061
rect 505591 376027 505609 376061
rect 505647 376027 505659 376061
rect 505659 376027 505681 376061
rect 505719 376027 505727 376061
rect 505727 376027 505753 376061
rect 505791 376027 505795 376061
rect 505795 376027 505825 376061
rect 505863 376027 505897 376061
rect 504639 375569 504673 375603
rect 504711 375569 504741 375603
rect 504741 375569 504745 375603
rect 504783 375569 504809 375603
rect 504809 375569 504817 375603
rect 504855 375569 504877 375603
rect 504877 375569 504889 375603
rect 504927 375569 504945 375603
rect 504945 375569 504961 375603
rect 504999 375569 505013 375603
rect 505013 375569 505033 375603
rect 505071 375569 505081 375603
rect 505081 375569 505105 375603
rect 505143 375569 505149 375603
rect 505149 375569 505177 375603
rect 505215 375569 505217 375603
rect 505217 375569 505249 375603
rect 505287 375569 505319 375603
rect 505319 375569 505321 375603
rect 505359 375569 505387 375603
rect 505387 375569 505393 375603
rect 505431 375569 505455 375603
rect 505455 375569 505465 375603
rect 505503 375569 505523 375603
rect 505523 375569 505537 375603
rect 505575 375569 505591 375603
rect 505591 375569 505609 375603
rect 505647 375569 505659 375603
rect 505659 375569 505681 375603
rect 505719 375569 505727 375603
rect 505727 375569 505753 375603
rect 505791 375569 505795 375603
rect 505795 375569 505825 375603
rect 505863 375569 505897 375603
rect 504639 375111 504673 375145
rect 504711 375111 504741 375145
rect 504741 375111 504745 375145
rect 504783 375111 504809 375145
rect 504809 375111 504817 375145
rect 504855 375111 504877 375145
rect 504877 375111 504889 375145
rect 504927 375111 504945 375145
rect 504945 375111 504961 375145
rect 504999 375111 505013 375145
rect 505013 375111 505033 375145
rect 505071 375111 505081 375145
rect 505081 375111 505105 375145
rect 505143 375111 505149 375145
rect 505149 375111 505177 375145
rect 505215 375111 505217 375145
rect 505217 375111 505249 375145
rect 505287 375111 505319 375145
rect 505319 375111 505321 375145
rect 505359 375111 505387 375145
rect 505387 375111 505393 375145
rect 505431 375111 505455 375145
rect 505455 375111 505465 375145
rect 505503 375111 505523 375145
rect 505523 375111 505537 375145
rect 505575 375111 505591 375145
rect 505591 375111 505609 375145
rect 505647 375111 505659 375145
rect 505659 375111 505681 375145
rect 505719 375111 505727 375145
rect 505727 375111 505753 375145
rect 505791 375111 505795 375145
rect 505795 375111 505825 375145
rect 505863 375111 505897 375145
rect 504639 374653 504673 374687
rect 504711 374653 504741 374687
rect 504741 374653 504745 374687
rect 504783 374653 504809 374687
rect 504809 374653 504817 374687
rect 504855 374653 504877 374687
rect 504877 374653 504889 374687
rect 504927 374653 504945 374687
rect 504945 374653 504961 374687
rect 504999 374653 505013 374687
rect 505013 374653 505033 374687
rect 505071 374653 505081 374687
rect 505081 374653 505105 374687
rect 505143 374653 505149 374687
rect 505149 374653 505177 374687
rect 505215 374653 505217 374687
rect 505217 374653 505249 374687
rect 505287 374653 505319 374687
rect 505319 374653 505321 374687
rect 505359 374653 505387 374687
rect 505387 374653 505393 374687
rect 505431 374653 505455 374687
rect 505455 374653 505465 374687
rect 505503 374653 505523 374687
rect 505523 374653 505537 374687
rect 505575 374653 505591 374687
rect 505591 374653 505609 374687
rect 505647 374653 505659 374687
rect 505659 374653 505681 374687
rect 505719 374653 505727 374687
rect 505727 374653 505753 374687
rect 505791 374653 505795 374687
rect 505795 374653 505825 374687
rect 505863 374653 505897 374687
rect 506105 376343 506139 376377
rect 506251 377265 506285 377299
rect 506251 376865 506285 376899
rect 506251 376465 506285 376499
rect 506251 376065 506285 376099
rect 506251 375665 506285 375699
rect 506251 375265 506285 375299
rect 506251 374865 506285 374899
rect 508131 377485 508165 377519
rect 508131 377085 508165 377119
rect 508131 376685 508165 376719
rect 508131 376285 508165 376319
rect 508131 375885 508165 375919
rect 508131 375485 508165 375519
rect 508131 375085 508165 375119
rect 508131 374685 508165 374719
rect 502491 374261 502525 374295
rect 508131 374285 508165 374319
rect 510011 381085 510045 381119
rect 510011 380685 510045 380719
rect 510011 380285 510045 380319
rect 510011 379885 510045 379919
rect 510011 379485 510045 379519
rect 510011 379085 510045 379119
rect 510011 378685 510045 378719
rect 510011 378285 510045 378319
rect 510011 377885 510045 377919
rect 511891 381209 511925 381243
rect 511891 380809 511925 380843
rect 511891 380409 511925 380443
rect 511891 380009 511925 380043
rect 511891 379609 511925 379643
rect 511891 379209 511925 379243
rect 511891 378809 511925 378843
rect 511891 378409 511925 378443
rect 511891 378009 511925 378043
rect 513771 384809 513805 384843
rect 513771 384409 513805 384443
rect 513771 384009 513805 384043
rect 513771 383609 513805 383643
rect 513771 383209 513805 383243
rect 513771 382809 513805 382843
rect 513771 382409 513805 382443
rect 513771 382009 513805 382043
rect 513771 381609 513805 381643
rect 513771 381209 513805 381243
rect 513771 380809 513805 380843
rect 513771 380409 513805 380443
rect 513771 380009 513805 380043
rect 513771 379609 513805 379643
rect 513771 379209 513805 379243
rect 513771 378809 513805 378843
rect 513771 378409 513805 378443
rect 513771 378009 513805 378043
rect 515651 384809 515685 384843
rect 515651 384409 515685 384443
rect 515651 384009 515685 384043
rect 515651 383609 515685 383643
rect 515651 383209 515685 383243
rect 515651 382809 515685 382843
rect 515651 382409 515685 382443
rect 515651 382009 515685 382043
rect 515651 381609 515685 381643
rect 515651 381209 515685 381243
rect 515651 380809 515685 380843
rect 515651 380409 515685 380443
rect 515651 380009 515685 380043
rect 515651 379609 515685 379643
rect 515651 379209 515685 379243
rect 515651 378809 515685 378843
rect 515651 378409 515685 378443
rect 515651 378009 515685 378043
rect 517531 384809 517565 384843
rect 517531 384409 517565 384443
rect 517531 384009 517565 384043
rect 517531 383609 517565 383643
rect 517531 383209 517565 383243
rect 517531 382809 517565 382843
rect 519411 384791 519445 384825
rect 519411 384591 519445 384625
rect 519679 384595 520217 384989
rect 520639 384595 521177 384989
rect 521291 384791 521325 384825
rect 521291 384591 521325 384625
rect 519411 384391 519445 384425
rect 519411 384191 519445 384225
rect 521291 384391 521325 384425
rect 521291 384191 521325 384225
rect 519411 383991 519445 384025
rect 519411 383791 519445 383825
rect 519411 383591 519445 383625
rect 521291 383991 521325 384025
rect 521291 383791 521325 383825
rect 521291 383591 521325 383625
rect 519411 383391 519445 383425
rect 519411 383191 519445 383225
rect 519411 382991 519445 383025
rect 521291 383391 521325 383425
rect 521291 383191 521325 383225
rect 519411 382791 519445 382825
rect 519679 382588 520217 382982
rect 520639 382588 521177 382982
rect 521291 382991 521325 383025
rect 521291 382791 521325 382825
rect 523171 384707 523205 384741
rect 523171 384307 523205 384341
rect 523439 385463 523473 385497
rect 523511 385463 523541 385497
rect 523541 385463 523545 385497
rect 523583 385463 523609 385497
rect 523609 385463 523617 385497
rect 523655 385463 523677 385497
rect 523677 385463 523689 385497
rect 523727 385463 523745 385497
rect 523745 385463 523761 385497
rect 523799 385463 523813 385497
rect 523813 385463 523833 385497
rect 523871 385463 523881 385497
rect 523881 385463 523905 385497
rect 523943 385463 523949 385497
rect 523949 385463 523977 385497
rect 524015 385463 524017 385497
rect 524017 385463 524049 385497
rect 524087 385463 524119 385497
rect 524119 385463 524121 385497
rect 524159 385463 524187 385497
rect 524187 385463 524193 385497
rect 524231 385463 524255 385497
rect 524255 385463 524265 385497
rect 524303 385463 524323 385497
rect 524323 385463 524337 385497
rect 524375 385463 524391 385497
rect 524391 385463 524409 385497
rect 524447 385463 524459 385497
rect 524459 385463 524481 385497
rect 524519 385463 524527 385497
rect 524527 385463 524553 385497
rect 524591 385463 524595 385497
rect 524595 385463 524625 385497
rect 524663 385463 524697 385497
rect 523439 385005 523473 385039
rect 523511 385005 523541 385039
rect 523541 385005 523545 385039
rect 523583 385005 523609 385039
rect 523609 385005 523617 385039
rect 523655 385005 523677 385039
rect 523677 385005 523689 385039
rect 523727 385005 523745 385039
rect 523745 385005 523761 385039
rect 523799 385005 523813 385039
rect 523813 385005 523833 385039
rect 523871 385005 523881 385039
rect 523881 385005 523905 385039
rect 523943 385005 523949 385039
rect 523949 385005 523977 385039
rect 524015 385005 524017 385039
rect 524017 385005 524049 385039
rect 524087 385005 524119 385039
rect 524119 385005 524121 385039
rect 524159 385005 524187 385039
rect 524187 385005 524193 385039
rect 524231 385005 524255 385039
rect 524255 385005 524265 385039
rect 524303 385005 524323 385039
rect 524323 385005 524337 385039
rect 524375 385005 524391 385039
rect 524391 385005 524409 385039
rect 524447 385005 524459 385039
rect 524459 385005 524481 385039
rect 524519 385005 524527 385039
rect 524527 385005 524553 385039
rect 524591 385005 524595 385039
rect 524595 385005 524625 385039
rect 524663 385005 524697 385039
rect 523439 384547 523473 384581
rect 523511 384547 523541 384581
rect 523541 384547 523545 384581
rect 523583 384547 523609 384581
rect 523609 384547 523617 384581
rect 523655 384547 523677 384581
rect 523677 384547 523689 384581
rect 523727 384547 523745 384581
rect 523745 384547 523761 384581
rect 523799 384547 523813 384581
rect 523813 384547 523833 384581
rect 523871 384547 523881 384581
rect 523881 384547 523905 384581
rect 523943 384547 523949 384581
rect 523949 384547 523977 384581
rect 524015 384547 524017 384581
rect 524017 384547 524049 384581
rect 524087 384547 524119 384581
rect 524119 384547 524121 384581
rect 524159 384547 524187 384581
rect 524187 384547 524193 384581
rect 524231 384547 524255 384581
rect 524255 384547 524265 384581
rect 524303 384547 524323 384581
rect 524323 384547 524337 384581
rect 524375 384547 524391 384581
rect 524391 384547 524409 384581
rect 524447 384547 524459 384581
rect 524459 384547 524481 384581
rect 524519 384547 524527 384581
rect 524527 384547 524553 384581
rect 524591 384547 524595 384581
rect 524595 384547 524625 384581
rect 524663 384547 524697 384581
rect 523439 384089 523473 384123
rect 523511 384089 523541 384123
rect 523541 384089 523545 384123
rect 523583 384089 523609 384123
rect 523609 384089 523617 384123
rect 523655 384089 523677 384123
rect 523677 384089 523689 384123
rect 523727 384089 523745 384123
rect 523745 384089 523761 384123
rect 523799 384089 523813 384123
rect 523813 384089 523833 384123
rect 523871 384089 523881 384123
rect 523881 384089 523905 384123
rect 523943 384089 523949 384123
rect 523949 384089 523977 384123
rect 524015 384089 524017 384123
rect 524017 384089 524049 384123
rect 524087 384089 524119 384123
rect 524119 384089 524121 384123
rect 524159 384089 524187 384123
rect 524187 384089 524193 384123
rect 524231 384089 524255 384123
rect 524255 384089 524265 384123
rect 524303 384089 524323 384123
rect 524323 384089 524337 384123
rect 524375 384089 524391 384123
rect 524391 384089 524409 384123
rect 524447 384089 524459 384123
rect 524459 384089 524481 384123
rect 524519 384089 524527 384123
rect 524527 384089 524553 384123
rect 524591 384089 524595 384123
rect 524595 384089 524625 384123
rect 524663 384089 524697 384123
rect 523171 383907 523205 383941
rect 523171 383507 523205 383541
rect 523171 383107 523205 383141
rect 523171 382707 523205 382741
rect 523439 383631 523473 383665
rect 523511 383631 523541 383665
rect 523541 383631 523545 383665
rect 523583 383631 523609 383665
rect 523609 383631 523617 383665
rect 523655 383631 523677 383665
rect 523677 383631 523689 383665
rect 523727 383631 523745 383665
rect 523745 383631 523761 383665
rect 523799 383631 523813 383665
rect 523813 383631 523833 383665
rect 523871 383631 523881 383665
rect 523881 383631 523905 383665
rect 523943 383631 523949 383665
rect 523949 383631 523977 383665
rect 524015 383631 524017 383665
rect 524017 383631 524049 383665
rect 524087 383631 524119 383665
rect 524119 383631 524121 383665
rect 524159 383631 524187 383665
rect 524187 383631 524193 383665
rect 524231 383631 524255 383665
rect 524255 383631 524265 383665
rect 524303 383631 524323 383665
rect 524323 383631 524337 383665
rect 524375 383631 524391 383665
rect 524391 383631 524409 383665
rect 524447 383631 524459 383665
rect 524459 383631 524481 383665
rect 524519 383631 524527 383665
rect 524527 383631 524553 383665
rect 524591 383631 524595 383665
rect 524595 383631 524625 383665
rect 524663 383631 524697 383665
rect 523439 383173 523473 383207
rect 523511 383173 523541 383207
rect 523541 383173 523545 383207
rect 523583 383173 523609 383207
rect 523609 383173 523617 383207
rect 523655 383173 523677 383207
rect 523677 383173 523689 383207
rect 523727 383173 523745 383207
rect 523745 383173 523761 383207
rect 523799 383173 523813 383207
rect 523813 383173 523833 383207
rect 523871 383173 523881 383207
rect 523881 383173 523905 383207
rect 523943 383173 523949 383207
rect 523949 383173 523977 383207
rect 524015 383173 524017 383207
rect 524017 383173 524049 383207
rect 524087 383173 524119 383207
rect 524119 383173 524121 383207
rect 524159 383173 524187 383207
rect 524187 383173 524193 383207
rect 524231 383173 524255 383207
rect 524255 383173 524265 383207
rect 524303 383173 524323 383207
rect 524323 383173 524337 383207
rect 524375 383173 524391 383207
rect 524391 383173 524409 383207
rect 524447 383173 524459 383207
rect 524459 383173 524481 383207
rect 524519 383173 524527 383207
rect 524527 383173 524553 383207
rect 524591 383173 524595 383207
rect 524595 383173 524625 383207
rect 524663 383173 524697 383207
rect 517531 382409 517565 382443
rect 517531 382009 517565 382043
rect 523171 382307 523205 382341
rect 523171 381907 523205 381941
rect 517531 381609 517565 381643
rect 517531 381209 517565 381243
rect 517531 380809 517565 380843
rect 517531 380409 517565 380443
rect 517531 380009 517565 380043
rect 517531 379609 517565 379643
rect 519411 381557 519445 381591
rect 519411 381357 519445 381391
rect 519679 381361 520217 381755
rect 520639 381361 521177 381755
rect 521291 381557 521325 381591
rect 521291 381357 521325 381391
rect 519411 381157 519445 381191
rect 519411 380957 519445 380991
rect 521291 381157 521325 381191
rect 521291 380957 521325 380991
rect 519411 380757 519445 380791
rect 519411 380557 519445 380591
rect 519411 380357 519445 380391
rect 521291 380757 521325 380791
rect 521291 380557 521325 380591
rect 521291 380357 521325 380391
rect 519411 380157 519445 380191
rect 519411 379957 519445 379991
rect 519411 379757 519445 379791
rect 521291 380157 521325 380191
rect 521291 379957 521325 379991
rect 519411 379557 519445 379591
rect 519679 379354 520217 379748
rect 520639 379354 521177 379748
rect 521291 379757 521325 379791
rect 521291 379557 521325 379591
rect 523171 381507 523205 381541
rect 523439 382715 523473 382749
rect 523511 382715 523541 382749
rect 523541 382715 523545 382749
rect 523583 382715 523609 382749
rect 523609 382715 523617 382749
rect 523655 382715 523677 382749
rect 523677 382715 523689 382749
rect 523727 382715 523745 382749
rect 523745 382715 523761 382749
rect 523799 382715 523813 382749
rect 523813 382715 523833 382749
rect 523871 382715 523881 382749
rect 523881 382715 523905 382749
rect 523943 382715 523949 382749
rect 523949 382715 523977 382749
rect 524015 382715 524017 382749
rect 524017 382715 524049 382749
rect 524087 382715 524119 382749
rect 524119 382715 524121 382749
rect 524159 382715 524187 382749
rect 524187 382715 524193 382749
rect 524231 382715 524255 382749
rect 524255 382715 524265 382749
rect 524303 382715 524323 382749
rect 524323 382715 524337 382749
rect 524375 382715 524391 382749
rect 524391 382715 524409 382749
rect 524447 382715 524459 382749
rect 524459 382715 524481 382749
rect 524519 382715 524527 382749
rect 524527 382715 524553 382749
rect 524591 382715 524595 382749
rect 524595 382715 524625 382749
rect 524663 382715 524697 382749
rect 523439 382257 523473 382291
rect 523511 382257 523541 382291
rect 523541 382257 523545 382291
rect 523583 382257 523609 382291
rect 523609 382257 523617 382291
rect 523655 382257 523677 382291
rect 523677 382257 523689 382291
rect 523727 382257 523745 382291
rect 523745 382257 523761 382291
rect 523799 382257 523813 382291
rect 523813 382257 523833 382291
rect 523871 382257 523881 382291
rect 523881 382257 523905 382291
rect 523943 382257 523949 382291
rect 523949 382257 523977 382291
rect 524015 382257 524017 382291
rect 524017 382257 524049 382291
rect 524087 382257 524119 382291
rect 524119 382257 524121 382291
rect 524159 382257 524187 382291
rect 524187 382257 524193 382291
rect 524231 382257 524255 382291
rect 524255 382257 524265 382291
rect 524303 382257 524323 382291
rect 524323 382257 524337 382291
rect 524375 382257 524391 382291
rect 524391 382257 524409 382291
rect 524447 382257 524459 382291
rect 524459 382257 524481 382291
rect 524519 382257 524527 382291
rect 524527 382257 524553 382291
rect 524591 382257 524595 382291
rect 524595 382257 524625 382291
rect 524663 382257 524697 382291
rect 523439 381799 523473 381833
rect 523511 381799 523541 381833
rect 523541 381799 523545 381833
rect 523583 381799 523609 381833
rect 523609 381799 523617 381833
rect 523655 381799 523677 381833
rect 523677 381799 523689 381833
rect 523727 381799 523745 381833
rect 523745 381799 523761 381833
rect 523799 381799 523813 381833
rect 523813 381799 523833 381833
rect 523871 381799 523881 381833
rect 523881 381799 523905 381833
rect 523943 381799 523949 381833
rect 523949 381799 523977 381833
rect 524015 381799 524017 381833
rect 524017 381799 524049 381833
rect 524087 381799 524119 381833
rect 524119 381799 524121 381833
rect 524159 381799 524187 381833
rect 524187 381799 524193 381833
rect 524231 381799 524255 381833
rect 524255 381799 524265 381833
rect 524303 381799 524323 381833
rect 524323 381799 524337 381833
rect 524375 381799 524391 381833
rect 524391 381799 524409 381833
rect 524447 381799 524459 381833
rect 524459 381799 524481 381833
rect 524519 381799 524527 381833
rect 524527 381799 524553 381833
rect 524591 381799 524595 381833
rect 524595 381799 524625 381833
rect 524663 381799 524697 381833
rect 523439 381341 523473 381375
rect 523511 381341 523541 381375
rect 523541 381341 523545 381375
rect 523583 381341 523609 381375
rect 523609 381341 523617 381375
rect 523655 381341 523677 381375
rect 523677 381341 523689 381375
rect 523727 381341 523745 381375
rect 523745 381341 523761 381375
rect 523799 381341 523813 381375
rect 523813 381341 523833 381375
rect 523871 381341 523881 381375
rect 523881 381341 523905 381375
rect 523943 381341 523949 381375
rect 523949 381341 523977 381375
rect 524015 381341 524017 381375
rect 524017 381341 524049 381375
rect 524087 381341 524119 381375
rect 524119 381341 524121 381375
rect 524159 381341 524187 381375
rect 524187 381341 524193 381375
rect 524231 381341 524255 381375
rect 524255 381341 524265 381375
rect 524303 381341 524323 381375
rect 524323 381341 524337 381375
rect 524375 381341 524391 381375
rect 524391 381341 524409 381375
rect 524447 381341 524459 381375
rect 524459 381341 524481 381375
rect 524519 381341 524527 381375
rect 524527 381341 524553 381375
rect 524591 381341 524595 381375
rect 524595 381341 524625 381375
rect 524663 381341 524697 381375
rect 523171 381107 523205 381141
rect 523171 380707 523205 380741
rect 523171 380307 523205 380341
rect 523439 380883 523473 380917
rect 523511 380883 523541 380917
rect 523541 380883 523545 380917
rect 523583 380883 523609 380917
rect 523609 380883 523617 380917
rect 523655 380883 523677 380917
rect 523677 380883 523689 380917
rect 523727 380883 523745 380917
rect 523745 380883 523761 380917
rect 523799 380883 523813 380917
rect 523813 380883 523833 380917
rect 523871 380883 523881 380917
rect 523881 380883 523905 380917
rect 523943 380883 523949 380917
rect 523949 380883 523977 380917
rect 524015 380883 524017 380917
rect 524017 380883 524049 380917
rect 524087 380883 524119 380917
rect 524119 380883 524121 380917
rect 524159 380883 524187 380917
rect 524187 380883 524193 380917
rect 524231 380883 524255 380917
rect 524255 380883 524265 380917
rect 524303 380883 524323 380917
rect 524323 380883 524337 380917
rect 524375 380883 524391 380917
rect 524391 380883 524409 380917
rect 524447 380883 524459 380917
rect 524459 380883 524481 380917
rect 524519 380883 524527 380917
rect 524527 380883 524553 380917
rect 524591 380883 524595 380917
rect 524595 380883 524625 380917
rect 524663 380883 524697 380917
rect 524805 380575 524839 380609
rect 523439 380425 523473 380459
rect 523511 380425 523541 380459
rect 523541 380425 523545 380459
rect 523583 380425 523609 380459
rect 523609 380425 523617 380459
rect 523655 380425 523677 380459
rect 523677 380425 523689 380459
rect 523727 380425 523745 380459
rect 523745 380425 523761 380459
rect 523799 380425 523813 380459
rect 523813 380425 523833 380459
rect 523871 380425 523881 380459
rect 523881 380425 523905 380459
rect 523943 380425 523949 380459
rect 523949 380425 523977 380459
rect 524015 380425 524017 380459
rect 524017 380425 524049 380459
rect 524087 380425 524119 380459
rect 524119 380425 524121 380459
rect 524159 380425 524187 380459
rect 524187 380425 524193 380459
rect 524231 380425 524255 380459
rect 524255 380425 524265 380459
rect 524303 380425 524323 380459
rect 524323 380425 524337 380459
rect 524375 380425 524391 380459
rect 524391 380425 524409 380459
rect 524447 380425 524459 380459
rect 524459 380425 524481 380459
rect 524519 380425 524527 380459
rect 524527 380425 524553 380459
rect 524591 380425 524595 380459
rect 524595 380425 524625 380459
rect 524663 380425 524697 380459
rect 523171 379907 523205 379941
rect 523171 379507 523205 379541
rect 517531 379209 517565 379243
rect 517531 378809 517565 378843
rect 517531 378409 517565 378443
rect 517531 378009 517565 378043
rect 523171 379107 523205 379141
rect 523439 379967 523473 380001
rect 523511 379967 523541 380001
rect 523541 379967 523545 380001
rect 523583 379967 523609 380001
rect 523609 379967 523617 380001
rect 523655 379967 523677 380001
rect 523677 379967 523689 380001
rect 523727 379967 523745 380001
rect 523745 379967 523761 380001
rect 523799 379967 523813 380001
rect 523813 379967 523833 380001
rect 523871 379967 523881 380001
rect 523881 379967 523905 380001
rect 523943 379967 523949 380001
rect 523949 379967 523977 380001
rect 524015 379967 524017 380001
rect 524017 379967 524049 380001
rect 524087 379967 524119 380001
rect 524119 379967 524121 380001
rect 524159 379967 524187 380001
rect 524187 379967 524193 380001
rect 524231 379967 524255 380001
rect 524255 379967 524265 380001
rect 524303 379967 524323 380001
rect 524323 379967 524337 380001
rect 524375 379967 524391 380001
rect 524391 379967 524409 380001
rect 524447 379967 524459 380001
rect 524459 379967 524481 380001
rect 524519 379967 524527 380001
rect 524527 379967 524553 380001
rect 524591 379967 524595 380001
rect 524595 379967 524625 380001
rect 524663 379967 524697 380001
rect 523439 379509 523473 379543
rect 523511 379509 523541 379543
rect 523541 379509 523545 379543
rect 523583 379509 523609 379543
rect 523609 379509 523617 379543
rect 523655 379509 523677 379543
rect 523677 379509 523689 379543
rect 523727 379509 523745 379543
rect 523745 379509 523761 379543
rect 523799 379509 523813 379543
rect 523813 379509 523833 379543
rect 523871 379509 523881 379543
rect 523881 379509 523905 379543
rect 523943 379509 523949 379543
rect 523949 379509 523977 379543
rect 524015 379509 524017 379543
rect 524017 379509 524049 379543
rect 524087 379509 524119 379543
rect 524119 379509 524121 379543
rect 524159 379509 524187 379543
rect 524187 379509 524193 379543
rect 524231 379509 524255 379543
rect 524255 379509 524265 379543
rect 524303 379509 524323 379543
rect 524323 379509 524337 379543
rect 524375 379509 524391 379543
rect 524391 379509 524409 379543
rect 524447 379509 524459 379543
rect 524459 379509 524481 379543
rect 524519 379509 524527 379543
rect 524527 379509 524553 379543
rect 524591 379509 524595 379543
rect 524595 379509 524625 379543
rect 524663 379509 524697 379543
rect 523171 378707 523205 378741
rect 523439 379051 523473 379085
rect 523511 379051 523541 379085
rect 523541 379051 523545 379085
rect 523583 379051 523609 379085
rect 523609 379051 523617 379085
rect 523655 379051 523677 379085
rect 523677 379051 523689 379085
rect 523727 379051 523745 379085
rect 523745 379051 523761 379085
rect 523799 379051 523813 379085
rect 523813 379051 523833 379085
rect 523871 379051 523881 379085
rect 523881 379051 523905 379085
rect 523943 379051 523949 379085
rect 523949 379051 523977 379085
rect 524015 379051 524017 379085
rect 524017 379051 524049 379085
rect 524087 379051 524119 379085
rect 524119 379051 524121 379085
rect 524159 379051 524187 379085
rect 524187 379051 524193 379085
rect 524231 379051 524255 379085
rect 524255 379051 524265 379085
rect 524303 379051 524323 379085
rect 524323 379051 524337 379085
rect 524375 379051 524391 379085
rect 524391 379051 524409 379085
rect 524447 379051 524459 379085
rect 524459 379051 524481 379085
rect 524519 379051 524527 379085
rect 524527 379051 524553 379085
rect 524591 379051 524595 379085
rect 524595 379051 524625 379085
rect 524663 379051 524697 379085
rect 523439 378593 523473 378627
rect 523511 378593 523541 378627
rect 523541 378593 523545 378627
rect 523583 378593 523609 378627
rect 523609 378593 523617 378627
rect 523655 378593 523677 378627
rect 523677 378593 523689 378627
rect 523727 378593 523745 378627
rect 523745 378593 523761 378627
rect 523799 378593 523813 378627
rect 523813 378593 523833 378627
rect 523871 378593 523881 378627
rect 523881 378593 523905 378627
rect 523943 378593 523949 378627
rect 523949 378593 523977 378627
rect 524015 378593 524017 378627
rect 524017 378593 524049 378627
rect 524087 378593 524119 378627
rect 524119 378593 524121 378627
rect 524159 378593 524187 378627
rect 524187 378593 524193 378627
rect 524231 378593 524255 378627
rect 524255 378593 524265 378627
rect 524303 378593 524323 378627
rect 524323 378593 524337 378627
rect 524375 378593 524391 378627
rect 524391 378593 524409 378627
rect 524447 378593 524459 378627
rect 524459 378593 524481 378627
rect 524519 378593 524527 378627
rect 524527 378593 524553 378627
rect 524591 378593 524595 378627
rect 524595 378593 524625 378627
rect 524663 378593 524697 378627
rect 523171 378307 523205 378341
rect 523171 377907 523205 377941
rect 510011 377485 510045 377519
rect 510011 377085 510045 377119
rect 510011 376685 510045 376719
rect 510011 376285 510045 376319
rect 510011 375885 510045 375919
rect 510011 375485 510045 375519
rect 510011 375085 510045 375119
rect 510011 374685 510045 374719
rect 511891 377265 511925 377299
rect 511891 376865 511925 376899
rect 512159 377401 512193 377435
rect 512231 377401 512261 377435
rect 512261 377401 512265 377435
rect 512303 377401 512329 377435
rect 512329 377401 512337 377435
rect 512375 377401 512397 377435
rect 512397 377401 512409 377435
rect 512447 377401 512465 377435
rect 512465 377401 512481 377435
rect 512519 377401 512533 377435
rect 512533 377401 512553 377435
rect 512591 377401 512601 377435
rect 512601 377401 512625 377435
rect 512663 377401 512669 377435
rect 512669 377401 512697 377435
rect 512735 377401 512737 377435
rect 512737 377401 512769 377435
rect 512807 377401 512839 377435
rect 512839 377401 512841 377435
rect 512879 377401 512907 377435
rect 512907 377401 512913 377435
rect 512951 377401 512975 377435
rect 512975 377401 512985 377435
rect 513023 377401 513043 377435
rect 513043 377401 513057 377435
rect 513095 377401 513111 377435
rect 513111 377401 513129 377435
rect 513167 377401 513179 377435
rect 513179 377401 513201 377435
rect 513239 377401 513247 377435
rect 513247 377401 513273 377435
rect 513311 377401 513315 377435
rect 513315 377401 513345 377435
rect 513383 377401 513417 377435
rect 512159 376943 512193 376977
rect 512231 376943 512261 376977
rect 512261 376943 512265 376977
rect 512303 376943 512329 376977
rect 512329 376943 512337 376977
rect 512375 376943 512397 376977
rect 512397 376943 512409 376977
rect 512447 376943 512465 376977
rect 512465 376943 512481 376977
rect 512519 376943 512533 376977
rect 512533 376943 512553 376977
rect 512591 376943 512601 376977
rect 512601 376943 512625 376977
rect 512663 376943 512669 376977
rect 512669 376943 512697 376977
rect 512735 376943 512737 376977
rect 512737 376943 512769 376977
rect 512807 376943 512839 376977
rect 512839 376943 512841 376977
rect 512879 376943 512907 376977
rect 512907 376943 512913 376977
rect 512951 376943 512975 376977
rect 512975 376943 512985 376977
rect 513023 376943 513043 376977
rect 513043 376943 513057 376977
rect 513095 376943 513111 376977
rect 513111 376943 513129 376977
rect 513167 376943 513179 376977
rect 513179 376943 513201 376977
rect 513239 376943 513247 376977
rect 513247 376943 513273 376977
rect 513311 376943 513315 376977
rect 513315 376943 513345 376977
rect 513383 376943 513417 376977
rect 511891 376465 511925 376499
rect 511891 376065 511925 376099
rect 511891 375665 511925 375699
rect 511891 375265 511925 375299
rect 511891 374865 511925 374899
rect 512159 376485 512193 376519
rect 512231 376485 512261 376519
rect 512261 376485 512265 376519
rect 512303 376485 512329 376519
rect 512329 376485 512337 376519
rect 512375 376485 512397 376519
rect 512397 376485 512409 376519
rect 512447 376485 512465 376519
rect 512465 376485 512481 376519
rect 512519 376485 512533 376519
rect 512533 376485 512553 376519
rect 512591 376485 512601 376519
rect 512601 376485 512625 376519
rect 512663 376485 512669 376519
rect 512669 376485 512697 376519
rect 512735 376485 512737 376519
rect 512737 376485 512769 376519
rect 512807 376485 512839 376519
rect 512839 376485 512841 376519
rect 512879 376485 512907 376519
rect 512907 376485 512913 376519
rect 512951 376485 512975 376519
rect 512975 376485 512985 376519
rect 513023 376485 513043 376519
rect 513043 376485 513057 376519
rect 513095 376485 513111 376519
rect 513111 376485 513129 376519
rect 513167 376485 513179 376519
rect 513179 376485 513201 376519
rect 513239 376485 513247 376519
rect 513247 376485 513273 376519
rect 513311 376485 513315 376519
rect 513315 376485 513345 376519
rect 513383 376485 513417 376519
rect 513517 376343 513551 376377
rect 512159 376027 512193 376061
rect 512231 376027 512261 376061
rect 512261 376027 512265 376061
rect 512303 376027 512329 376061
rect 512329 376027 512337 376061
rect 512375 376027 512397 376061
rect 512397 376027 512409 376061
rect 512447 376027 512465 376061
rect 512465 376027 512481 376061
rect 512519 376027 512533 376061
rect 512533 376027 512553 376061
rect 512591 376027 512601 376061
rect 512601 376027 512625 376061
rect 512663 376027 512669 376061
rect 512669 376027 512697 376061
rect 512735 376027 512737 376061
rect 512737 376027 512769 376061
rect 512807 376027 512839 376061
rect 512839 376027 512841 376061
rect 512879 376027 512907 376061
rect 512907 376027 512913 376061
rect 512951 376027 512975 376061
rect 512975 376027 512985 376061
rect 513023 376027 513043 376061
rect 513043 376027 513057 376061
rect 513095 376027 513111 376061
rect 513111 376027 513129 376061
rect 513167 376027 513179 376061
rect 513179 376027 513201 376061
rect 513239 376027 513247 376061
rect 513247 376027 513273 376061
rect 513311 376027 513315 376061
rect 513315 376027 513345 376061
rect 513383 376027 513417 376061
rect 512159 375569 512193 375603
rect 512231 375569 512261 375603
rect 512261 375569 512265 375603
rect 512303 375569 512329 375603
rect 512329 375569 512337 375603
rect 512375 375569 512397 375603
rect 512397 375569 512409 375603
rect 512447 375569 512465 375603
rect 512465 375569 512481 375603
rect 512519 375569 512533 375603
rect 512533 375569 512553 375603
rect 512591 375569 512601 375603
rect 512601 375569 512625 375603
rect 512663 375569 512669 375603
rect 512669 375569 512697 375603
rect 512735 375569 512737 375603
rect 512737 375569 512769 375603
rect 512807 375569 512839 375603
rect 512839 375569 512841 375603
rect 512879 375569 512907 375603
rect 512907 375569 512913 375603
rect 512951 375569 512975 375603
rect 512975 375569 512985 375603
rect 513023 375569 513043 375603
rect 513043 375569 513057 375603
rect 513095 375569 513111 375603
rect 513111 375569 513129 375603
rect 513167 375569 513179 375603
rect 513179 375569 513201 375603
rect 513239 375569 513247 375603
rect 513247 375569 513273 375603
rect 513311 375569 513315 375603
rect 513315 375569 513345 375603
rect 513383 375569 513417 375603
rect 512159 375111 512193 375145
rect 512231 375111 512261 375145
rect 512261 375111 512265 375145
rect 512303 375111 512329 375145
rect 512329 375111 512337 375145
rect 512375 375111 512397 375145
rect 512397 375111 512409 375145
rect 512447 375111 512465 375145
rect 512465 375111 512481 375145
rect 512519 375111 512533 375145
rect 512533 375111 512553 375145
rect 512591 375111 512601 375145
rect 512601 375111 512625 375145
rect 512663 375111 512669 375145
rect 512669 375111 512697 375145
rect 512735 375111 512737 375145
rect 512737 375111 512769 375145
rect 512807 375111 512839 375145
rect 512839 375111 512841 375145
rect 512879 375111 512907 375145
rect 512907 375111 512913 375145
rect 512951 375111 512975 375145
rect 512975 375111 512985 375145
rect 513023 375111 513043 375145
rect 513043 375111 513057 375145
rect 513095 375111 513111 375145
rect 513111 375111 513129 375145
rect 513167 375111 513179 375145
rect 513179 375111 513201 375145
rect 513239 375111 513247 375145
rect 513247 375111 513273 375145
rect 513311 375111 513315 375145
rect 513315 375111 513345 375145
rect 513383 375111 513417 375145
rect 512159 374653 512193 374687
rect 512231 374653 512261 374687
rect 512261 374653 512265 374687
rect 512303 374653 512329 374687
rect 512329 374653 512337 374687
rect 512375 374653 512397 374687
rect 512397 374653 512409 374687
rect 512447 374653 512465 374687
rect 512465 374653 512481 374687
rect 512519 374653 512533 374687
rect 512533 374653 512553 374687
rect 512591 374653 512601 374687
rect 512601 374653 512625 374687
rect 512663 374653 512669 374687
rect 512669 374653 512697 374687
rect 512735 374653 512737 374687
rect 512737 374653 512769 374687
rect 512807 374653 512839 374687
rect 512839 374653 512841 374687
rect 512879 374653 512907 374687
rect 512907 374653 512913 374687
rect 512951 374653 512975 374687
rect 512975 374653 512985 374687
rect 513023 374653 513043 374687
rect 513043 374653 513057 374687
rect 513095 374653 513111 374687
rect 513111 374653 513129 374687
rect 513167 374653 513179 374687
rect 513179 374653 513201 374687
rect 513239 374653 513247 374687
rect 513247 374653 513273 374687
rect 513311 374653 513315 374687
rect 513315 374653 513345 374687
rect 513383 374653 513417 374687
rect 512061 374595 512095 374629
rect 513771 377265 513805 377299
rect 513771 376865 513805 376899
rect 513771 376465 513805 376499
rect 513653 376343 513687 376377
rect 513771 376065 513805 376099
rect 513771 375665 513805 375699
rect 513771 375265 513805 375299
rect 515651 377343 515685 377377
rect 515651 377143 515685 377177
rect 515919 377147 516457 377541
rect 516879 377147 517417 377541
rect 517531 377343 517565 377377
rect 517531 377143 517565 377177
rect 515651 376943 515685 376977
rect 515651 376743 515685 376777
rect 517531 376943 517565 376977
rect 517531 376743 517565 376777
rect 515651 376543 515685 376577
rect 515651 376343 515685 376377
rect 515651 376143 515685 376177
rect 517531 376543 517565 376577
rect 517531 376343 517565 376377
rect 517531 376143 517565 376177
rect 515651 375943 515685 375977
rect 515651 375743 515685 375777
rect 515651 375543 515685 375577
rect 517531 375943 517565 375977
rect 517531 375743 517565 375777
rect 515651 375343 515685 375377
rect 515919 375140 516457 375534
rect 516879 375140 517417 375534
rect 517531 375543 517565 375577
rect 517531 375343 517565 375377
rect 519411 377343 519445 377377
rect 519411 377143 519445 377177
rect 519679 377147 520217 377541
rect 520639 377147 521177 377541
rect 521291 377343 521325 377377
rect 521291 377143 521325 377177
rect 519411 376943 519445 376977
rect 519411 376743 519445 376777
rect 521291 376943 521325 376977
rect 521291 376743 521325 376777
rect 519411 376543 519445 376577
rect 519411 376343 519445 376377
rect 519411 376143 519445 376177
rect 521291 376543 521325 376577
rect 521291 376343 521325 376377
rect 521291 376143 521325 376177
rect 519411 375943 519445 375977
rect 519411 375743 519445 375777
rect 519411 375543 519445 375577
rect 521291 375943 521325 375977
rect 521291 375743 521325 375777
rect 519411 375343 519445 375377
rect 519679 375140 520217 375534
rect 520639 375140 521177 375534
rect 521291 375543 521325 375577
rect 521291 375343 521325 375377
rect 523171 377507 523205 377541
rect 523439 378135 523473 378169
rect 523511 378135 523541 378169
rect 523541 378135 523545 378169
rect 523583 378135 523609 378169
rect 523609 378135 523617 378169
rect 523655 378135 523677 378169
rect 523677 378135 523689 378169
rect 523727 378135 523745 378169
rect 523745 378135 523761 378169
rect 523799 378135 523813 378169
rect 523813 378135 523833 378169
rect 523871 378135 523881 378169
rect 523881 378135 523905 378169
rect 523943 378135 523949 378169
rect 523949 378135 523977 378169
rect 524015 378135 524017 378169
rect 524017 378135 524049 378169
rect 524087 378135 524119 378169
rect 524119 378135 524121 378169
rect 524159 378135 524187 378169
rect 524187 378135 524193 378169
rect 524231 378135 524255 378169
rect 524255 378135 524265 378169
rect 524303 378135 524323 378169
rect 524323 378135 524337 378169
rect 524375 378135 524391 378169
rect 524391 378135 524409 378169
rect 524447 378135 524459 378169
rect 524459 378135 524481 378169
rect 524519 378135 524527 378169
rect 524527 378135 524553 378169
rect 524591 378135 524595 378169
rect 524595 378135 524625 378169
rect 524663 378135 524697 378169
rect 523439 377677 523473 377711
rect 523511 377677 523541 377711
rect 523541 377677 523545 377711
rect 523583 377677 523609 377711
rect 523609 377677 523617 377711
rect 523655 377677 523677 377711
rect 523677 377677 523689 377711
rect 523727 377677 523745 377711
rect 523745 377677 523761 377711
rect 523799 377677 523813 377711
rect 523813 377677 523833 377711
rect 523871 377677 523881 377711
rect 523881 377677 523905 377711
rect 523943 377677 523949 377711
rect 523949 377677 523977 377711
rect 524015 377677 524017 377711
rect 524017 377677 524049 377711
rect 524087 377677 524119 377711
rect 524119 377677 524121 377711
rect 524159 377677 524187 377711
rect 524187 377677 524193 377711
rect 524231 377677 524255 377711
rect 524255 377677 524265 377711
rect 524303 377677 524323 377711
rect 524323 377677 524337 377711
rect 524375 377677 524391 377711
rect 524391 377677 524409 377711
rect 524447 377677 524459 377711
rect 524459 377677 524481 377711
rect 524519 377677 524527 377711
rect 524527 377677 524553 377711
rect 524591 377677 524595 377711
rect 524595 377677 524625 377711
rect 524663 377677 524697 377711
rect 523171 377107 523205 377141
rect 523171 376707 523205 376741
rect 523171 376307 523205 376341
rect 523439 377219 523473 377253
rect 523511 377219 523541 377253
rect 523541 377219 523545 377253
rect 523583 377219 523609 377253
rect 523609 377219 523617 377253
rect 523655 377219 523677 377253
rect 523677 377219 523689 377253
rect 523727 377219 523745 377253
rect 523745 377219 523761 377253
rect 523799 377219 523813 377253
rect 523813 377219 523833 377253
rect 523871 377219 523881 377253
rect 523881 377219 523905 377253
rect 523943 377219 523949 377253
rect 523949 377219 523977 377253
rect 524015 377219 524017 377253
rect 524017 377219 524049 377253
rect 524087 377219 524119 377253
rect 524119 377219 524121 377253
rect 524159 377219 524187 377253
rect 524187 377219 524193 377253
rect 524231 377219 524255 377253
rect 524255 377219 524265 377253
rect 524303 377219 524323 377253
rect 524323 377219 524337 377253
rect 524375 377219 524391 377253
rect 524391 377219 524409 377253
rect 524447 377219 524459 377253
rect 524459 377219 524481 377253
rect 524519 377219 524527 377253
rect 524527 377219 524553 377253
rect 524591 377219 524595 377253
rect 524595 377219 524625 377253
rect 524663 377219 524697 377253
rect 523439 376761 523473 376795
rect 523511 376761 523541 376795
rect 523541 376761 523545 376795
rect 523583 376761 523609 376795
rect 523609 376761 523617 376795
rect 523655 376761 523677 376795
rect 523677 376761 523689 376795
rect 523727 376761 523745 376795
rect 523745 376761 523761 376795
rect 523799 376761 523813 376795
rect 523813 376761 523833 376795
rect 523871 376761 523881 376795
rect 523881 376761 523905 376795
rect 523943 376761 523949 376795
rect 523949 376761 523977 376795
rect 524015 376761 524017 376795
rect 524017 376761 524049 376795
rect 524087 376761 524119 376795
rect 524119 376761 524121 376795
rect 524159 376761 524187 376795
rect 524187 376761 524193 376795
rect 524231 376761 524255 376795
rect 524255 376761 524265 376795
rect 524303 376761 524323 376795
rect 524323 376761 524337 376795
rect 524375 376761 524391 376795
rect 524391 376761 524409 376795
rect 524447 376761 524459 376795
rect 524459 376761 524481 376795
rect 524519 376761 524527 376795
rect 524527 376761 524553 376795
rect 524591 376761 524595 376795
rect 524595 376761 524625 376795
rect 524663 376761 524697 376795
rect 523171 375907 523205 375941
rect 523171 375507 523205 375541
rect 513771 374865 513805 374899
rect 523171 375107 523205 375141
rect 523439 376303 523473 376337
rect 523511 376303 523541 376337
rect 523541 376303 523545 376337
rect 523583 376303 523609 376337
rect 523609 376303 523617 376337
rect 523655 376303 523677 376337
rect 523677 376303 523689 376337
rect 523727 376303 523745 376337
rect 523745 376303 523761 376337
rect 523799 376303 523813 376337
rect 523813 376303 523833 376337
rect 523871 376303 523881 376337
rect 523881 376303 523905 376337
rect 523943 376303 523949 376337
rect 523949 376303 523977 376337
rect 524015 376303 524017 376337
rect 524017 376303 524049 376337
rect 524087 376303 524119 376337
rect 524119 376303 524121 376337
rect 524159 376303 524187 376337
rect 524187 376303 524193 376337
rect 524231 376303 524255 376337
rect 524255 376303 524265 376337
rect 524303 376303 524323 376337
rect 524323 376303 524337 376337
rect 524375 376303 524391 376337
rect 524391 376303 524409 376337
rect 524447 376303 524459 376337
rect 524459 376303 524481 376337
rect 524519 376303 524527 376337
rect 524527 376303 524553 376337
rect 524591 376303 524595 376337
rect 524595 376303 524625 376337
rect 524663 376303 524697 376337
rect 523439 375845 523473 375879
rect 523511 375845 523541 375879
rect 523541 375845 523545 375879
rect 523583 375845 523609 375879
rect 523609 375845 523617 375879
rect 523655 375845 523677 375879
rect 523677 375845 523689 375879
rect 523727 375845 523745 375879
rect 523745 375845 523761 375879
rect 523799 375845 523813 375879
rect 523813 375845 523833 375879
rect 523871 375845 523881 375879
rect 523881 375845 523905 375879
rect 523943 375845 523949 375879
rect 523949 375845 523977 375879
rect 524015 375845 524017 375879
rect 524017 375845 524049 375879
rect 524087 375845 524119 375879
rect 524119 375845 524121 375879
rect 524159 375845 524187 375879
rect 524187 375845 524193 375879
rect 524231 375845 524255 375879
rect 524255 375845 524265 375879
rect 524303 375845 524323 375879
rect 524323 375845 524337 375879
rect 524375 375845 524391 375879
rect 524391 375845 524409 375879
rect 524447 375845 524459 375879
rect 524459 375845 524481 375879
rect 524519 375845 524527 375879
rect 524527 375845 524553 375879
rect 524591 375845 524595 375879
rect 524595 375845 524625 375879
rect 524663 375845 524697 375879
rect 523439 375387 523473 375421
rect 523511 375387 523541 375421
rect 523541 375387 523545 375421
rect 523583 375387 523609 375421
rect 523609 375387 523617 375421
rect 523655 375387 523677 375421
rect 523677 375387 523689 375421
rect 523727 375387 523745 375421
rect 523745 375387 523761 375421
rect 523799 375387 523813 375421
rect 523813 375387 523833 375421
rect 523871 375387 523881 375421
rect 523881 375387 523905 375421
rect 523943 375387 523949 375421
rect 523949 375387 523977 375421
rect 524015 375387 524017 375421
rect 524017 375387 524049 375421
rect 524087 375387 524119 375421
rect 524119 375387 524121 375421
rect 524159 375387 524187 375421
rect 524187 375387 524193 375421
rect 524231 375387 524255 375421
rect 524255 375387 524265 375421
rect 524303 375387 524323 375421
rect 524323 375387 524337 375421
rect 524375 375387 524391 375421
rect 524391 375387 524409 375421
rect 524447 375387 524459 375421
rect 524459 375387 524481 375421
rect 524519 375387 524527 375421
rect 524527 375387 524553 375421
rect 524591 375387 524595 375421
rect 524595 375387 524625 375421
rect 524663 375387 524697 375421
rect 523439 374929 523473 374963
rect 523511 374929 523541 374963
rect 523541 374929 523545 374963
rect 523583 374929 523609 374963
rect 523609 374929 523617 374963
rect 523655 374929 523677 374963
rect 523677 374929 523689 374963
rect 523727 374929 523745 374963
rect 523745 374929 523761 374963
rect 523799 374929 523813 374963
rect 523813 374929 523833 374963
rect 523871 374929 523881 374963
rect 523881 374929 523905 374963
rect 523943 374929 523949 374963
rect 523949 374929 523977 374963
rect 524015 374929 524017 374963
rect 524017 374929 524049 374963
rect 524087 374929 524119 374963
rect 524119 374929 524121 374963
rect 524159 374929 524187 374963
rect 524187 374929 524193 374963
rect 524231 374929 524255 374963
rect 524255 374929 524265 374963
rect 524303 374929 524323 374963
rect 524323 374929 524337 374963
rect 524375 374929 524391 374963
rect 524391 374929 524409 374963
rect 524447 374929 524459 374963
rect 524459 374929 524481 374963
rect 524519 374929 524527 374963
rect 524527 374929 524553 374963
rect 524591 374929 524595 374963
rect 524595 374929 524625 374963
rect 524663 374929 524697 374963
rect 515651 374599 515685 374633
rect 510011 374285 510045 374319
rect 515651 374399 515685 374433
rect 515919 374403 516457 374797
rect 516879 374403 517417 374797
rect 517531 374599 517565 374633
rect 517531 374399 517565 374433
rect 515651 374199 515685 374233
rect 502491 373861 502525 373895
rect 515651 373999 515685 374033
rect 517531 374199 517565 374233
rect 517531 373999 517565 374033
rect 515651 373799 515685 373833
rect 515651 373599 515685 373633
rect 498731 373307 498765 373341
rect 515651 373399 515685 373433
rect 517531 373799 517565 373833
rect 517531 373599 517565 373633
rect 517531 373399 517565 373433
rect 515651 373199 515685 373233
rect 498731 372907 498765 372941
rect 498731 372507 498765 372541
rect 500611 372953 500645 372987
rect 500611 372753 500645 372787
rect 500611 372553 500645 372587
rect 500611 372353 500645 372387
rect 500611 372153 500645 372187
rect 494971 371907 495005 371941
rect 494971 371507 495005 371541
rect 494971 371107 495005 371141
rect 494971 370707 495005 370741
rect 494971 370307 495005 370341
rect 494971 369907 495005 369941
rect 494971 369507 495005 369541
rect 494971 369107 495005 369141
rect 494971 368707 495005 368741
rect 494971 368307 495005 368341
rect 494971 367907 495005 367941
rect 494971 367507 495005 367541
rect 494971 367107 495005 367141
rect 494971 366707 495005 366741
rect 494971 366307 495005 366341
rect 494971 365907 495005 365941
rect 494971 365507 495005 365541
rect 494971 365107 495005 365141
rect 494971 364707 495005 364741
rect 494971 364307 495005 364341
rect 494971 363907 495005 363941
rect 494971 363507 495005 363541
rect 494971 363107 495005 363141
rect 494971 362707 495005 362741
rect 496851 371777 496885 371811
rect 496851 371577 496885 371611
rect 496851 371377 496885 371411
rect 496851 371177 496885 371211
rect 496851 370977 496885 371011
rect 496851 370777 496885 370811
rect 496851 370577 496885 370611
rect 496851 370377 496885 370411
rect 496851 370177 496885 370211
rect 496851 369977 496885 370011
rect 496851 369777 496885 369811
rect 496851 369577 496885 369611
rect 496851 369377 496885 369411
rect 496851 369177 496885 369211
rect 496851 368977 496885 369011
rect 496851 368777 496885 368811
rect 496851 368577 496885 368611
rect 496851 368377 496885 368411
rect 496851 368177 496885 368211
rect 496851 367977 496885 368011
rect 496851 367777 496885 367811
rect 496851 367577 496885 367611
rect 496851 367377 496885 367411
rect 496851 367177 496885 367211
rect 496851 366977 496885 367011
rect 496851 366777 496885 366811
rect 496851 366577 496885 366611
rect 496851 366377 496885 366411
rect 496851 366177 496885 366211
rect 496851 365977 496885 366011
rect 496851 365777 496885 365811
rect 496851 365577 496885 365611
rect 496851 365377 496885 365411
rect 496851 365177 496885 365211
rect 496851 364977 496885 365011
rect 496851 364777 496885 364811
rect 496851 364577 496885 364611
rect 496851 364377 496885 364411
rect 496851 364177 496885 364211
rect 496851 363977 496885 364011
rect 496851 363777 496885 363811
rect 496851 363577 496885 363611
rect 496851 363377 496885 363411
rect 496851 363177 496885 363211
rect 496851 362977 496885 363011
rect 496851 362777 496885 362811
rect 497184 371914 497218 371948
rect 497184 371838 497218 371858
rect 497184 371824 497199 371838
rect 497199 371824 497218 371838
rect 497184 371748 497218 371768
rect 497184 371734 497199 371748
rect 497199 371734 497218 371748
rect 497184 371658 497218 371678
rect 497184 371644 497199 371658
rect 497199 371644 497218 371658
rect 497184 371568 497218 371588
rect 497184 371554 497199 371568
rect 497199 371554 497218 371568
rect 497184 371478 497218 371498
rect 497184 371464 497199 371478
rect 497199 371464 497218 371478
rect 497184 371388 497218 371408
rect 497184 371374 497199 371388
rect 497199 371374 497218 371388
rect 497184 371298 497218 371318
rect 497184 371284 497199 371298
rect 497199 371284 497218 371298
rect 497184 371208 497218 371228
rect 497184 371194 497199 371208
rect 497199 371194 497218 371208
rect 497184 371118 497218 371138
rect 497184 371104 497199 371118
rect 497199 371104 497218 371118
rect 497184 371028 497218 371048
rect 497184 371014 497199 371028
rect 497199 371014 497218 371028
rect 497184 370938 497218 370958
rect 497184 370924 497199 370938
rect 497199 370924 497218 370938
rect 497184 370848 497218 370868
rect 497184 370834 497199 370848
rect 497199 370834 497218 370848
rect 497344 371750 497378 371784
rect 497344 371674 497378 371694
rect 497344 371660 497346 371674
rect 497346 371660 497378 371674
rect 497344 371584 497378 371604
rect 497344 371570 497346 371584
rect 497346 371570 497378 371584
rect 497344 371494 497378 371514
rect 497344 371480 497346 371494
rect 497346 371480 497378 371494
rect 497344 371404 497378 371424
rect 497344 371390 497346 371404
rect 497346 371390 497378 371404
rect 497344 371314 497378 371334
rect 497344 371300 497346 371314
rect 497346 371300 497378 371314
rect 497344 371224 497378 371244
rect 497344 371210 497346 371224
rect 497346 371210 497378 371224
rect 497344 371134 497378 371154
rect 497344 371120 497346 371134
rect 497346 371120 497378 371134
rect 497344 371044 497378 371064
rect 497344 371030 497346 371044
rect 497346 371030 497378 371044
rect 497548 371576 497554 371598
rect 497554 371576 497582 371598
rect 497548 371564 497582 371576
rect 497648 371564 497682 371598
rect 497748 371564 497782 371598
rect 497848 371576 497880 371598
rect 497880 371576 497882 371598
rect 497948 371576 497970 371598
rect 497970 371576 497982 371598
rect 498048 371576 498060 371598
rect 498060 371576 498082 371598
rect 497848 371564 497882 371576
rect 497948 371564 497982 371576
rect 498048 371564 498082 371576
rect 497548 371486 497554 371498
rect 497554 371486 497582 371498
rect 497548 371464 497582 371486
rect 497648 371464 497682 371498
rect 497748 371464 497782 371498
rect 497848 371486 497880 371498
rect 497880 371486 497882 371498
rect 497948 371486 497970 371498
rect 497970 371486 497982 371498
rect 498048 371486 498060 371498
rect 498060 371486 498082 371498
rect 497848 371464 497882 371486
rect 497948 371464 497982 371486
rect 498048 371464 498082 371486
rect 497548 371396 497554 371398
rect 497554 371396 497582 371398
rect 497548 371364 497582 371396
rect 497648 371364 497682 371398
rect 497748 371364 497782 371398
rect 497848 371396 497880 371398
rect 497880 371396 497882 371398
rect 497948 371396 497970 371398
rect 497970 371396 497982 371398
rect 498048 371396 498060 371398
rect 498060 371396 498082 371398
rect 497848 371364 497882 371396
rect 497948 371364 497982 371396
rect 498048 371364 498082 371396
rect 497548 371264 497582 371298
rect 497648 371264 497682 371298
rect 497748 371264 497782 371298
rect 497848 371264 497882 371298
rect 497948 371264 497982 371298
rect 498048 371264 498082 371298
rect 497548 371164 497582 371198
rect 497648 371164 497682 371198
rect 497748 371164 497782 371198
rect 497848 371164 497882 371198
rect 497948 371164 497982 371198
rect 498048 371164 498082 371198
rect 497548 371070 497582 371098
rect 497548 371064 497554 371070
rect 497554 371064 497582 371070
rect 497648 371064 497682 371098
rect 497748 371064 497782 371098
rect 497848 371070 497882 371098
rect 497948 371070 497982 371098
rect 498048 371070 498082 371098
rect 497848 371064 497880 371070
rect 497880 371064 497882 371070
rect 497948 371064 497970 371070
rect 497970 371064 497982 371070
rect 498048 371064 498060 371070
rect 498060 371064 498082 371070
rect 497344 370954 497378 370974
rect 497344 370940 497346 370954
rect 497346 370940 497378 370954
rect 497344 370850 497378 370884
rect 497184 370744 497218 370778
rect 497184 370574 497218 370608
rect 497184 370498 497218 370518
rect 497184 370484 497199 370498
rect 497199 370484 497218 370498
rect 497184 370408 497218 370428
rect 497184 370394 497199 370408
rect 497199 370394 497218 370408
rect 497184 370318 497218 370338
rect 497184 370304 497199 370318
rect 497199 370304 497218 370318
rect 497184 370228 497218 370248
rect 497184 370214 497199 370228
rect 497199 370214 497218 370228
rect 497184 370138 497218 370158
rect 497184 370124 497199 370138
rect 497199 370124 497218 370138
rect 497184 370048 497218 370068
rect 497184 370034 497199 370048
rect 497199 370034 497218 370048
rect 497184 369958 497218 369978
rect 497184 369944 497199 369958
rect 497199 369944 497218 369958
rect 497184 369868 497218 369888
rect 497184 369854 497199 369868
rect 497199 369854 497218 369868
rect 497184 369778 497218 369798
rect 497184 369764 497199 369778
rect 497199 369764 497218 369778
rect 497184 369688 497218 369708
rect 497184 369674 497199 369688
rect 497199 369674 497218 369688
rect 497184 369598 497218 369618
rect 497184 369584 497199 369598
rect 497199 369584 497218 369598
rect 497184 369508 497218 369528
rect 497184 369494 497199 369508
rect 497199 369494 497218 369508
rect 497344 370410 497378 370444
rect 497344 370334 497378 370354
rect 497344 370320 497346 370334
rect 497346 370320 497378 370334
rect 497344 370244 497378 370264
rect 497344 370230 497346 370244
rect 497346 370230 497378 370244
rect 497344 370154 497378 370174
rect 497344 370140 497346 370154
rect 497346 370140 497378 370154
rect 497344 370064 497378 370084
rect 497344 370050 497346 370064
rect 497346 370050 497378 370064
rect 497344 369974 497378 369994
rect 497344 369960 497346 369974
rect 497346 369960 497378 369974
rect 497344 369884 497378 369904
rect 497344 369870 497346 369884
rect 497346 369870 497378 369884
rect 497344 369794 497378 369814
rect 497344 369780 497346 369794
rect 497346 369780 497378 369794
rect 497344 369704 497378 369724
rect 497344 369690 497346 369704
rect 497346 369690 497378 369704
rect 497548 370236 497554 370258
rect 497554 370236 497582 370258
rect 497548 370224 497582 370236
rect 497648 370224 497682 370258
rect 497748 370224 497782 370258
rect 497848 370236 497880 370258
rect 497880 370236 497882 370258
rect 497948 370236 497970 370258
rect 497970 370236 497982 370258
rect 498048 370236 498060 370258
rect 498060 370236 498082 370258
rect 497848 370224 497882 370236
rect 497948 370224 497982 370236
rect 498048 370224 498082 370236
rect 497548 370146 497554 370158
rect 497554 370146 497582 370158
rect 497548 370124 497582 370146
rect 497648 370124 497682 370158
rect 497748 370124 497782 370158
rect 497848 370146 497880 370158
rect 497880 370146 497882 370158
rect 497948 370146 497970 370158
rect 497970 370146 497982 370158
rect 498048 370146 498060 370158
rect 498060 370146 498082 370158
rect 497848 370124 497882 370146
rect 497948 370124 497982 370146
rect 498048 370124 498082 370146
rect 497548 370056 497554 370058
rect 497554 370056 497582 370058
rect 497548 370024 497582 370056
rect 497648 370024 497682 370058
rect 497748 370024 497782 370058
rect 497848 370056 497880 370058
rect 497880 370056 497882 370058
rect 497948 370056 497970 370058
rect 497970 370056 497982 370058
rect 498048 370056 498060 370058
rect 498060 370056 498082 370058
rect 497848 370024 497882 370056
rect 497948 370024 497982 370056
rect 498048 370024 498082 370056
rect 497548 369924 497582 369958
rect 497648 369924 497682 369958
rect 497748 369924 497782 369958
rect 497848 369924 497882 369958
rect 497948 369924 497982 369958
rect 498048 369924 498082 369958
rect 497548 369824 497582 369858
rect 497648 369824 497682 369858
rect 497748 369824 497782 369858
rect 497848 369824 497882 369858
rect 497948 369824 497982 369858
rect 498048 369824 498082 369858
rect 497548 369730 497582 369758
rect 497548 369724 497554 369730
rect 497554 369724 497582 369730
rect 497648 369724 497682 369758
rect 497748 369724 497782 369758
rect 497848 369730 497882 369758
rect 497948 369730 497982 369758
rect 498048 369730 498082 369758
rect 497848 369724 497880 369730
rect 497880 369724 497882 369730
rect 497948 369724 497970 369730
rect 497970 369724 497982 369730
rect 498048 369724 498060 369730
rect 498060 369724 498082 369730
rect 497344 369614 497378 369634
rect 497344 369600 497346 369614
rect 497346 369600 497378 369614
rect 497344 369510 497378 369544
rect 497184 369404 497218 369438
rect 497184 369234 497218 369268
rect 497184 369158 497218 369178
rect 497184 369144 497199 369158
rect 497199 369144 497218 369158
rect 497184 369068 497218 369088
rect 497184 369054 497199 369068
rect 497199 369054 497218 369068
rect 497184 368978 497218 368998
rect 497184 368964 497199 368978
rect 497199 368964 497218 368978
rect 497184 368888 497218 368908
rect 497184 368874 497199 368888
rect 497199 368874 497218 368888
rect 497184 368798 497218 368818
rect 497184 368784 497199 368798
rect 497199 368784 497218 368798
rect 497184 368708 497218 368728
rect 497184 368694 497199 368708
rect 497199 368694 497218 368708
rect 497184 368618 497218 368638
rect 497184 368604 497199 368618
rect 497199 368604 497218 368618
rect 497184 368528 497218 368548
rect 497184 368514 497199 368528
rect 497199 368514 497218 368528
rect 497184 368438 497218 368458
rect 497184 368424 497199 368438
rect 497199 368424 497218 368438
rect 497184 368348 497218 368368
rect 497184 368334 497199 368348
rect 497199 368334 497218 368348
rect 497184 368258 497218 368278
rect 497184 368244 497199 368258
rect 497199 368244 497218 368258
rect 497184 368168 497218 368188
rect 497184 368154 497199 368168
rect 497199 368154 497218 368168
rect 497344 369070 497378 369104
rect 497344 368994 497378 369014
rect 497344 368980 497346 368994
rect 497346 368980 497378 368994
rect 497344 368904 497378 368924
rect 497344 368890 497346 368904
rect 497346 368890 497378 368904
rect 497344 368814 497378 368834
rect 497344 368800 497346 368814
rect 497346 368800 497378 368814
rect 497344 368724 497378 368744
rect 497344 368710 497346 368724
rect 497346 368710 497378 368724
rect 497344 368634 497378 368654
rect 497344 368620 497346 368634
rect 497346 368620 497378 368634
rect 497344 368544 497378 368564
rect 497344 368530 497346 368544
rect 497346 368530 497378 368544
rect 497344 368454 497378 368474
rect 497344 368440 497346 368454
rect 497346 368440 497378 368454
rect 497344 368364 497378 368384
rect 497344 368350 497346 368364
rect 497346 368350 497378 368364
rect 497548 368896 497554 368918
rect 497554 368896 497582 368918
rect 497548 368884 497582 368896
rect 497648 368884 497682 368918
rect 497748 368884 497782 368918
rect 497848 368896 497880 368918
rect 497880 368896 497882 368918
rect 497948 368896 497970 368918
rect 497970 368896 497982 368918
rect 498048 368896 498060 368918
rect 498060 368896 498082 368918
rect 497848 368884 497882 368896
rect 497948 368884 497982 368896
rect 498048 368884 498082 368896
rect 497548 368806 497554 368818
rect 497554 368806 497582 368818
rect 497548 368784 497582 368806
rect 497648 368784 497682 368818
rect 497748 368784 497782 368818
rect 497848 368806 497880 368818
rect 497880 368806 497882 368818
rect 497948 368806 497970 368818
rect 497970 368806 497982 368818
rect 498048 368806 498060 368818
rect 498060 368806 498082 368818
rect 497848 368784 497882 368806
rect 497948 368784 497982 368806
rect 498048 368784 498082 368806
rect 497548 368716 497554 368718
rect 497554 368716 497582 368718
rect 497548 368684 497582 368716
rect 497648 368684 497682 368718
rect 497748 368684 497782 368718
rect 497848 368716 497880 368718
rect 497880 368716 497882 368718
rect 497948 368716 497970 368718
rect 497970 368716 497982 368718
rect 498048 368716 498060 368718
rect 498060 368716 498082 368718
rect 497848 368684 497882 368716
rect 497948 368684 497982 368716
rect 498048 368684 498082 368716
rect 497548 368584 497582 368618
rect 497648 368584 497682 368618
rect 497748 368584 497782 368618
rect 497848 368584 497882 368618
rect 497948 368584 497982 368618
rect 498048 368584 498082 368618
rect 497548 368484 497582 368518
rect 497648 368484 497682 368518
rect 497748 368484 497782 368518
rect 497848 368484 497882 368518
rect 497948 368484 497982 368518
rect 498048 368484 498082 368518
rect 497548 368390 497582 368418
rect 497548 368384 497554 368390
rect 497554 368384 497582 368390
rect 497648 368384 497682 368418
rect 497748 368384 497782 368418
rect 497848 368390 497882 368418
rect 497948 368390 497982 368418
rect 498048 368390 498082 368418
rect 497848 368384 497880 368390
rect 497880 368384 497882 368390
rect 497948 368384 497970 368390
rect 497970 368384 497982 368390
rect 498048 368384 498060 368390
rect 498060 368384 498082 368390
rect 497344 368274 497378 368294
rect 497344 368260 497346 368274
rect 497346 368260 497378 368274
rect 497344 368170 497378 368204
rect 497184 368064 497218 368098
rect 497184 367894 497218 367928
rect 497184 367818 497218 367838
rect 497184 367804 497199 367818
rect 497199 367804 497218 367818
rect 497184 367728 497218 367748
rect 497184 367714 497199 367728
rect 497199 367714 497218 367728
rect 497184 367638 497218 367658
rect 497184 367624 497199 367638
rect 497199 367624 497218 367638
rect 497184 367548 497218 367568
rect 497184 367534 497199 367548
rect 497199 367534 497218 367548
rect 497184 367458 497218 367478
rect 497184 367444 497199 367458
rect 497199 367444 497218 367458
rect 497184 367368 497218 367388
rect 497184 367354 497199 367368
rect 497199 367354 497218 367368
rect 497184 367278 497218 367298
rect 497184 367264 497199 367278
rect 497199 367264 497218 367278
rect 497184 367188 497218 367208
rect 497184 367174 497199 367188
rect 497199 367174 497218 367188
rect 497184 367098 497218 367118
rect 497184 367084 497199 367098
rect 497199 367084 497218 367098
rect 497184 367008 497218 367028
rect 497184 366994 497199 367008
rect 497199 366994 497218 367008
rect 497184 366918 497218 366938
rect 497184 366904 497199 366918
rect 497199 366904 497218 366918
rect 497184 366828 497218 366848
rect 497184 366814 497199 366828
rect 497199 366814 497218 366828
rect 497344 367730 497378 367764
rect 497344 367654 497378 367674
rect 497344 367640 497346 367654
rect 497346 367640 497378 367654
rect 497344 367564 497378 367584
rect 497344 367550 497346 367564
rect 497346 367550 497378 367564
rect 497344 367474 497378 367494
rect 497344 367460 497346 367474
rect 497346 367460 497378 367474
rect 497344 367384 497378 367404
rect 497344 367370 497346 367384
rect 497346 367370 497378 367384
rect 497344 367294 497378 367314
rect 497344 367280 497346 367294
rect 497346 367280 497378 367294
rect 497344 367204 497378 367224
rect 497344 367190 497346 367204
rect 497346 367190 497378 367204
rect 497344 367114 497378 367134
rect 497344 367100 497346 367114
rect 497346 367100 497378 367114
rect 497344 367024 497378 367044
rect 497344 367010 497346 367024
rect 497346 367010 497378 367024
rect 497548 367556 497554 367578
rect 497554 367556 497582 367578
rect 497548 367544 497582 367556
rect 497648 367544 497682 367578
rect 497748 367544 497782 367578
rect 497848 367556 497880 367578
rect 497880 367556 497882 367578
rect 497948 367556 497970 367578
rect 497970 367556 497982 367578
rect 498048 367556 498060 367578
rect 498060 367556 498082 367578
rect 497848 367544 497882 367556
rect 497948 367544 497982 367556
rect 498048 367544 498082 367556
rect 497548 367466 497554 367478
rect 497554 367466 497582 367478
rect 497548 367444 497582 367466
rect 497648 367444 497682 367478
rect 497748 367444 497782 367478
rect 497848 367466 497880 367478
rect 497880 367466 497882 367478
rect 497948 367466 497970 367478
rect 497970 367466 497982 367478
rect 498048 367466 498060 367478
rect 498060 367466 498082 367478
rect 497848 367444 497882 367466
rect 497948 367444 497982 367466
rect 498048 367444 498082 367466
rect 497548 367376 497554 367378
rect 497554 367376 497582 367378
rect 497548 367344 497582 367376
rect 497648 367344 497682 367378
rect 497748 367344 497782 367378
rect 497848 367376 497880 367378
rect 497880 367376 497882 367378
rect 497948 367376 497970 367378
rect 497970 367376 497982 367378
rect 498048 367376 498060 367378
rect 498060 367376 498082 367378
rect 497848 367344 497882 367376
rect 497948 367344 497982 367376
rect 498048 367344 498082 367376
rect 497548 367244 497582 367278
rect 497648 367244 497682 367278
rect 497748 367244 497782 367278
rect 497848 367244 497882 367278
rect 497948 367244 497982 367278
rect 498048 367244 498082 367278
rect 497548 367144 497582 367178
rect 497648 367144 497682 367178
rect 497748 367144 497782 367178
rect 497848 367144 497882 367178
rect 497948 367144 497982 367178
rect 498048 367144 498082 367178
rect 497548 367050 497582 367078
rect 497548 367044 497554 367050
rect 497554 367044 497582 367050
rect 497648 367044 497682 367078
rect 497748 367044 497782 367078
rect 497848 367050 497882 367078
rect 497948 367050 497982 367078
rect 498048 367050 498082 367078
rect 497848 367044 497880 367050
rect 497880 367044 497882 367050
rect 497948 367044 497970 367050
rect 497970 367044 497982 367050
rect 498048 367044 498060 367050
rect 498060 367044 498082 367050
rect 497344 366934 497378 366954
rect 497344 366920 497346 366934
rect 497346 366920 497378 366934
rect 497344 366830 497378 366864
rect 497184 366724 497218 366758
rect 497184 366554 497218 366588
rect 497184 366478 497218 366498
rect 497184 366464 497199 366478
rect 497199 366464 497218 366478
rect 497184 366388 497218 366408
rect 497184 366374 497199 366388
rect 497199 366374 497218 366388
rect 497184 366298 497218 366318
rect 497184 366284 497199 366298
rect 497199 366284 497218 366298
rect 497184 366208 497218 366228
rect 497184 366194 497199 366208
rect 497199 366194 497218 366208
rect 497184 366118 497218 366138
rect 497184 366104 497199 366118
rect 497199 366104 497218 366118
rect 497184 366028 497218 366048
rect 497184 366014 497199 366028
rect 497199 366014 497218 366028
rect 497184 365938 497218 365958
rect 497184 365924 497199 365938
rect 497199 365924 497218 365938
rect 497184 365848 497218 365868
rect 497184 365834 497199 365848
rect 497199 365834 497218 365848
rect 497184 365758 497218 365778
rect 497184 365744 497199 365758
rect 497199 365744 497218 365758
rect 497184 365668 497218 365688
rect 497184 365654 497199 365668
rect 497199 365654 497218 365668
rect 497184 365578 497218 365598
rect 497184 365564 497199 365578
rect 497199 365564 497218 365578
rect 497184 365488 497218 365508
rect 497184 365474 497199 365488
rect 497199 365474 497218 365488
rect 497344 366390 497378 366424
rect 497344 366314 497378 366334
rect 497344 366300 497346 366314
rect 497346 366300 497378 366314
rect 497344 366224 497378 366244
rect 497344 366210 497346 366224
rect 497346 366210 497378 366224
rect 497344 366134 497378 366154
rect 497344 366120 497346 366134
rect 497346 366120 497378 366134
rect 497344 366044 497378 366064
rect 497344 366030 497346 366044
rect 497346 366030 497378 366044
rect 497344 365954 497378 365974
rect 497344 365940 497346 365954
rect 497346 365940 497378 365954
rect 497344 365864 497378 365884
rect 497344 365850 497346 365864
rect 497346 365850 497378 365864
rect 497344 365774 497378 365794
rect 497344 365760 497346 365774
rect 497346 365760 497378 365774
rect 497344 365684 497378 365704
rect 497344 365670 497346 365684
rect 497346 365670 497378 365684
rect 497548 366216 497554 366238
rect 497554 366216 497582 366238
rect 497548 366204 497582 366216
rect 497648 366204 497682 366238
rect 497748 366204 497782 366238
rect 497848 366216 497880 366238
rect 497880 366216 497882 366238
rect 497948 366216 497970 366238
rect 497970 366216 497982 366238
rect 498048 366216 498060 366238
rect 498060 366216 498082 366238
rect 497848 366204 497882 366216
rect 497948 366204 497982 366216
rect 498048 366204 498082 366216
rect 497548 366126 497554 366138
rect 497554 366126 497582 366138
rect 497548 366104 497582 366126
rect 497648 366104 497682 366138
rect 497748 366104 497782 366138
rect 497848 366126 497880 366138
rect 497880 366126 497882 366138
rect 497948 366126 497970 366138
rect 497970 366126 497982 366138
rect 498048 366126 498060 366138
rect 498060 366126 498082 366138
rect 497848 366104 497882 366126
rect 497948 366104 497982 366126
rect 498048 366104 498082 366126
rect 497548 366036 497554 366038
rect 497554 366036 497582 366038
rect 497548 366004 497582 366036
rect 497648 366004 497682 366038
rect 497748 366004 497782 366038
rect 497848 366036 497880 366038
rect 497880 366036 497882 366038
rect 497948 366036 497970 366038
rect 497970 366036 497982 366038
rect 498048 366036 498060 366038
rect 498060 366036 498082 366038
rect 497848 366004 497882 366036
rect 497948 366004 497982 366036
rect 498048 366004 498082 366036
rect 497548 365904 497582 365938
rect 497648 365904 497682 365938
rect 497748 365904 497782 365938
rect 497848 365904 497882 365938
rect 497948 365904 497982 365938
rect 498048 365904 498082 365938
rect 497548 365804 497582 365838
rect 497648 365804 497682 365838
rect 497748 365804 497782 365838
rect 497848 365804 497882 365838
rect 497948 365804 497982 365838
rect 498048 365804 498082 365838
rect 497548 365710 497582 365738
rect 497548 365704 497554 365710
rect 497554 365704 497582 365710
rect 497648 365704 497682 365738
rect 497748 365704 497782 365738
rect 497848 365710 497882 365738
rect 497948 365710 497982 365738
rect 498048 365710 498082 365738
rect 497848 365704 497880 365710
rect 497880 365704 497882 365710
rect 497948 365704 497970 365710
rect 497970 365704 497982 365710
rect 498048 365704 498060 365710
rect 498060 365704 498082 365710
rect 497344 365594 497378 365614
rect 497344 365580 497346 365594
rect 497346 365580 497378 365594
rect 497344 365490 497378 365524
rect 497184 365384 497218 365418
rect 497184 365214 497218 365248
rect 497184 365138 497218 365158
rect 497184 365124 497199 365138
rect 497199 365124 497218 365138
rect 497184 365048 497218 365068
rect 497184 365034 497199 365048
rect 497199 365034 497218 365048
rect 497184 364958 497218 364978
rect 497184 364944 497199 364958
rect 497199 364944 497218 364958
rect 497184 364868 497218 364888
rect 497184 364854 497199 364868
rect 497199 364854 497218 364868
rect 497184 364778 497218 364798
rect 497184 364764 497199 364778
rect 497199 364764 497218 364778
rect 497184 364688 497218 364708
rect 497184 364674 497199 364688
rect 497199 364674 497218 364688
rect 497184 364598 497218 364618
rect 497184 364584 497199 364598
rect 497199 364584 497218 364598
rect 497184 364508 497218 364528
rect 497184 364494 497199 364508
rect 497199 364494 497218 364508
rect 497184 364418 497218 364438
rect 497184 364404 497199 364418
rect 497199 364404 497218 364418
rect 497184 364328 497218 364348
rect 497184 364314 497199 364328
rect 497199 364314 497218 364328
rect 497184 364238 497218 364258
rect 497184 364224 497199 364238
rect 497199 364224 497218 364238
rect 497184 364148 497218 364168
rect 497184 364134 497199 364148
rect 497199 364134 497218 364148
rect 497344 365050 497378 365084
rect 497344 364974 497378 364994
rect 497344 364960 497346 364974
rect 497346 364960 497378 364974
rect 497344 364884 497378 364904
rect 497344 364870 497346 364884
rect 497346 364870 497378 364884
rect 497344 364794 497378 364814
rect 497344 364780 497346 364794
rect 497346 364780 497378 364794
rect 497344 364704 497378 364724
rect 497344 364690 497346 364704
rect 497346 364690 497378 364704
rect 497344 364614 497378 364634
rect 497344 364600 497346 364614
rect 497346 364600 497378 364614
rect 497344 364524 497378 364544
rect 497344 364510 497346 364524
rect 497346 364510 497378 364524
rect 497344 364434 497378 364454
rect 497344 364420 497346 364434
rect 497346 364420 497378 364434
rect 497344 364344 497378 364364
rect 497344 364330 497346 364344
rect 497346 364330 497378 364344
rect 497548 364876 497554 364898
rect 497554 364876 497582 364898
rect 497548 364864 497582 364876
rect 497648 364864 497682 364898
rect 497748 364864 497782 364898
rect 497848 364876 497880 364898
rect 497880 364876 497882 364898
rect 497948 364876 497970 364898
rect 497970 364876 497982 364898
rect 498048 364876 498060 364898
rect 498060 364876 498082 364898
rect 497848 364864 497882 364876
rect 497948 364864 497982 364876
rect 498048 364864 498082 364876
rect 497548 364786 497554 364798
rect 497554 364786 497582 364798
rect 497548 364764 497582 364786
rect 497648 364764 497682 364798
rect 497748 364764 497782 364798
rect 497848 364786 497880 364798
rect 497880 364786 497882 364798
rect 497948 364786 497970 364798
rect 497970 364786 497982 364798
rect 498048 364786 498060 364798
rect 498060 364786 498082 364798
rect 497848 364764 497882 364786
rect 497948 364764 497982 364786
rect 498048 364764 498082 364786
rect 497548 364696 497554 364698
rect 497554 364696 497582 364698
rect 497548 364664 497582 364696
rect 497648 364664 497682 364698
rect 497748 364664 497782 364698
rect 497848 364696 497880 364698
rect 497880 364696 497882 364698
rect 497948 364696 497970 364698
rect 497970 364696 497982 364698
rect 498048 364696 498060 364698
rect 498060 364696 498082 364698
rect 497848 364664 497882 364696
rect 497948 364664 497982 364696
rect 498048 364664 498082 364696
rect 497548 364564 497582 364598
rect 497648 364564 497682 364598
rect 497748 364564 497782 364598
rect 497848 364564 497882 364598
rect 497948 364564 497982 364598
rect 498048 364564 498082 364598
rect 497548 364464 497582 364498
rect 497648 364464 497682 364498
rect 497748 364464 497782 364498
rect 497848 364464 497882 364498
rect 497948 364464 497982 364498
rect 498048 364464 498082 364498
rect 497548 364370 497582 364398
rect 497548 364364 497554 364370
rect 497554 364364 497582 364370
rect 497648 364364 497682 364398
rect 497748 364364 497782 364398
rect 497848 364370 497882 364398
rect 497948 364370 497982 364398
rect 498048 364370 498082 364398
rect 497848 364364 497880 364370
rect 497880 364364 497882 364370
rect 497948 364364 497970 364370
rect 497970 364364 497982 364370
rect 498048 364364 498060 364370
rect 498060 364364 498082 364370
rect 497344 364254 497378 364274
rect 497344 364240 497346 364254
rect 497346 364240 497378 364254
rect 497344 364150 497378 364184
rect 497184 364044 497218 364078
rect 497184 363874 497218 363908
rect 497184 363798 497218 363818
rect 497184 363784 497199 363798
rect 497199 363784 497218 363798
rect 497184 363708 497218 363728
rect 497184 363694 497199 363708
rect 497199 363694 497218 363708
rect 497184 363618 497218 363638
rect 497184 363604 497199 363618
rect 497199 363604 497218 363618
rect 497184 363528 497218 363548
rect 497184 363514 497199 363528
rect 497199 363514 497218 363528
rect 497184 363438 497218 363458
rect 497184 363424 497199 363438
rect 497199 363424 497218 363438
rect 497184 363348 497218 363368
rect 497184 363334 497199 363348
rect 497199 363334 497218 363348
rect 497184 363258 497218 363278
rect 497184 363244 497199 363258
rect 497199 363244 497218 363258
rect 497184 363168 497218 363188
rect 497184 363154 497199 363168
rect 497199 363154 497218 363168
rect 497184 363078 497218 363098
rect 497184 363064 497199 363078
rect 497199 363064 497218 363078
rect 497184 362988 497218 363008
rect 497184 362974 497199 362988
rect 497199 362974 497218 362988
rect 497184 362898 497218 362918
rect 497184 362884 497199 362898
rect 497199 362884 497218 362898
rect 497184 362808 497218 362828
rect 497184 362794 497199 362808
rect 497199 362794 497218 362808
rect 497344 363710 497378 363744
rect 497344 363634 497378 363654
rect 497344 363620 497346 363634
rect 497346 363620 497378 363634
rect 497344 363544 497378 363564
rect 497344 363530 497346 363544
rect 497346 363530 497378 363544
rect 497344 363454 497378 363474
rect 497344 363440 497346 363454
rect 497346 363440 497378 363454
rect 497344 363364 497378 363384
rect 497344 363350 497346 363364
rect 497346 363350 497378 363364
rect 497344 363274 497378 363294
rect 497344 363260 497346 363274
rect 497346 363260 497378 363274
rect 497344 363184 497378 363204
rect 497344 363170 497346 363184
rect 497346 363170 497378 363184
rect 497344 363094 497378 363114
rect 497344 363080 497346 363094
rect 497346 363080 497378 363094
rect 497344 363004 497378 363024
rect 497344 362990 497346 363004
rect 497346 362990 497378 363004
rect 497548 363536 497554 363558
rect 497554 363536 497582 363558
rect 497548 363524 497582 363536
rect 497648 363524 497682 363558
rect 497748 363524 497782 363558
rect 497848 363536 497880 363558
rect 497880 363536 497882 363558
rect 497948 363536 497970 363558
rect 497970 363536 497982 363558
rect 498048 363536 498060 363558
rect 498060 363536 498082 363558
rect 497848 363524 497882 363536
rect 497948 363524 497982 363536
rect 498048 363524 498082 363536
rect 497548 363446 497554 363458
rect 497554 363446 497582 363458
rect 497548 363424 497582 363446
rect 497648 363424 497682 363458
rect 497748 363424 497782 363458
rect 497848 363446 497880 363458
rect 497880 363446 497882 363458
rect 497948 363446 497970 363458
rect 497970 363446 497982 363458
rect 498048 363446 498060 363458
rect 498060 363446 498082 363458
rect 497848 363424 497882 363446
rect 497948 363424 497982 363446
rect 498048 363424 498082 363446
rect 497548 363356 497554 363358
rect 497554 363356 497582 363358
rect 497548 363324 497582 363356
rect 497648 363324 497682 363358
rect 497748 363324 497782 363358
rect 497848 363356 497880 363358
rect 497880 363356 497882 363358
rect 497948 363356 497970 363358
rect 497970 363356 497982 363358
rect 498048 363356 498060 363358
rect 498060 363356 498082 363358
rect 497848 363324 497882 363356
rect 497948 363324 497982 363356
rect 498048 363324 498082 363356
rect 497548 363224 497582 363258
rect 497648 363224 497682 363258
rect 497748 363224 497782 363258
rect 497848 363224 497882 363258
rect 497948 363224 497982 363258
rect 498048 363224 498082 363258
rect 497548 363124 497582 363158
rect 497648 363124 497682 363158
rect 497748 363124 497782 363158
rect 497848 363124 497882 363158
rect 497948 363124 497982 363158
rect 498048 363124 498082 363158
rect 497548 363030 497582 363058
rect 497548 363024 497554 363030
rect 497554 363024 497582 363030
rect 497648 363024 497682 363058
rect 497748 363024 497782 363058
rect 497848 363030 497882 363058
rect 497948 363030 497982 363058
rect 498048 363030 498082 363058
rect 497848 363024 497880 363030
rect 497880 363024 497882 363030
rect 497948 363024 497970 363030
rect 497970 363024 497982 363030
rect 498048 363024 498060 363030
rect 498060 363024 498082 363030
rect 497344 362914 497378 362934
rect 497344 362900 497346 362914
rect 497346 362900 497378 362914
rect 497344 362810 497378 362844
rect 497184 362704 497218 362738
rect 498731 371777 498765 371811
rect 498731 371577 498765 371611
rect 498731 371377 498765 371411
rect 498731 371177 498765 371211
rect 498731 370977 498765 371011
rect 498731 370777 498765 370811
rect 498731 370577 498765 370611
rect 498731 370377 498765 370411
rect 498731 370177 498765 370211
rect 498731 369977 498765 370011
rect 498731 369777 498765 369811
rect 498731 369577 498765 369611
rect 498731 369377 498765 369411
rect 498731 369177 498765 369211
rect 498731 368977 498765 369011
rect 498731 368777 498765 368811
rect 498731 368577 498765 368611
rect 498731 368377 498765 368411
rect 498731 368177 498765 368211
rect 498731 367977 498765 368011
rect 498731 367777 498765 367811
rect 498731 367577 498765 367611
rect 498731 367377 498765 367411
rect 498731 367177 498765 367211
rect 498731 366977 498765 367011
rect 498731 366777 498765 366811
rect 498731 366577 498765 366611
rect 498731 366377 498765 366411
rect 498731 366177 498765 366211
rect 498731 365977 498765 366011
rect 498731 365777 498765 365811
rect 498731 365577 498765 365611
rect 498731 365377 498765 365411
rect 498731 365177 498765 365211
rect 498731 364977 498765 365011
rect 498731 364777 498765 364811
rect 498731 364577 498765 364611
rect 498731 364377 498765 364411
rect 498731 364177 498765 364211
rect 498731 363977 498765 364011
rect 498731 363777 498765 363811
rect 498731 363577 498765 363611
rect 498731 363377 498765 363411
rect 498731 363177 498765 363211
rect 498731 362977 498765 363011
rect 498731 362777 498765 362811
rect 500611 371953 500645 371987
rect 500611 371753 500645 371787
rect 500611 371553 500645 371587
rect 500611 371353 500645 371387
rect 500611 371153 500645 371187
rect 500611 370953 500645 370987
rect 500611 370753 500645 370787
rect 500611 370553 500645 370587
rect 500611 370353 500645 370387
rect 500611 370153 500645 370187
rect 500611 369953 500645 369987
rect 500611 369753 500645 369787
rect 500611 369553 500645 369587
rect 500611 369353 500645 369387
rect 500611 369153 500645 369187
rect 500611 368953 500645 368987
rect 500611 368753 500645 368787
rect 500611 368553 500645 368587
rect 500611 368353 500645 368387
rect 500611 368153 500645 368187
rect 500611 367953 500645 367987
rect 500611 367753 500645 367787
rect 500611 367553 500645 367587
rect 500611 367353 500645 367387
rect 500611 367153 500645 367187
rect 500611 366953 500645 366987
rect 500611 366753 500645 366787
rect 500611 366553 500645 366587
rect 500611 366353 500645 366387
rect 500611 366153 500645 366187
rect 500611 365953 500645 365987
rect 500611 365753 500645 365787
rect 500611 365553 500645 365587
rect 500611 365353 500645 365387
rect 500611 365153 500645 365187
rect 500611 364953 500645 364987
rect 500611 364753 500645 364787
rect 500611 364553 500645 364587
rect 500611 364353 500645 364387
rect 500611 364153 500645 364187
rect 500611 363953 500645 363987
rect 500611 363753 500645 363787
rect 500611 363553 500645 363587
rect 500611 363353 500645 363387
rect 500611 363153 500645 363187
rect 500611 362953 500645 362987
rect 500611 362753 500645 362787
rect 500611 362553 500645 362587
rect 500944 373090 500978 373124
rect 500944 373014 500978 373034
rect 500944 373000 500959 373014
rect 500959 373000 500978 373014
rect 500944 372924 500978 372944
rect 500944 372910 500959 372924
rect 500959 372910 500978 372924
rect 500944 372834 500978 372854
rect 500944 372820 500959 372834
rect 500959 372820 500978 372834
rect 500944 372744 500978 372764
rect 500944 372730 500959 372744
rect 500959 372730 500978 372744
rect 500944 372654 500978 372674
rect 500944 372640 500959 372654
rect 500959 372640 500978 372654
rect 500944 372564 500978 372584
rect 500944 372550 500959 372564
rect 500959 372550 500978 372564
rect 500944 372474 500978 372494
rect 500944 372460 500959 372474
rect 500959 372460 500978 372474
rect 500944 372384 500978 372404
rect 500944 372370 500959 372384
rect 500959 372370 500978 372384
rect 500944 372294 500978 372314
rect 500944 372280 500959 372294
rect 500959 372280 500978 372294
rect 500944 372204 500978 372224
rect 500944 372190 500959 372204
rect 500959 372190 500978 372204
rect 500944 372114 500978 372134
rect 500944 372100 500959 372114
rect 500959 372100 500978 372114
rect 500944 372024 500978 372044
rect 500944 372010 500959 372024
rect 500959 372010 500978 372024
rect 501104 372926 501138 372960
rect 501104 372850 501138 372870
rect 501104 372836 501106 372850
rect 501106 372836 501138 372850
rect 501104 372760 501138 372780
rect 501104 372746 501106 372760
rect 501106 372746 501138 372760
rect 501104 372670 501138 372690
rect 501104 372656 501106 372670
rect 501106 372656 501138 372670
rect 501104 372580 501138 372600
rect 501104 372566 501106 372580
rect 501106 372566 501138 372580
rect 501104 372490 501138 372510
rect 501104 372476 501106 372490
rect 501106 372476 501138 372490
rect 501104 372400 501138 372420
rect 501104 372386 501106 372400
rect 501106 372386 501138 372400
rect 501104 372310 501138 372330
rect 501104 372296 501106 372310
rect 501106 372296 501138 372310
rect 501104 372220 501138 372240
rect 501104 372206 501106 372220
rect 501106 372206 501138 372220
rect 501308 372752 501314 372774
rect 501314 372752 501342 372774
rect 501308 372740 501342 372752
rect 501408 372740 501442 372774
rect 501508 372740 501542 372774
rect 501608 372752 501640 372774
rect 501640 372752 501642 372774
rect 501708 372752 501730 372774
rect 501730 372752 501742 372774
rect 501808 372752 501820 372774
rect 501820 372752 501842 372774
rect 501608 372740 501642 372752
rect 501708 372740 501742 372752
rect 501808 372740 501842 372752
rect 501308 372662 501314 372674
rect 501314 372662 501342 372674
rect 501308 372640 501342 372662
rect 501408 372640 501442 372674
rect 501508 372640 501542 372674
rect 501608 372662 501640 372674
rect 501640 372662 501642 372674
rect 501708 372662 501730 372674
rect 501730 372662 501742 372674
rect 501808 372662 501820 372674
rect 501820 372662 501842 372674
rect 501608 372640 501642 372662
rect 501708 372640 501742 372662
rect 501808 372640 501842 372662
rect 501308 372572 501314 372574
rect 501314 372572 501342 372574
rect 501308 372540 501342 372572
rect 501408 372540 501442 372574
rect 501508 372540 501542 372574
rect 501608 372572 501640 372574
rect 501640 372572 501642 372574
rect 501708 372572 501730 372574
rect 501730 372572 501742 372574
rect 501808 372572 501820 372574
rect 501820 372572 501842 372574
rect 501608 372540 501642 372572
rect 501708 372540 501742 372572
rect 501808 372540 501842 372572
rect 501308 372440 501342 372474
rect 501408 372440 501442 372474
rect 501508 372440 501542 372474
rect 501608 372440 501642 372474
rect 501708 372440 501742 372474
rect 501808 372440 501842 372474
rect 501308 372340 501342 372374
rect 501408 372340 501442 372374
rect 501508 372340 501542 372374
rect 501608 372340 501642 372374
rect 501708 372340 501742 372374
rect 501808 372340 501842 372374
rect 501308 372246 501342 372274
rect 501308 372240 501314 372246
rect 501314 372240 501342 372246
rect 501408 372240 501442 372274
rect 501508 372240 501542 372274
rect 501608 372246 501642 372274
rect 501708 372246 501742 372274
rect 501808 372246 501842 372274
rect 501608 372240 501640 372246
rect 501640 372240 501642 372246
rect 501708 372240 501730 372246
rect 501730 372240 501742 372246
rect 501808 372240 501820 372246
rect 501820 372240 501842 372246
rect 501104 372130 501138 372150
rect 501104 372116 501106 372130
rect 501106 372116 501138 372130
rect 501104 372026 501138 372060
rect 500944 371920 500978 371954
rect 500944 371750 500978 371784
rect 500944 371674 500978 371694
rect 500944 371660 500959 371674
rect 500959 371660 500978 371674
rect 500944 371584 500978 371604
rect 500944 371570 500959 371584
rect 500959 371570 500978 371584
rect 500944 371494 500978 371514
rect 500944 371480 500959 371494
rect 500959 371480 500978 371494
rect 500944 371404 500978 371424
rect 500944 371390 500959 371404
rect 500959 371390 500978 371404
rect 500944 371314 500978 371334
rect 500944 371300 500959 371314
rect 500959 371300 500978 371314
rect 500944 371224 500978 371244
rect 500944 371210 500959 371224
rect 500959 371210 500978 371224
rect 500944 371134 500978 371154
rect 500944 371120 500959 371134
rect 500959 371120 500978 371134
rect 500944 371044 500978 371064
rect 500944 371030 500959 371044
rect 500959 371030 500978 371044
rect 500944 370954 500978 370974
rect 500944 370940 500959 370954
rect 500959 370940 500978 370954
rect 500944 370864 500978 370884
rect 500944 370850 500959 370864
rect 500959 370850 500978 370864
rect 500944 370774 500978 370794
rect 500944 370760 500959 370774
rect 500959 370760 500978 370774
rect 500944 370684 500978 370704
rect 500944 370670 500959 370684
rect 500959 370670 500978 370684
rect 501104 371586 501138 371620
rect 501104 371510 501138 371530
rect 501104 371496 501106 371510
rect 501106 371496 501138 371510
rect 501104 371420 501138 371440
rect 501104 371406 501106 371420
rect 501106 371406 501138 371420
rect 501104 371330 501138 371350
rect 501104 371316 501106 371330
rect 501106 371316 501138 371330
rect 501104 371240 501138 371260
rect 501104 371226 501106 371240
rect 501106 371226 501138 371240
rect 501104 371150 501138 371170
rect 501104 371136 501106 371150
rect 501106 371136 501138 371150
rect 501104 371060 501138 371080
rect 501104 371046 501106 371060
rect 501106 371046 501138 371060
rect 501104 370970 501138 370990
rect 501104 370956 501106 370970
rect 501106 370956 501138 370970
rect 501104 370880 501138 370900
rect 501104 370866 501106 370880
rect 501106 370866 501138 370880
rect 501308 371412 501314 371434
rect 501314 371412 501342 371434
rect 501308 371400 501342 371412
rect 501408 371400 501442 371434
rect 501508 371400 501542 371434
rect 501608 371412 501640 371434
rect 501640 371412 501642 371434
rect 501708 371412 501730 371434
rect 501730 371412 501742 371434
rect 501808 371412 501820 371434
rect 501820 371412 501842 371434
rect 501608 371400 501642 371412
rect 501708 371400 501742 371412
rect 501808 371400 501842 371412
rect 501308 371322 501314 371334
rect 501314 371322 501342 371334
rect 501308 371300 501342 371322
rect 501408 371300 501442 371334
rect 501508 371300 501542 371334
rect 501608 371322 501640 371334
rect 501640 371322 501642 371334
rect 501708 371322 501730 371334
rect 501730 371322 501742 371334
rect 501808 371322 501820 371334
rect 501820 371322 501842 371334
rect 501608 371300 501642 371322
rect 501708 371300 501742 371322
rect 501808 371300 501842 371322
rect 501308 371232 501314 371234
rect 501314 371232 501342 371234
rect 501308 371200 501342 371232
rect 501408 371200 501442 371234
rect 501508 371200 501542 371234
rect 501608 371232 501640 371234
rect 501640 371232 501642 371234
rect 501708 371232 501730 371234
rect 501730 371232 501742 371234
rect 501808 371232 501820 371234
rect 501820 371232 501842 371234
rect 501608 371200 501642 371232
rect 501708 371200 501742 371232
rect 501808 371200 501842 371232
rect 501308 371100 501342 371134
rect 501408 371100 501442 371134
rect 501508 371100 501542 371134
rect 501608 371100 501642 371134
rect 501708 371100 501742 371134
rect 501808 371100 501842 371134
rect 501308 371000 501342 371034
rect 501408 371000 501442 371034
rect 501508 371000 501542 371034
rect 501608 371000 501642 371034
rect 501708 371000 501742 371034
rect 501808 371000 501842 371034
rect 501308 370906 501342 370934
rect 501308 370900 501314 370906
rect 501314 370900 501342 370906
rect 501408 370900 501442 370934
rect 501508 370900 501542 370934
rect 501608 370906 501642 370934
rect 501708 370906 501742 370934
rect 501808 370906 501842 370934
rect 501608 370900 501640 370906
rect 501640 370900 501642 370906
rect 501708 370900 501730 370906
rect 501730 370900 501742 370906
rect 501808 370900 501820 370906
rect 501820 370900 501842 370906
rect 501104 370790 501138 370810
rect 501104 370776 501106 370790
rect 501106 370776 501138 370790
rect 501104 370686 501138 370720
rect 500944 370580 500978 370614
rect 500944 370410 500978 370444
rect 500944 370334 500978 370354
rect 500944 370320 500959 370334
rect 500959 370320 500978 370334
rect 500944 370244 500978 370264
rect 500944 370230 500959 370244
rect 500959 370230 500978 370244
rect 500944 370154 500978 370174
rect 500944 370140 500959 370154
rect 500959 370140 500978 370154
rect 500944 370064 500978 370084
rect 500944 370050 500959 370064
rect 500959 370050 500978 370064
rect 500944 369974 500978 369994
rect 500944 369960 500959 369974
rect 500959 369960 500978 369974
rect 500944 369884 500978 369904
rect 500944 369870 500959 369884
rect 500959 369870 500978 369884
rect 500944 369794 500978 369814
rect 500944 369780 500959 369794
rect 500959 369780 500978 369794
rect 500944 369704 500978 369724
rect 500944 369690 500959 369704
rect 500959 369690 500978 369704
rect 500944 369614 500978 369634
rect 500944 369600 500959 369614
rect 500959 369600 500978 369614
rect 500944 369524 500978 369544
rect 500944 369510 500959 369524
rect 500959 369510 500978 369524
rect 500944 369434 500978 369454
rect 500944 369420 500959 369434
rect 500959 369420 500978 369434
rect 500944 369344 500978 369364
rect 500944 369330 500959 369344
rect 500959 369330 500978 369344
rect 501104 370246 501138 370280
rect 501104 370170 501138 370190
rect 501104 370156 501106 370170
rect 501106 370156 501138 370170
rect 501104 370080 501138 370100
rect 501104 370066 501106 370080
rect 501106 370066 501138 370080
rect 501104 369990 501138 370010
rect 501104 369976 501106 369990
rect 501106 369976 501138 369990
rect 501104 369900 501138 369920
rect 501104 369886 501106 369900
rect 501106 369886 501138 369900
rect 501104 369810 501138 369830
rect 501104 369796 501106 369810
rect 501106 369796 501138 369810
rect 501104 369720 501138 369740
rect 501104 369706 501106 369720
rect 501106 369706 501138 369720
rect 501104 369630 501138 369650
rect 501104 369616 501106 369630
rect 501106 369616 501138 369630
rect 501104 369540 501138 369560
rect 501104 369526 501106 369540
rect 501106 369526 501138 369540
rect 501308 370072 501314 370094
rect 501314 370072 501342 370094
rect 501308 370060 501342 370072
rect 501408 370060 501442 370094
rect 501508 370060 501542 370094
rect 501608 370072 501640 370094
rect 501640 370072 501642 370094
rect 501708 370072 501730 370094
rect 501730 370072 501742 370094
rect 501808 370072 501820 370094
rect 501820 370072 501842 370094
rect 501608 370060 501642 370072
rect 501708 370060 501742 370072
rect 501808 370060 501842 370072
rect 501308 369982 501314 369994
rect 501314 369982 501342 369994
rect 501308 369960 501342 369982
rect 501408 369960 501442 369994
rect 501508 369960 501542 369994
rect 501608 369982 501640 369994
rect 501640 369982 501642 369994
rect 501708 369982 501730 369994
rect 501730 369982 501742 369994
rect 501808 369982 501820 369994
rect 501820 369982 501842 369994
rect 501608 369960 501642 369982
rect 501708 369960 501742 369982
rect 501808 369960 501842 369982
rect 501308 369892 501314 369894
rect 501314 369892 501342 369894
rect 501308 369860 501342 369892
rect 501408 369860 501442 369894
rect 501508 369860 501542 369894
rect 501608 369892 501640 369894
rect 501640 369892 501642 369894
rect 501708 369892 501730 369894
rect 501730 369892 501742 369894
rect 501808 369892 501820 369894
rect 501820 369892 501842 369894
rect 501608 369860 501642 369892
rect 501708 369860 501742 369892
rect 501808 369860 501842 369892
rect 501308 369760 501342 369794
rect 501408 369760 501442 369794
rect 501508 369760 501542 369794
rect 501608 369760 501642 369794
rect 501708 369760 501742 369794
rect 501808 369760 501842 369794
rect 501308 369660 501342 369694
rect 501408 369660 501442 369694
rect 501508 369660 501542 369694
rect 501608 369660 501642 369694
rect 501708 369660 501742 369694
rect 501808 369660 501842 369694
rect 501308 369566 501342 369594
rect 501308 369560 501314 369566
rect 501314 369560 501342 369566
rect 501408 369560 501442 369594
rect 501508 369560 501542 369594
rect 501608 369566 501642 369594
rect 501708 369566 501742 369594
rect 501808 369566 501842 369594
rect 501608 369560 501640 369566
rect 501640 369560 501642 369566
rect 501708 369560 501730 369566
rect 501730 369560 501742 369566
rect 501808 369560 501820 369566
rect 501820 369560 501842 369566
rect 501104 369450 501138 369470
rect 501104 369436 501106 369450
rect 501106 369436 501138 369450
rect 501104 369346 501138 369380
rect 500944 369240 500978 369274
rect 500944 369070 500978 369104
rect 500944 368994 500978 369014
rect 500944 368980 500959 368994
rect 500959 368980 500978 368994
rect 500944 368904 500978 368924
rect 500944 368890 500959 368904
rect 500959 368890 500978 368904
rect 500944 368814 500978 368834
rect 500944 368800 500959 368814
rect 500959 368800 500978 368814
rect 500944 368724 500978 368744
rect 500944 368710 500959 368724
rect 500959 368710 500978 368724
rect 500944 368634 500978 368654
rect 500944 368620 500959 368634
rect 500959 368620 500978 368634
rect 500944 368544 500978 368564
rect 500944 368530 500959 368544
rect 500959 368530 500978 368544
rect 500944 368454 500978 368474
rect 500944 368440 500959 368454
rect 500959 368440 500978 368454
rect 500944 368364 500978 368384
rect 500944 368350 500959 368364
rect 500959 368350 500978 368364
rect 500944 368274 500978 368294
rect 500944 368260 500959 368274
rect 500959 368260 500978 368274
rect 500944 368184 500978 368204
rect 500944 368170 500959 368184
rect 500959 368170 500978 368184
rect 500944 368094 500978 368114
rect 500944 368080 500959 368094
rect 500959 368080 500978 368094
rect 500944 368004 500978 368024
rect 500944 367990 500959 368004
rect 500959 367990 500978 368004
rect 501104 368906 501138 368940
rect 501104 368830 501138 368850
rect 501104 368816 501106 368830
rect 501106 368816 501138 368830
rect 501104 368740 501138 368760
rect 501104 368726 501106 368740
rect 501106 368726 501138 368740
rect 501104 368650 501138 368670
rect 501104 368636 501106 368650
rect 501106 368636 501138 368650
rect 501104 368560 501138 368580
rect 501104 368546 501106 368560
rect 501106 368546 501138 368560
rect 501104 368470 501138 368490
rect 501104 368456 501106 368470
rect 501106 368456 501138 368470
rect 501104 368380 501138 368400
rect 501104 368366 501106 368380
rect 501106 368366 501138 368380
rect 501104 368290 501138 368310
rect 501104 368276 501106 368290
rect 501106 368276 501138 368290
rect 501104 368200 501138 368220
rect 501104 368186 501106 368200
rect 501106 368186 501138 368200
rect 501308 368732 501314 368754
rect 501314 368732 501342 368754
rect 501308 368720 501342 368732
rect 501408 368720 501442 368754
rect 501508 368720 501542 368754
rect 501608 368732 501640 368754
rect 501640 368732 501642 368754
rect 501708 368732 501730 368754
rect 501730 368732 501742 368754
rect 501808 368732 501820 368754
rect 501820 368732 501842 368754
rect 501608 368720 501642 368732
rect 501708 368720 501742 368732
rect 501808 368720 501842 368732
rect 501308 368642 501314 368654
rect 501314 368642 501342 368654
rect 501308 368620 501342 368642
rect 501408 368620 501442 368654
rect 501508 368620 501542 368654
rect 501608 368642 501640 368654
rect 501640 368642 501642 368654
rect 501708 368642 501730 368654
rect 501730 368642 501742 368654
rect 501808 368642 501820 368654
rect 501820 368642 501842 368654
rect 501608 368620 501642 368642
rect 501708 368620 501742 368642
rect 501808 368620 501842 368642
rect 501308 368552 501314 368554
rect 501314 368552 501342 368554
rect 501308 368520 501342 368552
rect 501408 368520 501442 368554
rect 501508 368520 501542 368554
rect 501608 368552 501640 368554
rect 501640 368552 501642 368554
rect 501708 368552 501730 368554
rect 501730 368552 501742 368554
rect 501808 368552 501820 368554
rect 501820 368552 501842 368554
rect 501608 368520 501642 368552
rect 501708 368520 501742 368552
rect 501808 368520 501842 368552
rect 501308 368420 501342 368454
rect 501408 368420 501442 368454
rect 501508 368420 501542 368454
rect 501608 368420 501642 368454
rect 501708 368420 501742 368454
rect 501808 368420 501842 368454
rect 501308 368320 501342 368354
rect 501408 368320 501442 368354
rect 501508 368320 501542 368354
rect 501608 368320 501642 368354
rect 501708 368320 501742 368354
rect 501808 368320 501842 368354
rect 501308 368226 501342 368254
rect 501308 368220 501314 368226
rect 501314 368220 501342 368226
rect 501408 368220 501442 368254
rect 501508 368220 501542 368254
rect 501608 368226 501642 368254
rect 501708 368226 501742 368254
rect 501808 368226 501842 368254
rect 501608 368220 501640 368226
rect 501640 368220 501642 368226
rect 501708 368220 501730 368226
rect 501730 368220 501742 368226
rect 501808 368220 501820 368226
rect 501820 368220 501842 368226
rect 501104 368110 501138 368130
rect 501104 368096 501106 368110
rect 501106 368096 501138 368110
rect 501104 368006 501138 368040
rect 500944 367900 500978 367934
rect 500944 367730 500978 367764
rect 500944 367654 500978 367674
rect 500944 367640 500959 367654
rect 500959 367640 500978 367654
rect 500944 367564 500978 367584
rect 500944 367550 500959 367564
rect 500959 367550 500978 367564
rect 500944 367474 500978 367494
rect 500944 367460 500959 367474
rect 500959 367460 500978 367474
rect 500944 367384 500978 367404
rect 500944 367370 500959 367384
rect 500959 367370 500978 367384
rect 500944 367294 500978 367314
rect 500944 367280 500959 367294
rect 500959 367280 500978 367294
rect 500944 367204 500978 367224
rect 500944 367190 500959 367204
rect 500959 367190 500978 367204
rect 500944 367114 500978 367134
rect 500944 367100 500959 367114
rect 500959 367100 500978 367114
rect 500944 367024 500978 367044
rect 500944 367010 500959 367024
rect 500959 367010 500978 367024
rect 500944 366934 500978 366954
rect 500944 366920 500959 366934
rect 500959 366920 500978 366934
rect 500944 366844 500978 366864
rect 500944 366830 500959 366844
rect 500959 366830 500978 366844
rect 500944 366754 500978 366774
rect 500944 366740 500959 366754
rect 500959 366740 500978 366754
rect 500944 366664 500978 366684
rect 500944 366650 500959 366664
rect 500959 366650 500978 366664
rect 501104 367566 501138 367600
rect 501104 367490 501138 367510
rect 501104 367476 501106 367490
rect 501106 367476 501138 367490
rect 501104 367400 501138 367420
rect 501104 367386 501106 367400
rect 501106 367386 501138 367400
rect 501104 367310 501138 367330
rect 501104 367296 501106 367310
rect 501106 367296 501138 367310
rect 501104 367220 501138 367240
rect 501104 367206 501106 367220
rect 501106 367206 501138 367220
rect 501104 367130 501138 367150
rect 501104 367116 501106 367130
rect 501106 367116 501138 367130
rect 501104 367040 501138 367060
rect 501104 367026 501106 367040
rect 501106 367026 501138 367040
rect 501104 366950 501138 366970
rect 501104 366936 501106 366950
rect 501106 366936 501138 366950
rect 501104 366860 501138 366880
rect 501104 366846 501106 366860
rect 501106 366846 501138 366860
rect 501308 367392 501314 367414
rect 501314 367392 501342 367414
rect 501308 367380 501342 367392
rect 501408 367380 501442 367414
rect 501508 367380 501542 367414
rect 501608 367392 501640 367414
rect 501640 367392 501642 367414
rect 501708 367392 501730 367414
rect 501730 367392 501742 367414
rect 501808 367392 501820 367414
rect 501820 367392 501842 367414
rect 501608 367380 501642 367392
rect 501708 367380 501742 367392
rect 501808 367380 501842 367392
rect 501308 367302 501314 367314
rect 501314 367302 501342 367314
rect 501308 367280 501342 367302
rect 501408 367280 501442 367314
rect 501508 367280 501542 367314
rect 501608 367302 501640 367314
rect 501640 367302 501642 367314
rect 501708 367302 501730 367314
rect 501730 367302 501742 367314
rect 501808 367302 501820 367314
rect 501820 367302 501842 367314
rect 501608 367280 501642 367302
rect 501708 367280 501742 367302
rect 501808 367280 501842 367302
rect 501308 367212 501314 367214
rect 501314 367212 501342 367214
rect 501308 367180 501342 367212
rect 501408 367180 501442 367214
rect 501508 367180 501542 367214
rect 501608 367212 501640 367214
rect 501640 367212 501642 367214
rect 501708 367212 501730 367214
rect 501730 367212 501742 367214
rect 501808 367212 501820 367214
rect 501820 367212 501842 367214
rect 501608 367180 501642 367212
rect 501708 367180 501742 367212
rect 501808 367180 501842 367212
rect 501308 367080 501342 367114
rect 501408 367080 501442 367114
rect 501508 367080 501542 367114
rect 501608 367080 501642 367114
rect 501708 367080 501742 367114
rect 501808 367080 501842 367114
rect 501308 366980 501342 367014
rect 501408 366980 501442 367014
rect 501508 366980 501542 367014
rect 501608 366980 501642 367014
rect 501708 366980 501742 367014
rect 501808 366980 501842 367014
rect 501308 366886 501342 366914
rect 501308 366880 501314 366886
rect 501314 366880 501342 366886
rect 501408 366880 501442 366914
rect 501508 366880 501542 366914
rect 501608 366886 501642 366914
rect 501708 366886 501742 366914
rect 501808 366886 501842 366914
rect 501608 366880 501640 366886
rect 501640 366880 501642 366886
rect 501708 366880 501730 366886
rect 501730 366880 501742 366886
rect 501808 366880 501820 366886
rect 501820 366880 501842 366886
rect 501104 366770 501138 366790
rect 501104 366756 501106 366770
rect 501106 366756 501138 366770
rect 501104 366666 501138 366700
rect 500944 366560 500978 366594
rect 500944 366390 500978 366424
rect 500944 366314 500978 366334
rect 500944 366300 500959 366314
rect 500959 366300 500978 366314
rect 500944 366224 500978 366244
rect 500944 366210 500959 366224
rect 500959 366210 500978 366224
rect 500944 366134 500978 366154
rect 500944 366120 500959 366134
rect 500959 366120 500978 366134
rect 500944 366044 500978 366064
rect 500944 366030 500959 366044
rect 500959 366030 500978 366044
rect 500944 365954 500978 365974
rect 500944 365940 500959 365954
rect 500959 365940 500978 365954
rect 500944 365864 500978 365884
rect 500944 365850 500959 365864
rect 500959 365850 500978 365864
rect 500944 365774 500978 365794
rect 500944 365760 500959 365774
rect 500959 365760 500978 365774
rect 500944 365684 500978 365704
rect 500944 365670 500959 365684
rect 500959 365670 500978 365684
rect 500944 365594 500978 365614
rect 500944 365580 500959 365594
rect 500959 365580 500978 365594
rect 500944 365504 500978 365524
rect 500944 365490 500959 365504
rect 500959 365490 500978 365504
rect 500944 365414 500978 365434
rect 500944 365400 500959 365414
rect 500959 365400 500978 365414
rect 500944 365324 500978 365344
rect 500944 365310 500959 365324
rect 500959 365310 500978 365324
rect 501104 366226 501138 366260
rect 501104 366150 501138 366170
rect 501104 366136 501106 366150
rect 501106 366136 501138 366150
rect 501104 366060 501138 366080
rect 501104 366046 501106 366060
rect 501106 366046 501138 366060
rect 501104 365970 501138 365990
rect 501104 365956 501106 365970
rect 501106 365956 501138 365970
rect 501104 365880 501138 365900
rect 501104 365866 501106 365880
rect 501106 365866 501138 365880
rect 501104 365790 501138 365810
rect 501104 365776 501106 365790
rect 501106 365776 501138 365790
rect 501104 365700 501138 365720
rect 501104 365686 501106 365700
rect 501106 365686 501138 365700
rect 501104 365610 501138 365630
rect 501104 365596 501106 365610
rect 501106 365596 501138 365610
rect 501104 365520 501138 365540
rect 501104 365506 501106 365520
rect 501106 365506 501138 365520
rect 501308 366052 501314 366074
rect 501314 366052 501342 366074
rect 501308 366040 501342 366052
rect 501408 366040 501442 366074
rect 501508 366040 501542 366074
rect 501608 366052 501640 366074
rect 501640 366052 501642 366074
rect 501708 366052 501730 366074
rect 501730 366052 501742 366074
rect 501808 366052 501820 366074
rect 501820 366052 501842 366074
rect 501608 366040 501642 366052
rect 501708 366040 501742 366052
rect 501808 366040 501842 366052
rect 501308 365962 501314 365974
rect 501314 365962 501342 365974
rect 501308 365940 501342 365962
rect 501408 365940 501442 365974
rect 501508 365940 501542 365974
rect 501608 365962 501640 365974
rect 501640 365962 501642 365974
rect 501708 365962 501730 365974
rect 501730 365962 501742 365974
rect 501808 365962 501820 365974
rect 501820 365962 501842 365974
rect 501608 365940 501642 365962
rect 501708 365940 501742 365962
rect 501808 365940 501842 365962
rect 501308 365872 501314 365874
rect 501314 365872 501342 365874
rect 501308 365840 501342 365872
rect 501408 365840 501442 365874
rect 501508 365840 501542 365874
rect 501608 365872 501640 365874
rect 501640 365872 501642 365874
rect 501708 365872 501730 365874
rect 501730 365872 501742 365874
rect 501808 365872 501820 365874
rect 501820 365872 501842 365874
rect 501608 365840 501642 365872
rect 501708 365840 501742 365872
rect 501808 365840 501842 365872
rect 501308 365740 501342 365774
rect 501408 365740 501442 365774
rect 501508 365740 501542 365774
rect 501608 365740 501642 365774
rect 501708 365740 501742 365774
rect 501808 365740 501842 365774
rect 501308 365640 501342 365674
rect 501408 365640 501442 365674
rect 501508 365640 501542 365674
rect 501608 365640 501642 365674
rect 501708 365640 501742 365674
rect 501808 365640 501842 365674
rect 501308 365546 501342 365574
rect 501308 365540 501314 365546
rect 501314 365540 501342 365546
rect 501408 365540 501442 365574
rect 501508 365540 501542 365574
rect 501608 365546 501642 365574
rect 501708 365546 501742 365574
rect 501808 365546 501842 365574
rect 501608 365540 501640 365546
rect 501640 365540 501642 365546
rect 501708 365540 501730 365546
rect 501730 365540 501742 365546
rect 501808 365540 501820 365546
rect 501820 365540 501842 365546
rect 501104 365430 501138 365450
rect 501104 365416 501106 365430
rect 501106 365416 501138 365430
rect 501104 365326 501138 365360
rect 500944 365220 500978 365254
rect 500944 365050 500978 365084
rect 500944 364974 500978 364994
rect 500944 364960 500959 364974
rect 500959 364960 500978 364974
rect 500944 364884 500978 364904
rect 500944 364870 500959 364884
rect 500959 364870 500978 364884
rect 500944 364794 500978 364814
rect 500944 364780 500959 364794
rect 500959 364780 500978 364794
rect 500944 364704 500978 364724
rect 500944 364690 500959 364704
rect 500959 364690 500978 364704
rect 500944 364614 500978 364634
rect 500944 364600 500959 364614
rect 500959 364600 500978 364614
rect 500944 364524 500978 364544
rect 500944 364510 500959 364524
rect 500959 364510 500978 364524
rect 500944 364434 500978 364454
rect 500944 364420 500959 364434
rect 500959 364420 500978 364434
rect 500944 364344 500978 364364
rect 500944 364330 500959 364344
rect 500959 364330 500978 364344
rect 500944 364254 500978 364274
rect 500944 364240 500959 364254
rect 500959 364240 500978 364254
rect 500944 364164 500978 364184
rect 500944 364150 500959 364164
rect 500959 364150 500978 364164
rect 500944 364074 500978 364094
rect 500944 364060 500959 364074
rect 500959 364060 500978 364074
rect 500944 363984 500978 364004
rect 500944 363970 500959 363984
rect 500959 363970 500978 363984
rect 501104 364886 501138 364920
rect 501104 364810 501138 364830
rect 501104 364796 501106 364810
rect 501106 364796 501138 364810
rect 501104 364720 501138 364740
rect 501104 364706 501106 364720
rect 501106 364706 501138 364720
rect 501104 364630 501138 364650
rect 501104 364616 501106 364630
rect 501106 364616 501138 364630
rect 501104 364540 501138 364560
rect 501104 364526 501106 364540
rect 501106 364526 501138 364540
rect 501104 364450 501138 364470
rect 501104 364436 501106 364450
rect 501106 364436 501138 364450
rect 501104 364360 501138 364380
rect 501104 364346 501106 364360
rect 501106 364346 501138 364360
rect 501104 364270 501138 364290
rect 501104 364256 501106 364270
rect 501106 364256 501138 364270
rect 501104 364180 501138 364200
rect 501104 364166 501106 364180
rect 501106 364166 501138 364180
rect 501308 364712 501314 364734
rect 501314 364712 501342 364734
rect 501308 364700 501342 364712
rect 501408 364700 501442 364734
rect 501508 364700 501542 364734
rect 501608 364712 501640 364734
rect 501640 364712 501642 364734
rect 501708 364712 501730 364734
rect 501730 364712 501742 364734
rect 501808 364712 501820 364734
rect 501820 364712 501842 364734
rect 501608 364700 501642 364712
rect 501708 364700 501742 364712
rect 501808 364700 501842 364712
rect 501308 364622 501314 364634
rect 501314 364622 501342 364634
rect 501308 364600 501342 364622
rect 501408 364600 501442 364634
rect 501508 364600 501542 364634
rect 501608 364622 501640 364634
rect 501640 364622 501642 364634
rect 501708 364622 501730 364634
rect 501730 364622 501742 364634
rect 501808 364622 501820 364634
rect 501820 364622 501842 364634
rect 501608 364600 501642 364622
rect 501708 364600 501742 364622
rect 501808 364600 501842 364622
rect 501308 364532 501314 364534
rect 501314 364532 501342 364534
rect 501308 364500 501342 364532
rect 501408 364500 501442 364534
rect 501508 364500 501542 364534
rect 501608 364532 501640 364534
rect 501640 364532 501642 364534
rect 501708 364532 501730 364534
rect 501730 364532 501742 364534
rect 501808 364532 501820 364534
rect 501820 364532 501842 364534
rect 501608 364500 501642 364532
rect 501708 364500 501742 364532
rect 501808 364500 501842 364532
rect 501308 364400 501342 364434
rect 501408 364400 501442 364434
rect 501508 364400 501542 364434
rect 501608 364400 501642 364434
rect 501708 364400 501742 364434
rect 501808 364400 501842 364434
rect 501308 364300 501342 364334
rect 501408 364300 501442 364334
rect 501508 364300 501542 364334
rect 501608 364300 501642 364334
rect 501708 364300 501742 364334
rect 501808 364300 501842 364334
rect 501308 364206 501342 364234
rect 501308 364200 501314 364206
rect 501314 364200 501342 364206
rect 501408 364200 501442 364234
rect 501508 364200 501542 364234
rect 501608 364206 501642 364234
rect 501708 364206 501742 364234
rect 501808 364206 501842 364234
rect 501608 364200 501640 364206
rect 501640 364200 501642 364206
rect 501708 364200 501730 364206
rect 501730 364200 501742 364206
rect 501808 364200 501820 364206
rect 501820 364200 501842 364206
rect 501104 364090 501138 364110
rect 501104 364076 501106 364090
rect 501106 364076 501138 364090
rect 501104 363986 501138 364020
rect 500944 363880 500978 363914
rect 500944 363710 500978 363744
rect 500944 363634 500978 363654
rect 500944 363620 500959 363634
rect 500959 363620 500978 363634
rect 500944 363544 500978 363564
rect 500944 363530 500959 363544
rect 500959 363530 500978 363544
rect 500944 363454 500978 363474
rect 500944 363440 500959 363454
rect 500959 363440 500978 363454
rect 500944 363364 500978 363384
rect 500944 363350 500959 363364
rect 500959 363350 500978 363364
rect 500944 363274 500978 363294
rect 500944 363260 500959 363274
rect 500959 363260 500978 363274
rect 500944 363184 500978 363204
rect 500944 363170 500959 363184
rect 500959 363170 500978 363184
rect 500944 363094 500978 363114
rect 500944 363080 500959 363094
rect 500959 363080 500978 363094
rect 500944 363004 500978 363024
rect 500944 362990 500959 363004
rect 500959 362990 500978 363004
rect 500944 362914 500978 362934
rect 500944 362900 500959 362914
rect 500959 362900 500978 362914
rect 500944 362824 500978 362844
rect 500944 362810 500959 362824
rect 500959 362810 500978 362824
rect 500944 362734 500978 362754
rect 500944 362720 500959 362734
rect 500959 362720 500978 362734
rect 500944 362644 500978 362664
rect 500944 362630 500959 362644
rect 500959 362630 500978 362644
rect 501104 363546 501138 363580
rect 501104 363470 501138 363490
rect 501104 363456 501106 363470
rect 501106 363456 501138 363470
rect 501104 363380 501138 363400
rect 501104 363366 501106 363380
rect 501106 363366 501138 363380
rect 501104 363290 501138 363310
rect 501104 363276 501106 363290
rect 501106 363276 501138 363290
rect 501104 363200 501138 363220
rect 501104 363186 501106 363200
rect 501106 363186 501138 363200
rect 501104 363110 501138 363130
rect 501104 363096 501106 363110
rect 501106 363096 501138 363110
rect 501104 363020 501138 363040
rect 501104 363006 501106 363020
rect 501106 363006 501138 363020
rect 501104 362930 501138 362950
rect 501104 362916 501106 362930
rect 501106 362916 501138 362930
rect 501104 362840 501138 362860
rect 501104 362826 501106 362840
rect 501106 362826 501138 362840
rect 501308 363372 501314 363394
rect 501314 363372 501342 363394
rect 501308 363360 501342 363372
rect 501408 363360 501442 363394
rect 501508 363360 501542 363394
rect 501608 363372 501640 363394
rect 501640 363372 501642 363394
rect 501708 363372 501730 363394
rect 501730 363372 501742 363394
rect 501808 363372 501820 363394
rect 501820 363372 501842 363394
rect 501608 363360 501642 363372
rect 501708 363360 501742 363372
rect 501808 363360 501842 363372
rect 501308 363282 501314 363294
rect 501314 363282 501342 363294
rect 501308 363260 501342 363282
rect 501408 363260 501442 363294
rect 501508 363260 501542 363294
rect 501608 363282 501640 363294
rect 501640 363282 501642 363294
rect 501708 363282 501730 363294
rect 501730 363282 501742 363294
rect 501808 363282 501820 363294
rect 501820 363282 501842 363294
rect 501608 363260 501642 363282
rect 501708 363260 501742 363282
rect 501808 363260 501842 363282
rect 501308 363192 501314 363194
rect 501314 363192 501342 363194
rect 501308 363160 501342 363192
rect 501408 363160 501442 363194
rect 501508 363160 501542 363194
rect 501608 363192 501640 363194
rect 501640 363192 501642 363194
rect 501708 363192 501730 363194
rect 501730 363192 501742 363194
rect 501808 363192 501820 363194
rect 501820 363192 501842 363194
rect 501608 363160 501642 363192
rect 501708 363160 501742 363192
rect 501808 363160 501842 363192
rect 501308 363060 501342 363094
rect 501408 363060 501442 363094
rect 501508 363060 501542 363094
rect 501608 363060 501642 363094
rect 501708 363060 501742 363094
rect 501808 363060 501842 363094
rect 501308 362960 501342 362994
rect 501408 362960 501442 362994
rect 501508 362960 501542 362994
rect 501608 362960 501642 362994
rect 501708 362960 501742 362994
rect 501808 362960 501842 362994
rect 501308 362866 501342 362894
rect 501308 362860 501314 362866
rect 501314 362860 501342 362866
rect 501408 362860 501442 362894
rect 501508 362860 501542 362894
rect 501608 362866 501642 362894
rect 501708 362866 501742 362894
rect 501808 362866 501842 362894
rect 501608 362860 501640 362866
rect 501640 362860 501642 362866
rect 501708 362860 501730 362866
rect 501730 362860 501742 362866
rect 501808 362860 501820 362866
rect 501820 362860 501842 362866
rect 501104 362750 501138 362770
rect 501104 362736 501106 362750
rect 501106 362736 501138 362750
rect 501104 362646 501138 362680
rect 500944 362540 500978 362574
rect 502491 372953 502525 372987
rect 502491 372753 502525 372787
rect 502491 372553 502525 372587
rect 502491 372353 502525 372387
rect 502491 372153 502525 372187
rect 502491 371953 502525 371987
rect 502491 371753 502525 371787
rect 502491 371553 502525 371587
rect 502491 371353 502525 371387
rect 502491 371153 502525 371187
rect 502491 370953 502525 370987
rect 502491 370753 502525 370787
rect 502491 370553 502525 370587
rect 502491 370353 502525 370387
rect 502491 370153 502525 370187
rect 502491 369953 502525 369987
rect 502491 369753 502525 369787
rect 502491 369553 502525 369587
rect 502491 369353 502525 369387
rect 502491 369153 502525 369187
rect 502491 368953 502525 368987
rect 502491 368753 502525 368787
rect 502491 368553 502525 368587
rect 502491 368353 502525 368387
rect 502491 368153 502525 368187
rect 502491 367953 502525 367987
rect 502491 367753 502525 367787
rect 502491 367553 502525 367587
rect 502491 367353 502525 367387
rect 502491 367153 502525 367187
rect 502491 366953 502525 366987
rect 502491 366753 502525 366787
rect 502491 366553 502525 366587
rect 502491 366353 502525 366387
rect 502491 366153 502525 366187
rect 502491 365953 502525 365987
rect 502491 365753 502525 365787
rect 502491 365553 502525 365587
rect 502491 365353 502525 365387
rect 502491 365153 502525 365187
rect 502491 364953 502525 364987
rect 502491 364753 502525 364787
rect 502491 364553 502525 364587
rect 502491 364353 502525 364387
rect 502491 364153 502525 364187
rect 502491 363953 502525 363987
rect 502491 363753 502525 363787
rect 502491 363553 502525 363587
rect 502491 363353 502525 363387
rect 502491 363153 502525 363187
rect 502491 362953 502525 362987
rect 502491 362753 502525 362787
rect 502491 362553 502525 362587
rect 504371 372953 504405 372987
rect 504371 372753 504405 372787
rect 504371 372553 504405 372587
rect 504371 372353 504405 372387
rect 504371 372153 504405 372187
rect 504371 371953 504405 371987
rect 504371 371753 504405 371787
rect 504371 371553 504405 371587
rect 504371 371353 504405 371387
rect 504371 371153 504405 371187
rect 504371 370953 504405 370987
rect 504371 370753 504405 370787
rect 504371 370553 504405 370587
rect 504371 370353 504405 370387
rect 504371 370153 504405 370187
rect 504371 369953 504405 369987
rect 504371 369753 504405 369787
rect 504371 369553 504405 369587
rect 504371 369353 504405 369387
rect 504371 369153 504405 369187
rect 504371 368953 504405 368987
rect 504371 368753 504405 368787
rect 504371 368553 504405 368587
rect 504371 368353 504405 368387
rect 504371 368153 504405 368187
rect 504371 367953 504405 367987
rect 504371 367753 504405 367787
rect 504371 367553 504405 367587
rect 504371 367353 504405 367387
rect 504371 367153 504405 367187
rect 504371 366953 504405 366987
rect 504371 366753 504405 366787
rect 504371 366553 504405 366587
rect 504371 366353 504405 366387
rect 504371 366153 504405 366187
rect 504371 365953 504405 365987
rect 504371 365753 504405 365787
rect 504371 365553 504405 365587
rect 504371 365353 504405 365387
rect 504371 365153 504405 365187
rect 504371 364953 504405 364987
rect 504371 364753 504405 364787
rect 504371 364553 504405 364587
rect 504371 364353 504405 364387
rect 504371 364153 504405 364187
rect 504371 363953 504405 363987
rect 504371 363753 504405 363787
rect 504371 363553 504405 363587
rect 504371 363353 504405 363387
rect 504371 363153 504405 363187
rect 504371 362953 504405 362987
rect 504371 362753 504405 362787
rect 504371 362553 504405 362587
rect 504704 373090 504738 373124
rect 504704 373014 504738 373034
rect 504704 373000 504719 373014
rect 504719 373000 504738 373014
rect 504704 372924 504738 372944
rect 504704 372910 504719 372924
rect 504719 372910 504738 372924
rect 504704 372834 504738 372854
rect 504704 372820 504719 372834
rect 504719 372820 504738 372834
rect 504704 372744 504738 372764
rect 504704 372730 504719 372744
rect 504719 372730 504738 372744
rect 504704 372654 504738 372674
rect 504704 372640 504719 372654
rect 504719 372640 504738 372654
rect 504704 372564 504738 372584
rect 504704 372550 504719 372564
rect 504719 372550 504738 372564
rect 504704 372474 504738 372494
rect 504704 372460 504719 372474
rect 504719 372460 504738 372474
rect 504704 372384 504738 372404
rect 504704 372370 504719 372384
rect 504719 372370 504738 372384
rect 504704 372294 504738 372314
rect 504704 372280 504719 372294
rect 504719 372280 504738 372294
rect 504704 372204 504738 372224
rect 504704 372190 504719 372204
rect 504719 372190 504738 372204
rect 504704 372114 504738 372134
rect 504704 372100 504719 372114
rect 504719 372100 504738 372114
rect 504704 372024 504738 372044
rect 504704 372010 504719 372024
rect 504719 372010 504738 372024
rect 504864 372926 504898 372960
rect 504864 372850 504898 372870
rect 504864 372836 504866 372850
rect 504866 372836 504898 372850
rect 504864 372760 504898 372780
rect 504864 372746 504866 372760
rect 504866 372746 504898 372760
rect 504864 372670 504898 372690
rect 504864 372656 504866 372670
rect 504866 372656 504898 372670
rect 504864 372580 504898 372600
rect 504864 372566 504866 372580
rect 504866 372566 504898 372580
rect 504864 372490 504898 372510
rect 504864 372476 504866 372490
rect 504866 372476 504898 372490
rect 504864 372400 504898 372420
rect 504864 372386 504866 372400
rect 504866 372386 504898 372400
rect 504864 372310 504898 372330
rect 504864 372296 504866 372310
rect 504866 372296 504898 372310
rect 504864 372220 504898 372240
rect 504864 372206 504866 372220
rect 504866 372206 504898 372220
rect 505068 372752 505074 372774
rect 505074 372752 505102 372774
rect 505068 372740 505102 372752
rect 505168 372740 505202 372774
rect 505268 372740 505302 372774
rect 505368 372752 505400 372774
rect 505400 372752 505402 372774
rect 505468 372752 505490 372774
rect 505490 372752 505502 372774
rect 505568 372752 505580 372774
rect 505580 372752 505602 372774
rect 505368 372740 505402 372752
rect 505468 372740 505502 372752
rect 505568 372740 505602 372752
rect 505068 372662 505074 372674
rect 505074 372662 505102 372674
rect 505068 372640 505102 372662
rect 505168 372640 505202 372674
rect 505268 372640 505302 372674
rect 505368 372662 505400 372674
rect 505400 372662 505402 372674
rect 505468 372662 505490 372674
rect 505490 372662 505502 372674
rect 505568 372662 505580 372674
rect 505580 372662 505602 372674
rect 505368 372640 505402 372662
rect 505468 372640 505502 372662
rect 505568 372640 505602 372662
rect 505068 372572 505074 372574
rect 505074 372572 505102 372574
rect 505068 372540 505102 372572
rect 505168 372540 505202 372574
rect 505268 372540 505302 372574
rect 505368 372572 505400 372574
rect 505400 372572 505402 372574
rect 505468 372572 505490 372574
rect 505490 372572 505502 372574
rect 505568 372572 505580 372574
rect 505580 372572 505602 372574
rect 505368 372540 505402 372572
rect 505468 372540 505502 372572
rect 505568 372540 505602 372572
rect 505068 372440 505102 372474
rect 505168 372440 505202 372474
rect 505268 372440 505302 372474
rect 505368 372440 505402 372474
rect 505468 372440 505502 372474
rect 505568 372440 505602 372474
rect 505068 372340 505102 372374
rect 505168 372340 505202 372374
rect 505268 372340 505302 372374
rect 505368 372340 505402 372374
rect 505468 372340 505502 372374
rect 505568 372340 505602 372374
rect 505068 372246 505102 372274
rect 505068 372240 505074 372246
rect 505074 372240 505102 372246
rect 505168 372240 505202 372274
rect 505268 372240 505302 372274
rect 505368 372246 505402 372274
rect 505468 372246 505502 372274
rect 505568 372246 505602 372274
rect 505368 372240 505400 372246
rect 505400 372240 505402 372246
rect 505468 372240 505490 372246
rect 505490 372240 505502 372246
rect 505568 372240 505580 372246
rect 505580 372240 505602 372246
rect 504864 372130 504898 372150
rect 504864 372116 504866 372130
rect 504866 372116 504898 372130
rect 504864 372026 504898 372060
rect 504704 371920 504738 371954
rect 504704 371750 504738 371784
rect 504704 371674 504738 371694
rect 504704 371660 504719 371674
rect 504719 371660 504738 371674
rect 504704 371584 504738 371604
rect 504704 371570 504719 371584
rect 504719 371570 504738 371584
rect 504704 371494 504738 371514
rect 504704 371480 504719 371494
rect 504719 371480 504738 371494
rect 504704 371404 504738 371424
rect 504704 371390 504719 371404
rect 504719 371390 504738 371404
rect 504704 371314 504738 371334
rect 504704 371300 504719 371314
rect 504719 371300 504738 371314
rect 504704 371224 504738 371244
rect 504704 371210 504719 371224
rect 504719 371210 504738 371224
rect 504704 371134 504738 371154
rect 504704 371120 504719 371134
rect 504719 371120 504738 371134
rect 504704 371044 504738 371064
rect 504704 371030 504719 371044
rect 504719 371030 504738 371044
rect 504704 370954 504738 370974
rect 504704 370940 504719 370954
rect 504719 370940 504738 370954
rect 504704 370864 504738 370884
rect 504704 370850 504719 370864
rect 504719 370850 504738 370864
rect 504704 370774 504738 370794
rect 504704 370760 504719 370774
rect 504719 370760 504738 370774
rect 504704 370684 504738 370704
rect 504704 370670 504719 370684
rect 504719 370670 504738 370684
rect 504864 371586 504898 371620
rect 504864 371510 504898 371530
rect 504864 371496 504866 371510
rect 504866 371496 504898 371510
rect 504864 371420 504898 371440
rect 504864 371406 504866 371420
rect 504866 371406 504898 371420
rect 504864 371330 504898 371350
rect 504864 371316 504866 371330
rect 504866 371316 504898 371330
rect 504864 371240 504898 371260
rect 504864 371226 504866 371240
rect 504866 371226 504898 371240
rect 504864 371150 504898 371170
rect 504864 371136 504866 371150
rect 504866 371136 504898 371150
rect 504864 371060 504898 371080
rect 504864 371046 504866 371060
rect 504866 371046 504898 371060
rect 504864 370970 504898 370990
rect 504864 370956 504866 370970
rect 504866 370956 504898 370970
rect 504864 370880 504898 370900
rect 504864 370866 504866 370880
rect 504866 370866 504898 370880
rect 505068 371412 505074 371434
rect 505074 371412 505102 371434
rect 505068 371400 505102 371412
rect 505168 371400 505202 371434
rect 505268 371400 505302 371434
rect 505368 371412 505400 371434
rect 505400 371412 505402 371434
rect 505468 371412 505490 371434
rect 505490 371412 505502 371434
rect 505568 371412 505580 371434
rect 505580 371412 505602 371434
rect 505368 371400 505402 371412
rect 505468 371400 505502 371412
rect 505568 371400 505602 371412
rect 505068 371322 505074 371334
rect 505074 371322 505102 371334
rect 505068 371300 505102 371322
rect 505168 371300 505202 371334
rect 505268 371300 505302 371334
rect 505368 371322 505400 371334
rect 505400 371322 505402 371334
rect 505468 371322 505490 371334
rect 505490 371322 505502 371334
rect 505568 371322 505580 371334
rect 505580 371322 505602 371334
rect 505368 371300 505402 371322
rect 505468 371300 505502 371322
rect 505568 371300 505602 371322
rect 505068 371232 505074 371234
rect 505074 371232 505102 371234
rect 505068 371200 505102 371232
rect 505168 371200 505202 371234
rect 505268 371200 505302 371234
rect 505368 371232 505400 371234
rect 505400 371232 505402 371234
rect 505468 371232 505490 371234
rect 505490 371232 505502 371234
rect 505568 371232 505580 371234
rect 505580 371232 505602 371234
rect 505368 371200 505402 371232
rect 505468 371200 505502 371232
rect 505568 371200 505602 371232
rect 505068 371100 505102 371134
rect 505168 371100 505202 371134
rect 505268 371100 505302 371134
rect 505368 371100 505402 371134
rect 505468 371100 505502 371134
rect 505568 371100 505602 371134
rect 505068 371000 505102 371034
rect 505168 371000 505202 371034
rect 505268 371000 505302 371034
rect 505368 371000 505402 371034
rect 505468 371000 505502 371034
rect 505568 371000 505602 371034
rect 505068 370906 505102 370934
rect 505068 370900 505074 370906
rect 505074 370900 505102 370906
rect 505168 370900 505202 370934
rect 505268 370900 505302 370934
rect 505368 370906 505402 370934
rect 505468 370906 505502 370934
rect 505568 370906 505602 370934
rect 505368 370900 505400 370906
rect 505400 370900 505402 370906
rect 505468 370900 505490 370906
rect 505490 370900 505502 370906
rect 505568 370900 505580 370906
rect 505580 370900 505602 370906
rect 504864 370790 504898 370810
rect 504864 370776 504866 370790
rect 504866 370776 504898 370790
rect 504864 370686 504898 370720
rect 504704 370580 504738 370614
rect 504704 370410 504738 370444
rect 504704 370334 504738 370354
rect 504704 370320 504719 370334
rect 504719 370320 504738 370334
rect 504704 370244 504738 370264
rect 504704 370230 504719 370244
rect 504719 370230 504738 370244
rect 504704 370154 504738 370174
rect 504704 370140 504719 370154
rect 504719 370140 504738 370154
rect 504704 370064 504738 370084
rect 504704 370050 504719 370064
rect 504719 370050 504738 370064
rect 504704 369974 504738 369994
rect 504704 369960 504719 369974
rect 504719 369960 504738 369974
rect 504704 369884 504738 369904
rect 504704 369870 504719 369884
rect 504719 369870 504738 369884
rect 504704 369794 504738 369814
rect 504704 369780 504719 369794
rect 504719 369780 504738 369794
rect 504704 369704 504738 369724
rect 504704 369690 504719 369704
rect 504719 369690 504738 369704
rect 504704 369614 504738 369634
rect 504704 369600 504719 369614
rect 504719 369600 504738 369614
rect 504704 369524 504738 369544
rect 504704 369510 504719 369524
rect 504719 369510 504738 369524
rect 504704 369434 504738 369454
rect 504704 369420 504719 369434
rect 504719 369420 504738 369434
rect 504704 369344 504738 369364
rect 504704 369330 504719 369344
rect 504719 369330 504738 369344
rect 504864 370246 504898 370280
rect 504864 370170 504898 370190
rect 504864 370156 504866 370170
rect 504866 370156 504898 370170
rect 504864 370080 504898 370100
rect 504864 370066 504866 370080
rect 504866 370066 504898 370080
rect 504864 369990 504898 370010
rect 504864 369976 504866 369990
rect 504866 369976 504898 369990
rect 504864 369900 504898 369920
rect 504864 369886 504866 369900
rect 504866 369886 504898 369900
rect 504864 369810 504898 369830
rect 504864 369796 504866 369810
rect 504866 369796 504898 369810
rect 504864 369720 504898 369740
rect 504864 369706 504866 369720
rect 504866 369706 504898 369720
rect 504864 369630 504898 369650
rect 504864 369616 504866 369630
rect 504866 369616 504898 369630
rect 504864 369540 504898 369560
rect 504864 369526 504866 369540
rect 504866 369526 504898 369540
rect 505068 370072 505074 370094
rect 505074 370072 505102 370094
rect 505068 370060 505102 370072
rect 505168 370060 505202 370094
rect 505268 370060 505302 370094
rect 505368 370072 505400 370094
rect 505400 370072 505402 370094
rect 505468 370072 505490 370094
rect 505490 370072 505502 370094
rect 505568 370072 505580 370094
rect 505580 370072 505602 370094
rect 505368 370060 505402 370072
rect 505468 370060 505502 370072
rect 505568 370060 505602 370072
rect 505068 369982 505074 369994
rect 505074 369982 505102 369994
rect 505068 369960 505102 369982
rect 505168 369960 505202 369994
rect 505268 369960 505302 369994
rect 505368 369982 505400 369994
rect 505400 369982 505402 369994
rect 505468 369982 505490 369994
rect 505490 369982 505502 369994
rect 505568 369982 505580 369994
rect 505580 369982 505602 369994
rect 505368 369960 505402 369982
rect 505468 369960 505502 369982
rect 505568 369960 505602 369982
rect 505068 369892 505074 369894
rect 505074 369892 505102 369894
rect 505068 369860 505102 369892
rect 505168 369860 505202 369894
rect 505268 369860 505302 369894
rect 505368 369892 505400 369894
rect 505400 369892 505402 369894
rect 505468 369892 505490 369894
rect 505490 369892 505502 369894
rect 505568 369892 505580 369894
rect 505580 369892 505602 369894
rect 505368 369860 505402 369892
rect 505468 369860 505502 369892
rect 505568 369860 505602 369892
rect 505068 369760 505102 369794
rect 505168 369760 505202 369794
rect 505268 369760 505302 369794
rect 505368 369760 505402 369794
rect 505468 369760 505502 369794
rect 505568 369760 505602 369794
rect 505068 369660 505102 369694
rect 505168 369660 505202 369694
rect 505268 369660 505302 369694
rect 505368 369660 505402 369694
rect 505468 369660 505502 369694
rect 505568 369660 505602 369694
rect 505068 369566 505102 369594
rect 505068 369560 505074 369566
rect 505074 369560 505102 369566
rect 505168 369560 505202 369594
rect 505268 369560 505302 369594
rect 505368 369566 505402 369594
rect 505468 369566 505502 369594
rect 505568 369566 505602 369594
rect 505368 369560 505400 369566
rect 505400 369560 505402 369566
rect 505468 369560 505490 369566
rect 505490 369560 505502 369566
rect 505568 369560 505580 369566
rect 505580 369560 505602 369566
rect 504864 369450 504898 369470
rect 504864 369436 504866 369450
rect 504866 369436 504898 369450
rect 504864 369346 504898 369380
rect 504704 369240 504738 369274
rect 504704 369070 504738 369104
rect 504704 368994 504738 369014
rect 504704 368980 504719 368994
rect 504719 368980 504738 368994
rect 504704 368904 504738 368924
rect 504704 368890 504719 368904
rect 504719 368890 504738 368904
rect 504704 368814 504738 368834
rect 504704 368800 504719 368814
rect 504719 368800 504738 368814
rect 504704 368724 504738 368744
rect 504704 368710 504719 368724
rect 504719 368710 504738 368724
rect 504704 368634 504738 368654
rect 504704 368620 504719 368634
rect 504719 368620 504738 368634
rect 504704 368544 504738 368564
rect 504704 368530 504719 368544
rect 504719 368530 504738 368544
rect 504704 368454 504738 368474
rect 504704 368440 504719 368454
rect 504719 368440 504738 368454
rect 504704 368364 504738 368384
rect 504704 368350 504719 368364
rect 504719 368350 504738 368364
rect 504704 368274 504738 368294
rect 504704 368260 504719 368274
rect 504719 368260 504738 368274
rect 504704 368184 504738 368204
rect 504704 368170 504719 368184
rect 504719 368170 504738 368184
rect 504704 368094 504738 368114
rect 504704 368080 504719 368094
rect 504719 368080 504738 368094
rect 504704 368004 504738 368024
rect 504704 367990 504719 368004
rect 504719 367990 504738 368004
rect 504864 368906 504898 368940
rect 504864 368830 504898 368850
rect 504864 368816 504866 368830
rect 504866 368816 504898 368830
rect 504864 368740 504898 368760
rect 504864 368726 504866 368740
rect 504866 368726 504898 368740
rect 504864 368650 504898 368670
rect 504864 368636 504866 368650
rect 504866 368636 504898 368650
rect 504864 368560 504898 368580
rect 504864 368546 504866 368560
rect 504866 368546 504898 368560
rect 504864 368470 504898 368490
rect 504864 368456 504866 368470
rect 504866 368456 504898 368470
rect 504864 368380 504898 368400
rect 504864 368366 504866 368380
rect 504866 368366 504898 368380
rect 504864 368290 504898 368310
rect 504864 368276 504866 368290
rect 504866 368276 504898 368290
rect 504864 368200 504898 368220
rect 504864 368186 504866 368200
rect 504866 368186 504898 368200
rect 505068 368732 505074 368754
rect 505074 368732 505102 368754
rect 505068 368720 505102 368732
rect 505168 368720 505202 368754
rect 505268 368720 505302 368754
rect 505368 368732 505400 368754
rect 505400 368732 505402 368754
rect 505468 368732 505490 368754
rect 505490 368732 505502 368754
rect 505568 368732 505580 368754
rect 505580 368732 505602 368754
rect 505368 368720 505402 368732
rect 505468 368720 505502 368732
rect 505568 368720 505602 368732
rect 505068 368642 505074 368654
rect 505074 368642 505102 368654
rect 505068 368620 505102 368642
rect 505168 368620 505202 368654
rect 505268 368620 505302 368654
rect 505368 368642 505400 368654
rect 505400 368642 505402 368654
rect 505468 368642 505490 368654
rect 505490 368642 505502 368654
rect 505568 368642 505580 368654
rect 505580 368642 505602 368654
rect 505368 368620 505402 368642
rect 505468 368620 505502 368642
rect 505568 368620 505602 368642
rect 505068 368552 505074 368554
rect 505074 368552 505102 368554
rect 505068 368520 505102 368552
rect 505168 368520 505202 368554
rect 505268 368520 505302 368554
rect 505368 368552 505400 368554
rect 505400 368552 505402 368554
rect 505468 368552 505490 368554
rect 505490 368552 505502 368554
rect 505568 368552 505580 368554
rect 505580 368552 505602 368554
rect 505368 368520 505402 368552
rect 505468 368520 505502 368552
rect 505568 368520 505602 368552
rect 505068 368420 505102 368454
rect 505168 368420 505202 368454
rect 505268 368420 505302 368454
rect 505368 368420 505402 368454
rect 505468 368420 505502 368454
rect 505568 368420 505602 368454
rect 505068 368320 505102 368354
rect 505168 368320 505202 368354
rect 505268 368320 505302 368354
rect 505368 368320 505402 368354
rect 505468 368320 505502 368354
rect 505568 368320 505602 368354
rect 505068 368226 505102 368254
rect 505068 368220 505074 368226
rect 505074 368220 505102 368226
rect 505168 368220 505202 368254
rect 505268 368220 505302 368254
rect 505368 368226 505402 368254
rect 505468 368226 505502 368254
rect 505568 368226 505602 368254
rect 505368 368220 505400 368226
rect 505400 368220 505402 368226
rect 505468 368220 505490 368226
rect 505490 368220 505502 368226
rect 505568 368220 505580 368226
rect 505580 368220 505602 368226
rect 504864 368110 504898 368130
rect 504864 368096 504866 368110
rect 504866 368096 504898 368110
rect 504864 368006 504898 368040
rect 504704 367900 504738 367934
rect 504704 367730 504738 367764
rect 504704 367654 504738 367674
rect 504704 367640 504719 367654
rect 504719 367640 504738 367654
rect 504704 367564 504738 367584
rect 504704 367550 504719 367564
rect 504719 367550 504738 367564
rect 504704 367474 504738 367494
rect 504704 367460 504719 367474
rect 504719 367460 504738 367474
rect 504704 367384 504738 367404
rect 504704 367370 504719 367384
rect 504719 367370 504738 367384
rect 504704 367294 504738 367314
rect 504704 367280 504719 367294
rect 504719 367280 504738 367294
rect 504704 367204 504738 367224
rect 504704 367190 504719 367204
rect 504719 367190 504738 367204
rect 504704 367114 504738 367134
rect 504704 367100 504719 367114
rect 504719 367100 504738 367114
rect 504704 367024 504738 367044
rect 504704 367010 504719 367024
rect 504719 367010 504738 367024
rect 504704 366934 504738 366954
rect 504704 366920 504719 366934
rect 504719 366920 504738 366934
rect 504704 366844 504738 366864
rect 504704 366830 504719 366844
rect 504719 366830 504738 366844
rect 504704 366754 504738 366774
rect 504704 366740 504719 366754
rect 504719 366740 504738 366754
rect 504704 366664 504738 366684
rect 504704 366650 504719 366664
rect 504719 366650 504738 366664
rect 504864 367566 504898 367600
rect 504864 367490 504898 367510
rect 504864 367476 504866 367490
rect 504866 367476 504898 367490
rect 504864 367400 504898 367420
rect 504864 367386 504866 367400
rect 504866 367386 504898 367400
rect 504864 367310 504898 367330
rect 504864 367296 504866 367310
rect 504866 367296 504898 367310
rect 504864 367220 504898 367240
rect 504864 367206 504866 367220
rect 504866 367206 504898 367220
rect 504864 367130 504898 367150
rect 504864 367116 504866 367130
rect 504866 367116 504898 367130
rect 504864 367040 504898 367060
rect 504864 367026 504866 367040
rect 504866 367026 504898 367040
rect 504864 366950 504898 366970
rect 504864 366936 504866 366950
rect 504866 366936 504898 366950
rect 504864 366860 504898 366880
rect 504864 366846 504866 366860
rect 504866 366846 504898 366860
rect 505068 367392 505074 367414
rect 505074 367392 505102 367414
rect 505068 367380 505102 367392
rect 505168 367380 505202 367414
rect 505268 367380 505302 367414
rect 505368 367392 505400 367414
rect 505400 367392 505402 367414
rect 505468 367392 505490 367414
rect 505490 367392 505502 367414
rect 505568 367392 505580 367414
rect 505580 367392 505602 367414
rect 505368 367380 505402 367392
rect 505468 367380 505502 367392
rect 505568 367380 505602 367392
rect 505068 367302 505074 367314
rect 505074 367302 505102 367314
rect 505068 367280 505102 367302
rect 505168 367280 505202 367314
rect 505268 367280 505302 367314
rect 505368 367302 505400 367314
rect 505400 367302 505402 367314
rect 505468 367302 505490 367314
rect 505490 367302 505502 367314
rect 505568 367302 505580 367314
rect 505580 367302 505602 367314
rect 505368 367280 505402 367302
rect 505468 367280 505502 367302
rect 505568 367280 505602 367302
rect 505068 367212 505074 367214
rect 505074 367212 505102 367214
rect 505068 367180 505102 367212
rect 505168 367180 505202 367214
rect 505268 367180 505302 367214
rect 505368 367212 505400 367214
rect 505400 367212 505402 367214
rect 505468 367212 505490 367214
rect 505490 367212 505502 367214
rect 505568 367212 505580 367214
rect 505580 367212 505602 367214
rect 505368 367180 505402 367212
rect 505468 367180 505502 367212
rect 505568 367180 505602 367212
rect 505068 367080 505102 367114
rect 505168 367080 505202 367114
rect 505268 367080 505302 367114
rect 505368 367080 505402 367114
rect 505468 367080 505502 367114
rect 505568 367080 505602 367114
rect 505068 366980 505102 367014
rect 505168 366980 505202 367014
rect 505268 366980 505302 367014
rect 505368 366980 505402 367014
rect 505468 366980 505502 367014
rect 505568 366980 505602 367014
rect 505068 366886 505102 366914
rect 505068 366880 505074 366886
rect 505074 366880 505102 366886
rect 505168 366880 505202 366914
rect 505268 366880 505302 366914
rect 505368 366886 505402 366914
rect 505468 366886 505502 366914
rect 505568 366886 505602 366914
rect 505368 366880 505400 366886
rect 505400 366880 505402 366886
rect 505468 366880 505490 366886
rect 505490 366880 505502 366886
rect 505568 366880 505580 366886
rect 505580 366880 505602 366886
rect 504864 366770 504898 366790
rect 504864 366756 504866 366770
rect 504866 366756 504898 366770
rect 504864 366666 504898 366700
rect 504704 366560 504738 366594
rect 504704 366390 504738 366424
rect 504704 366314 504738 366334
rect 504704 366300 504719 366314
rect 504719 366300 504738 366314
rect 504704 366224 504738 366244
rect 504704 366210 504719 366224
rect 504719 366210 504738 366224
rect 504704 366134 504738 366154
rect 504704 366120 504719 366134
rect 504719 366120 504738 366134
rect 504704 366044 504738 366064
rect 504704 366030 504719 366044
rect 504719 366030 504738 366044
rect 504704 365954 504738 365974
rect 504704 365940 504719 365954
rect 504719 365940 504738 365954
rect 504704 365864 504738 365884
rect 504704 365850 504719 365864
rect 504719 365850 504738 365864
rect 504704 365774 504738 365794
rect 504704 365760 504719 365774
rect 504719 365760 504738 365774
rect 504704 365684 504738 365704
rect 504704 365670 504719 365684
rect 504719 365670 504738 365684
rect 504704 365594 504738 365614
rect 504704 365580 504719 365594
rect 504719 365580 504738 365594
rect 504704 365504 504738 365524
rect 504704 365490 504719 365504
rect 504719 365490 504738 365504
rect 504704 365414 504738 365434
rect 504704 365400 504719 365414
rect 504719 365400 504738 365414
rect 504704 365324 504738 365344
rect 504704 365310 504719 365324
rect 504719 365310 504738 365324
rect 504864 366226 504898 366260
rect 504864 366150 504898 366170
rect 504864 366136 504866 366150
rect 504866 366136 504898 366150
rect 504864 366060 504898 366080
rect 504864 366046 504866 366060
rect 504866 366046 504898 366060
rect 504864 365970 504898 365990
rect 504864 365956 504866 365970
rect 504866 365956 504898 365970
rect 504864 365880 504898 365900
rect 504864 365866 504866 365880
rect 504866 365866 504898 365880
rect 504864 365790 504898 365810
rect 504864 365776 504866 365790
rect 504866 365776 504898 365790
rect 504864 365700 504898 365720
rect 504864 365686 504866 365700
rect 504866 365686 504898 365700
rect 504864 365610 504898 365630
rect 504864 365596 504866 365610
rect 504866 365596 504898 365610
rect 504864 365520 504898 365540
rect 504864 365506 504866 365520
rect 504866 365506 504898 365520
rect 505068 366052 505074 366074
rect 505074 366052 505102 366074
rect 505068 366040 505102 366052
rect 505168 366040 505202 366074
rect 505268 366040 505302 366074
rect 505368 366052 505400 366074
rect 505400 366052 505402 366074
rect 505468 366052 505490 366074
rect 505490 366052 505502 366074
rect 505568 366052 505580 366074
rect 505580 366052 505602 366074
rect 505368 366040 505402 366052
rect 505468 366040 505502 366052
rect 505568 366040 505602 366052
rect 505068 365962 505074 365974
rect 505074 365962 505102 365974
rect 505068 365940 505102 365962
rect 505168 365940 505202 365974
rect 505268 365940 505302 365974
rect 505368 365962 505400 365974
rect 505400 365962 505402 365974
rect 505468 365962 505490 365974
rect 505490 365962 505502 365974
rect 505568 365962 505580 365974
rect 505580 365962 505602 365974
rect 505368 365940 505402 365962
rect 505468 365940 505502 365962
rect 505568 365940 505602 365962
rect 505068 365872 505074 365874
rect 505074 365872 505102 365874
rect 505068 365840 505102 365872
rect 505168 365840 505202 365874
rect 505268 365840 505302 365874
rect 505368 365872 505400 365874
rect 505400 365872 505402 365874
rect 505468 365872 505490 365874
rect 505490 365872 505502 365874
rect 505568 365872 505580 365874
rect 505580 365872 505602 365874
rect 505368 365840 505402 365872
rect 505468 365840 505502 365872
rect 505568 365840 505602 365872
rect 505068 365740 505102 365774
rect 505168 365740 505202 365774
rect 505268 365740 505302 365774
rect 505368 365740 505402 365774
rect 505468 365740 505502 365774
rect 505568 365740 505602 365774
rect 505068 365640 505102 365674
rect 505168 365640 505202 365674
rect 505268 365640 505302 365674
rect 505368 365640 505402 365674
rect 505468 365640 505502 365674
rect 505568 365640 505602 365674
rect 505068 365546 505102 365574
rect 505068 365540 505074 365546
rect 505074 365540 505102 365546
rect 505168 365540 505202 365574
rect 505268 365540 505302 365574
rect 505368 365546 505402 365574
rect 505468 365546 505502 365574
rect 505568 365546 505602 365574
rect 505368 365540 505400 365546
rect 505400 365540 505402 365546
rect 505468 365540 505490 365546
rect 505490 365540 505502 365546
rect 505568 365540 505580 365546
rect 505580 365540 505602 365546
rect 504864 365430 504898 365450
rect 504864 365416 504866 365430
rect 504866 365416 504898 365430
rect 504864 365326 504898 365360
rect 504704 365220 504738 365254
rect 504704 365050 504738 365084
rect 504704 364974 504738 364994
rect 504704 364960 504719 364974
rect 504719 364960 504738 364974
rect 504704 364884 504738 364904
rect 504704 364870 504719 364884
rect 504719 364870 504738 364884
rect 504704 364794 504738 364814
rect 504704 364780 504719 364794
rect 504719 364780 504738 364794
rect 504704 364704 504738 364724
rect 504704 364690 504719 364704
rect 504719 364690 504738 364704
rect 504704 364614 504738 364634
rect 504704 364600 504719 364614
rect 504719 364600 504738 364614
rect 504704 364524 504738 364544
rect 504704 364510 504719 364524
rect 504719 364510 504738 364524
rect 504704 364434 504738 364454
rect 504704 364420 504719 364434
rect 504719 364420 504738 364434
rect 504704 364344 504738 364364
rect 504704 364330 504719 364344
rect 504719 364330 504738 364344
rect 504704 364254 504738 364274
rect 504704 364240 504719 364254
rect 504719 364240 504738 364254
rect 504704 364164 504738 364184
rect 504704 364150 504719 364164
rect 504719 364150 504738 364164
rect 504704 364074 504738 364094
rect 504704 364060 504719 364074
rect 504719 364060 504738 364074
rect 504704 363984 504738 364004
rect 504704 363970 504719 363984
rect 504719 363970 504738 363984
rect 504864 364886 504898 364920
rect 504864 364810 504898 364830
rect 504864 364796 504866 364810
rect 504866 364796 504898 364810
rect 504864 364720 504898 364740
rect 504864 364706 504866 364720
rect 504866 364706 504898 364720
rect 504864 364630 504898 364650
rect 504864 364616 504866 364630
rect 504866 364616 504898 364630
rect 504864 364540 504898 364560
rect 504864 364526 504866 364540
rect 504866 364526 504898 364540
rect 504864 364450 504898 364470
rect 504864 364436 504866 364450
rect 504866 364436 504898 364450
rect 504864 364360 504898 364380
rect 504864 364346 504866 364360
rect 504866 364346 504898 364360
rect 504864 364270 504898 364290
rect 504864 364256 504866 364270
rect 504866 364256 504898 364270
rect 504864 364180 504898 364200
rect 504864 364166 504866 364180
rect 504866 364166 504898 364180
rect 505068 364712 505074 364734
rect 505074 364712 505102 364734
rect 505068 364700 505102 364712
rect 505168 364700 505202 364734
rect 505268 364700 505302 364734
rect 505368 364712 505400 364734
rect 505400 364712 505402 364734
rect 505468 364712 505490 364734
rect 505490 364712 505502 364734
rect 505568 364712 505580 364734
rect 505580 364712 505602 364734
rect 505368 364700 505402 364712
rect 505468 364700 505502 364712
rect 505568 364700 505602 364712
rect 505068 364622 505074 364634
rect 505074 364622 505102 364634
rect 505068 364600 505102 364622
rect 505168 364600 505202 364634
rect 505268 364600 505302 364634
rect 505368 364622 505400 364634
rect 505400 364622 505402 364634
rect 505468 364622 505490 364634
rect 505490 364622 505502 364634
rect 505568 364622 505580 364634
rect 505580 364622 505602 364634
rect 505368 364600 505402 364622
rect 505468 364600 505502 364622
rect 505568 364600 505602 364622
rect 505068 364532 505074 364534
rect 505074 364532 505102 364534
rect 505068 364500 505102 364532
rect 505168 364500 505202 364534
rect 505268 364500 505302 364534
rect 505368 364532 505400 364534
rect 505400 364532 505402 364534
rect 505468 364532 505490 364534
rect 505490 364532 505502 364534
rect 505568 364532 505580 364534
rect 505580 364532 505602 364534
rect 505368 364500 505402 364532
rect 505468 364500 505502 364532
rect 505568 364500 505602 364532
rect 505068 364400 505102 364434
rect 505168 364400 505202 364434
rect 505268 364400 505302 364434
rect 505368 364400 505402 364434
rect 505468 364400 505502 364434
rect 505568 364400 505602 364434
rect 505068 364300 505102 364334
rect 505168 364300 505202 364334
rect 505268 364300 505302 364334
rect 505368 364300 505402 364334
rect 505468 364300 505502 364334
rect 505568 364300 505602 364334
rect 505068 364206 505102 364234
rect 505068 364200 505074 364206
rect 505074 364200 505102 364206
rect 505168 364200 505202 364234
rect 505268 364200 505302 364234
rect 505368 364206 505402 364234
rect 505468 364206 505502 364234
rect 505568 364206 505602 364234
rect 505368 364200 505400 364206
rect 505400 364200 505402 364206
rect 505468 364200 505490 364206
rect 505490 364200 505502 364206
rect 505568 364200 505580 364206
rect 505580 364200 505602 364206
rect 504864 364090 504898 364110
rect 504864 364076 504866 364090
rect 504866 364076 504898 364090
rect 504864 363986 504898 364020
rect 504704 363880 504738 363914
rect 504704 363710 504738 363744
rect 504704 363634 504738 363654
rect 504704 363620 504719 363634
rect 504719 363620 504738 363634
rect 504704 363544 504738 363564
rect 504704 363530 504719 363544
rect 504719 363530 504738 363544
rect 504704 363454 504738 363474
rect 504704 363440 504719 363454
rect 504719 363440 504738 363454
rect 504704 363364 504738 363384
rect 504704 363350 504719 363364
rect 504719 363350 504738 363364
rect 504704 363274 504738 363294
rect 504704 363260 504719 363274
rect 504719 363260 504738 363274
rect 504704 363184 504738 363204
rect 504704 363170 504719 363184
rect 504719 363170 504738 363184
rect 504704 363094 504738 363114
rect 504704 363080 504719 363094
rect 504719 363080 504738 363094
rect 504704 363004 504738 363024
rect 504704 362990 504719 363004
rect 504719 362990 504738 363004
rect 504704 362914 504738 362934
rect 504704 362900 504719 362914
rect 504719 362900 504738 362914
rect 504704 362824 504738 362844
rect 504704 362810 504719 362824
rect 504719 362810 504738 362824
rect 504704 362734 504738 362754
rect 504704 362720 504719 362734
rect 504719 362720 504738 362734
rect 504704 362644 504738 362664
rect 504704 362630 504719 362644
rect 504719 362630 504738 362644
rect 504864 363546 504898 363580
rect 504864 363470 504898 363490
rect 504864 363456 504866 363470
rect 504866 363456 504898 363470
rect 504864 363380 504898 363400
rect 504864 363366 504866 363380
rect 504866 363366 504898 363380
rect 504864 363290 504898 363310
rect 504864 363276 504866 363290
rect 504866 363276 504898 363290
rect 504864 363200 504898 363220
rect 504864 363186 504866 363200
rect 504866 363186 504898 363200
rect 504864 363110 504898 363130
rect 504864 363096 504866 363110
rect 504866 363096 504898 363110
rect 504864 363020 504898 363040
rect 504864 363006 504866 363020
rect 504866 363006 504898 363020
rect 504864 362930 504898 362950
rect 504864 362916 504866 362930
rect 504866 362916 504898 362930
rect 504864 362840 504898 362860
rect 504864 362826 504866 362840
rect 504866 362826 504898 362840
rect 505068 363372 505074 363394
rect 505074 363372 505102 363394
rect 505068 363360 505102 363372
rect 505168 363360 505202 363394
rect 505268 363360 505302 363394
rect 505368 363372 505400 363394
rect 505400 363372 505402 363394
rect 505468 363372 505490 363394
rect 505490 363372 505502 363394
rect 505568 363372 505580 363394
rect 505580 363372 505602 363394
rect 505368 363360 505402 363372
rect 505468 363360 505502 363372
rect 505568 363360 505602 363372
rect 505068 363282 505074 363294
rect 505074 363282 505102 363294
rect 505068 363260 505102 363282
rect 505168 363260 505202 363294
rect 505268 363260 505302 363294
rect 505368 363282 505400 363294
rect 505400 363282 505402 363294
rect 505468 363282 505490 363294
rect 505490 363282 505502 363294
rect 505568 363282 505580 363294
rect 505580 363282 505602 363294
rect 505368 363260 505402 363282
rect 505468 363260 505502 363282
rect 505568 363260 505602 363282
rect 505068 363192 505074 363194
rect 505074 363192 505102 363194
rect 505068 363160 505102 363192
rect 505168 363160 505202 363194
rect 505268 363160 505302 363194
rect 505368 363192 505400 363194
rect 505400 363192 505402 363194
rect 505468 363192 505490 363194
rect 505490 363192 505502 363194
rect 505568 363192 505580 363194
rect 505580 363192 505602 363194
rect 505368 363160 505402 363192
rect 505468 363160 505502 363192
rect 505568 363160 505602 363192
rect 505068 363060 505102 363094
rect 505168 363060 505202 363094
rect 505268 363060 505302 363094
rect 505368 363060 505402 363094
rect 505468 363060 505502 363094
rect 505568 363060 505602 363094
rect 505068 362960 505102 362994
rect 505168 362960 505202 362994
rect 505268 362960 505302 362994
rect 505368 362960 505402 362994
rect 505468 362960 505502 362994
rect 505568 362960 505602 362994
rect 505068 362866 505102 362894
rect 505068 362860 505074 362866
rect 505074 362860 505102 362866
rect 505168 362860 505202 362894
rect 505268 362860 505302 362894
rect 505368 362866 505402 362894
rect 505468 362866 505502 362894
rect 505568 362866 505602 362894
rect 505368 362860 505400 362866
rect 505400 362860 505402 362866
rect 505468 362860 505490 362866
rect 505490 362860 505502 362866
rect 505568 362860 505580 362866
rect 505580 362860 505602 362866
rect 504864 362750 504898 362770
rect 504864 362736 504866 362750
rect 504866 362736 504898 362750
rect 504864 362646 504898 362680
rect 504704 362540 504738 362574
rect 506251 372953 506285 372987
rect 506251 372753 506285 372787
rect 506251 372553 506285 372587
rect 506251 372353 506285 372387
rect 506251 372153 506285 372187
rect 506251 371953 506285 371987
rect 506251 371753 506285 371787
rect 506251 371553 506285 371587
rect 506251 371353 506285 371387
rect 506251 371153 506285 371187
rect 506251 370953 506285 370987
rect 506251 370753 506285 370787
rect 506251 370553 506285 370587
rect 506251 370353 506285 370387
rect 506251 370153 506285 370187
rect 506251 369953 506285 369987
rect 506251 369753 506285 369787
rect 506251 369553 506285 369587
rect 506251 369353 506285 369387
rect 506251 369153 506285 369187
rect 506251 368953 506285 368987
rect 506251 368753 506285 368787
rect 506251 368553 506285 368587
rect 506251 368353 506285 368387
rect 506251 368153 506285 368187
rect 506251 367953 506285 367987
rect 506251 367753 506285 367787
rect 506251 367553 506285 367587
rect 506251 367353 506285 367387
rect 506251 367153 506285 367187
rect 506251 366953 506285 366987
rect 506251 366753 506285 366787
rect 506251 366553 506285 366587
rect 506251 366353 506285 366387
rect 506251 366153 506285 366187
rect 506251 365953 506285 365987
rect 506251 365753 506285 365787
rect 506251 365553 506285 365587
rect 506251 365353 506285 365387
rect 506251 365153 506285 365187
rect 506251 364953 506285 364987
rect 506251 364753 506285 364787
rect 506251 364553 506285 364587
rect 506251 364353 506285 364387
rect 506251 364153 506285 364187
rect 506251 363953 506285 363987
rect 506251 363753 506285 363787
rect 506251 363553 506285 363587
rect 506251 363353 506285 363387
rect 506251 363153 506285 363187
rect 506251 362953 506285 362987
rect 506251 362753 506285 362787
rect 506251 362553 506285 362587
rect 508131 372953 508165 372987
rect 508131 372753 508165 372787
rect 508131 372553 508165 372587
rect 508131 372353 508165 372387
rect 508131 372153 508165 372187
rect 508131 371953 508165 371987
rect 508131 371753 508165 371787
rect 508131 371553 508165 371587
rect 508131 371353 508165 371387
rect 508131 371153 508165 371187
rect 508131 370953 508165 370987
rect 508131 370753 508165 370787
rect 508131 370553 508165 370587
rect 508131 370353 508165 370387
rect 508131 370153 508165 370187
rect 508131 369953 508165 369987
rect 508131 369753 508165 369787
rect 508131 369553 508165 369587
rect 508131 369353 508165 369387
rect 508131 369153 508165 369187
rect 508131 368953 508165 368987
rect 508131 368753 508165 368787
rect 508131 368553 508165 368587
rect 508131 368353 508165 368387
rect 508131 368153 508165 368187
rect 508131 367953 508165 367987
rect 508131 367753 508165 367787
rect 508131 367553 508165 367587
rect 508131 367353 508165 367387
rect 508131 367153 508165 367187
rect 508131 366953 508165 366987
rect 508131 366753 508165 366787
rect 508131 366553 508165 366587
rect 508131 366353 508165 366387
rect 508131 366153 508165 366187
rect 508131 365953 508165 365987
rect 508131 365753 508165 365787
rect 508131 365553 508165 365587
rect 508131 365353 508165 365387
rect 508131 365153 508165 365187
rect 508131 364953 508165 364987
rect 508131 364753 508165 364787
rect 508131 364553 508165 364587
rect 508131 364353 508165 364387
rect 508131 364153 508165 364187
rect 508131 363953 508165 363987
rect 508131 363753 508165 363787
rect 508131 363553 508165 363587
rect 508131 363353 508165 363387
rect 508131 363153 508165 363187
rect 508131 362953 508165 362987
rect 508131 362753 508165 362787
rect 508131 362553 508165 362587
rect 508464 373090 508498 373124
rect 508464 373014 508498 373034
rect 508464 373000 508479 373014
rect 508479 373000 508498 373014
rect 508464 372924 508498 372944
rect 508464 372910 508479 372924
rect 508479 372910 508498 372924
rect 508464 372834 508498 372854
rect 508464 372820 508479 372834
rect 508479 372820 508498 372834
rect 508464 372744 508498 372764
rect 508464 372730 508479 372744
rect 508479 372730 508498 372744
rect 508464 372654 508498 372674
rect 508464 372640 508479 372654
rect 508479 372640 508498 372654
rect 508464 372564 508498 372584
rect 508464 372550 508479 372564
rect 508479 372550 508498 372564
rect 508464 372474 508498 372494
rect 508464 372460 508479 372474
rect 508479 372460 508498 372474
rect 508464 372384 508498 372404
rect 508464 372370 508479 372384
rect 508479 372370 508498 372384
rect 508464 372294 508498 372314
rect 508464 372280 508479 372294
rect 508479 372280 508498 372294
rect 508464 372204 508498 372224
rect 508464 372190 508479 372204
rect 508479 372190 508498 372204
rect 508464 372114 508498 372134
rect 508464 372100 508479 372114
rect 508479 372100 508498 372114
rect 508464 372024 508498 372044
rect 508464 372010 508479 372024
rect 508479 372010 508498 372024
rect 508624 372926 508658 372960
rect 508624 372850 508658 372870
rect 508624 372836 508626 372850
rect 508626 372836 508658 372850
rect 508624 372760 508658 372780
rect 508624 372746 508626 372760
rect 508626 372746 508658 372760
rect 508624 372670 508658 372690
rect 508624 372656 508626 372670
rect 508626 372656 508658 372670
rect 508624 372580 508658 372600
rect 508624 372566 508626 372580
rect 508626 372566 508658 372580
rect 508624 372490 508658 372510
rect 508624 372476 508626 372490
rect 508626 372476 508658 372490
rect 508624 372400 508658 372420
rect 508624 372386 508626 372400
rect 508626 372386 508658 372400
rect 508624 372310 508658 372330
rect 508624 372296 508626 372310
rect 508626 372296 508658 372310
rect 508624 372220 508658 372240
rect 508624 372206 508626 372220
rect 508626 372206 508658 372220
rect 508828 372752 508834 372774
rect 508834 372752 508862 372774
rect 508828 372740 508862 372752
rect 508928 372740 508962 372774
rect 509028 372740 509062 372774
rect 509128 372752 509160 372774
rect 509160 372752 509162 372774
rect 509228 372752 509250 372774
rect 509250 372752 509262 372774
rect 509328 372752 509340 372774
rect 509340 372752 509362 372774
rect 509128 372740 509162 372752
rect 509228 372740 509262 372752
rect 509328 372740 509362 372752
rect 508828 372662 508834 372674
rect 508834 372662 508862 372674
rect 508828 372640 508862 372662
rect 508928 372640 508962 372674
rect 509028 372640 509062 372674
rect 509128 372662 509160 372674
rect 509160 372662 509162 372674
rect 509228 372662 509250 372674
rect 509250 372662 509262 372674
rect 509328 372662 509340 372674
rect 509340 372662 509362 372674
rect 509128 372640 509162 372662
rect 509228 372640 509262 372662
rect 509328 372640 509362 372662
rect 508828 372572 508834 372574
rect 508834 372572 508862 372574
rect 508828 372540 508862 372572
rect 508928 372540 508962 372574
rect 509028 372540 509062 372574
rect 509128 372572 509160 372574
rect 509160 372572 509162 372574
rect 509228 372572 509250 372574
rect 509250 372572 509262 372574
rect 509328 372572 509340 372574
rect 509340 372572 509362 372574
rect 509128 372540 509162 372572
rect 509228 372540 509262 372572
rect 509328 372540 509362 372572
rect 508828 372440 508862 372474
rect 508928 372440 508962 372474
rect 509028 372440 509062 372474
rect 509128 372440 509162 372474
rect 509228 372440 509262 372474
rect 509328 372440 509362 372474
rect 508828 372340 508862 372374
rect 508928 372340 508962 372374
rect 509028 372340 509062 372374
rect 509128 372340 509162 372374
rect 509228 372340 509262 372374
rect 509328 372340 509362 372374
rect 508828 372246 508862 372274
rect 508828 372240 508834 372246
rect 508834 372240 508862 372246
rect 508928 372240 508962 372274
rect 509028 372240 509062 372274
rect 509128 372246 509162 372274
rect 509228 372246 509262 372274
rect 509328 372246 509362 372274
rect 509128 372240 509160 372246
rect 509160 372240 509162 372246
rect 509228 372240 509250 372246
rect 509250 372240 509262 372246
rect 509328 372240 509340 372246
rect 509340 372240 509362 372246
rect 508624 372130 508658 372150
rect 508624 372116 508626 372130
rect 508626 372116 508658 372130
rect 508624 372026 508658 372060
rect 508464 371920 508498 371954
rect 508464 371750 508498 371784
rect 508464 371674 508498 371694
rect 508464 371660 508479 371674
rect 508479 371660 508498 371674
rect 508464 371584 508498 371604
rect 508464 371570 508479 371584
rect 508479 371570 508498 371584
rect 508464 371494 508498 371514
rect 508464 371480 508479 371494
rect 508479 371480 508498 371494
rect 508464 371404 508498 371424
rect 508464 371390 508479 371404
rect 508479 371390 508498 371404
rect 508464 371314 508498 371334
rect 508464 371300 508479 371314
rect 508479 371300 508498 371314
rect 508464 371224 508498 371244
rect 508464 371210 508479 371224
rect 508479 371210 508498 371224
rect 508464 371134 508498 371154
rect 508464 371120 508479 371134
rect 508479 371120 508498 371134
rect 508464 371044 508498 371064
rect 508464 371030 508479 371044
rect 508479 371030 508498 371044
rect 508464 370954 508498 370974
rect 508464 370940 508479 370954
rect 508479 370940 508498 370954
rect 508464 370864 508498 370884
rect 508464 370850 508479 370864
rect 508479 370850 508498 370864
rect 508464 370774 508498 370794
rect 508464 370760 508479 370774
rect 508479 370760 508498 370774
rect 508464 370684 508498 370704
rect 508464 370670 508479 370684
rect 508479 370670 508498 370684
rect 508624 371586 508658 371620
rect 508624 371510 508658 371530
rect 508624 371496 508626 371510
rect 508626 371496 508658 371510
rect 508624 371420 508658 371440
rect 508624 371406 508626 371420
rect 508626 371406 508658 371420
rect 508624 371330 508658 371350
rect 508624 371316 508626 371330
rect 508626 371316 508658 371330
rect 508624 371240 508658 371260
rect 508624 371226 508626 371240
rect 508626 371226 508658 371240
rect 508624 371150 508658 371170
rect 508624 371136 508626 371150
rect 508626 371136 508658 371150
rect 508624 371060 508658 371080
rect 508624 371046 508626 371060
rect 508626 371046 508658 371060
rect 508624 370970 508658 370990
rect 508624 370956 508626 370970
rect 508626 370956 508658 370970
rect 508624 370880 508658 370900
rect 508624 370866 508626 370880
rect 508626 370866 508658 370880
rect 508828 371412 508834 371434
rect 508834 371412 508862 371434
rect 508828 371400 508862 371412
rect 508928 371400 508962 371434
rect 509028 371400 509062 371434
rect 509128 371412 509160 371434
rect 509160 371412 509162 371434
rect 509228 371412 509250 371434
rect 509250 371412 509262 371434
rect 509328 371412 509340 371434
rect 509340 371412 509362 371434
rect 509128 371400 509162 371412
rect 509228 371400 509262 371412
rect 509328 371400 509362 371412
rect 508828 371322 508834 371334
rect 508834 371322 508862 371334
rect 508828 371300 508862 371322
rect 508928 371300 508962 371334
rect 509028 371300 509062 371334
rect 509128 371322 509160 371334
rect 509160 371322 509162 371334
rect 509228 371322 509250 371334
rect 509250 371322 509262 371334
rect 509328 371322 509340 371334
rect 509340 371322 509362 371334
rect 509128 371300 509162 371322
rect 509228 371300 509262 371322
rect 509328 371300 509362 371322
rect 508828 371232 508834 371234
rect 508834 371232 508862 371234
rect 508828 371200 508862 371232
rect 508928 371200 508962 371234
rect 509028 371200 509062 371234
rect 509128 371232 509160 371234
rect 509160 371232 509162 371234
rect 509228 371232 509250 371234
rect 509250 371232 509262 371234
rect 509328 371232 509340 371234
rect 509340 371232 509362 371234
rect 509128 371200 509162 371232
rect 509228 371200 509262 371232
rect 509328 371200 509362 371232
rect 508828 371100 508862 371134
rect 508928 371100 508962 371134
rect 509028 371100 509062 371134
rect 509128 371100 509162 371134
rect 509228 371100 509262 371134
rect 509328 371100 509362 371134
rect 508828 371000 508862 371034
rect 508928 371000 508962 371034
rect 509028 371000 509062 371034
rect 509128 371000 509162 371034
rect 509228 371000 509262 371034
rect 509328 371000 509362 371034
rect 508828 370906 508862 370934
rect 508828 370900 508834 370906
rect 508834 370900 508862 370906
rect 508928 370900 508962 370934
rect 509028 370900 509062 370934
rect 509128 370906 509162 370934
rect 509228 370906 509262 370934
rect 509328 370906 509362 370934
rect 509128 370900 509160 370906
rect 509160 370900 509162 370906
rect 509228 370900 509250 370906
rect 509250 370900 509262 370906
rect 509328 370900 509340 370906
rect 509340 370900 509362 370906
rect 508624 370790 508658 370810
rect 508624 370776 508626 370790
rect 508626 370776 508658 370790
rect 508624 370686 508658 370720
rect 508464 370580 508498 370614
rect 508464 370410 508498 370444
rect 508464 370334 508498 370354
rect 508464 370320 508479 370334
rect 508479 370320 508498 370334
rect 508464 370244 508498 370264
rect 508464 370230 508479 370244
rect 508479 370230 508498 370244
rect 508464 370154 508498 370174
rect 508464 370140 508479 370154
rect 508479 370140 508498 370154
rect 508464 370064 508498 370084
rect 508464 370050 508479 370064
rect 508479 370050 508498 370064
rect 508464 369974 508498 369994
rect 508464 369960 508479 369974
rect 508479 369960 508498 369974
rect 508464 369884 508498 369904
rect 508464 369870 508479 369884
rect 508479 369870 508498 369884
rect 508464 369794 508498 369814
rect 508464 369780 508479 369794
rect 508479 369780 508498 369794
rect 508464 369704 508498 369724
rect 508464 369690 508479 369704
rect 508479 369690 508498 369704
rect 508464 369614 508498 369634
rect 508464 369600 508479 369614
rect 508479 369600 508498 369614
rect 508464 369524 508498 369544
rect 508464 369510 508479 369524
rect 508479 369510 508498 369524
rect 508464 369434 508498 369454
rect 508464 369420 508479 369434
rect 508479 369420 508498 369434
rect 508464 369344 508498 369364
rect 508464 369330 508479 369344
rect 508479 369330 508498 369344
rect 508624 370246 508658 370280
rect 508624 370170 508658 370190
rect 508624 370156 508626 370170
rect 508626 370156 508658 370170
rect 508624 370080 508658 370100
rect 508624 370066 508626 370080
rect 508626 370066 508658 370080
rect 508624 369990 508658 370010
rect 508624 369976 508626 369990
rect 508626 369976 508658 369990
rect 508624 369900 508658 369920
rect 508624 369886 508626 369900
rect 508626 369886 508658 369900
rect 508624 369810 508658 369830
rect 508624 369796 508626 369810
rect 508626 369796 508658 369810
rect 508624 369720 508658 369740
rect 508624 369706 508626 369720
rect 508626 369706 508658 369720
rect 508624 369630 508658 369650
rect 508624 369616 508626 369630
rect 508626 369616 508658 369630
rect 508624 369540 508658 369560
rect 508624 369526 508626 369540
rect 508626 369526 508658 369540
rect 508828 370072 508834 370094
rect 508834 370072 508862 370094
rect 508828 370060 508862 370072
rect 508928 370060 508962 370094
rect 509028 370060 509062 370094
rect 509128 370072 509160 370094
rect 509160 370072 509162 370094
rect 509228 370072 509250 370094
rect 509250 370072 509262 370094
rect 509328 370072 509340 370094
rect 509340 370072 509362 370094
rect 509128 370060 509162 370072
rect 509228 370060 509262 370072
rect 509328 370060 509362 370072
rect 508828 369982 508834 369994
rect 508834 369982 508862 369994
rect 508828 369960 508862 369982
rect 508928 369960 508962 369994
rect 509028 369960 509062 369994
rect 509128 369982 509160 369994
rect 509160 369982 509162 369994
rect 509228 369982 509250 369994
rect 509250 369982 509262 369994
rect 509328 369982 509340 369994
rect 509340 369982 509362 369994
rect 509128 369960 509162 369982
rect 509228 369960 509262 369982
rect 509328 369960 509362 369982
rect 508828 369892 508834 369894
rect 508834 369892 508862 369894
rect 508828 369860 508862 369892
rect 508928 369860 508962 369894
rect 509028 369860 509062 369894
rect 509128 369892 509160 369894
rect 509160 369892 509162 369894
rect 509228 369892 509250 369894
rect 509250 369892 509262 369894
rect 509328 369892 509340 369894
rect 509340 369892 509362 369894
rect 509128 369860 509162 369892
rect 509228 369860 509262 369892
rect 509328 369860 509362 369892
rect 508828 369760 508862 369794
rect 508928 369760 508962 369794
rect 509028 369760 509062 369794
rect 509128 369760 509162 369794
rect 509228 369760 509262 369794
rect 509328 369760 509362 369794
rect 508828 369660 508862 369694
rect 508928 369660 508962 369694
rect 509028 369660 509062 369694
rect 509128 369660 509162 369694
rect 509228 369660 509262 369694
rect 509328 369660 509362 369694
rect 508828 369566 508862 369594
rect 508828 369560 508834 369566
rect 508834 369560 508862 369566
rect 508928 369560 508962 369594
rect 509028 369560 509062 369594
rect 509128 369566 509162 369594
rect 509228 369566 509262 369594
rect 509328 369566 509362 369594
rect 509128 369560 509160 369566
rect 509160 369560 509162 369566
rect 509228 369560 509250 369566
rect 509250 369560 509262 369566
rect 509328 369560 509340 369566
rect 509340 369560 509362 369566
rect 508624 369450 508658 369470
rect 508624 369436 508626 369450
rect 508626 369436 508658 369450
rect 508624 369346 508658 369380
rect 508464 369240 508498 369274
rect 508464 369070 508498 369104
rect 508464 368994 508498 369014
rect 508464 368980 508479 368994
rect 508479 368980 508498 368994
rect 508464 368904 508498 368924
rect 508464 368890 508479 368904
rect 508479 368890 508498 368904
rect 508464 368814 508498 368834
rect 508464 368800 508479 368814
rect 508479 368800 508498 368814
rect 508464 368724 508498 368744
rect 508464 368710 508479 368724
rect 508479 368710 508498 368724
rect 508464 368634 508498 368654
rect 508464 368620 508479 368634
rect 508479 368620 508498 368634
rect 508464 368544 508498 368564
rect 508464 368530 508479 368544
rect 508479 368530 508498 368544
rect 508464 368454 508498 368474
rect 508464 368440 508479 368454
rect 508479 368440 508498 368454
rect 508464 368364 508498 368384
rect 508464 368350 508479 368364
rect 508479 368350 508498 368364
rect 508464 368274 508498 368294
rect 508464 368260 508479 368274
rect 508479 368260 508498 368274
rect 508464 368184 508498 368204
rect 508464 368170 508479 368184
rect 508479 368170 508498 368184
rect 508464 368094 508498 368114
rect 508464 368080 508479 368094
rect 508479 368080 508498 368094
rect 508464 368004 508498 368024
rect 508464 367990 508479 368004
rect 508479 367990 508498 368004
rect 508624 368906 508658 368940
rect 508624 368830 508658 368850
rect 508624 368816 508626 368830
rect 508626 368816 508658 368830
rect 508624 368740 508658 368760
rect 508624 368726 508626 368740
rect 508626 368726 508658 368740
rect 508624 368650 508658 368670
rect 508624 368636 508626 368650
rect 508626 368636 508658 368650
rect 508624 368560 508658 368580
rect 508624 368546 508626 368560
rect 508626 368546 508658 368560
rect 508624 368470 508658 368490
rect 508624 368456 508626 368470
rect 508626 368456 508658 368470
rect 508624 368380 508658 368400
rect 508624 368366 508626 368380
rect 508626 368366 508658 368380
rect 508624 368290 508658 368310
rect 508624 368276 508626 368290
rect 508626 368276 508658 368290
rect 508624 368200 508658 368220
rect 508624 368186 508626 368200
rect 508626 368186 508658 368200
rect 508828 368732 508834 368754
rect 508834 368732 508862 368754
rect 508828 368720 508862 368732
rect 508928 368720 508962 368754
rect 509028 368720 509062 368754
rect 509128 368732 509160 368754
rect 509160 368732 509162 368754
rect 509228 368732 509250 368754
rect 509250 368732 509262 368754
rect 509328 368732 509340 368754
rect 509340 368732 509362 368754
rect 509128 368720 509162 368732
rect 509228 368720 509262 368732
rect 509328 368720 509362 368732
rect 508828 368642 508834 368654
rect 508834 368642 508862 368654
rect 508828 368620 508862 368642
rect 508928 368620 508962 368654
rect 509028 368620 509062 368654
rect 509128 368642 509160 368654
rect 509160 368642 509162 368654
rect 509228 368642 509250 368654
rect 509250 368642 509262 368654
rect 509328 368642 509340 368654
rect 509340 368642 509362 368654
rect 509128 368620 509162 368642
rect 509228 368620 509262 368642
rect 509328 368620 509362 368642
rect 508828 368552 508834 368554
rect 508834 368552 508862 368554
rect 508828 368520 508862 368552
rect 508928 368520 508962 368554
rect 509028 368520 509062 368554
rect 509128 368552 509160 368554
rect 509160 368552 509162 368554
rect 509228 368552 509250 368554
rect 509250 368552 509262 368554
rect 509328 368552 509340 368554
rect 509340 368552 509362 368554
rect 509128 368520 509162 368552
rect 509228 368520 509262 368552
rect 509328 368520 509362 368552
rect 508828 368420 508862 368454
rect 508928 368420 508962 368454
rect 509028 368420 509062 368454
rect 509128 368420 509162 368454
rect 509228 368420 509262 368454
rect 509328 368420 509362 368454
rect 508828 368320 508862 368354
rect 508928 368320 508962 368354
rect 509028 368320 509062 368354
rect 509128 368320 509162 368354
rect 509228 368320 509262 368354
rect 509328 368320 509362 368354
rect 508828 368226 508862 368254
rect 508828 368220 508834 368226
rect 508834 368220 508862 368226
rect 508928 368220 508962 368254
rect 509028 368220 509062 368254
rect 509128 368226 509162 368254
rect 509228 368226 509262 368254
rect 509328 368226 509362 368254
rect 509128 368220 509160 368226
rect 509160 368220 509162 368226
rect 509228 368220 509250 368226
rect 509250 368220 509262 368226
rect 509328 368220 509340 368226
rect 509340 368220 509362 368226
rect 508624 368110 508658 368130
rect 508624 368096 508626 368110
rect 508626 368096 508658 368110
rect 508624 368006 508658 368040
rect 508464 367900 508498 367934
rect 508464 367730 508498 367764
rect 508464 367654 508498 367674
rect 508464 367640 508479 367654
rect 508479 367640 508498 367654
rect 508464 367564 508498 367584
rect 508464 367550 508479 367564
rect 508479 367550 508498 367564
rect 508464 367474 508498 367494
rect 508464 367460 508479 367474
rect 508479 367460 508498 367474
rect 508464 367384 508498 367404
rect 508464 367370 508479 367384
rect 508479 367370 508498 367384
rect 508464 367294 508498 367314
rect 508464 367280 508479 367294
rect 508479 367280 508498 367294
rect 508464 367204 508498 367224
rect 508464 367190 508479 367204
rect 508479 367190 508498 367204
rect 508464 367114 508498 367134
rect 508464 367100 508479 367114
rect 508479 367100 508498 367114
rect 508464 367024 508498 367044
rect 508464 367010 508479 367024
rect 508479 367010 508498 367024
rect 508464 366934 508498 366954
rect 508464 366920 508479 366934
rect 508479 366920 508498 366934
rect 508464 366844 508498 366864
rect 508464 366830 508479 366844
rect 508479 366830 508498 366844
rect 508464 366754 508498 366774
rect 508464 366740 508479 366754
rect 508479 366740 508498 366754
rect 508464 366664 508498 366684
rect 508464 366650 508479 366664
rect 508479 366650 508498 366664
rect 508624 367566 508658 367600
rect 508624 367490 508658 367510
rect 508624 367476 508626 367490
rect 508626 367476 508658 367490
rect 508624 367400 508658 367420
rect 508624 367386 508626 367400
rect 508626 367386 508658 367400
rect 508624 367310 508658 367330
rect 508624 367296 508626 367310
rect 508626 367296 508658 367310
rect 508624 367220 508658 367240
rect 508624 367206 508626 367220
rect 508626 367206 508658 367220
rect 508624 367130 508658 367150
rect 508624 367116 508626 367130
rect 508626 367116 508658 367130
rect 508624 367040 508658 367060
rect 508624 367026 508626 367040
rect 508626 367026 508658 367040
rect 508624 366950 508658 366970
rect 508624 366936 508626 366950
rect 508626 366936 508658 366950
rect 508624 366860 508658 366880
rect 508624 366846 508626 366860
rect 508626 366846 508658 366860
rect 508828 367392 508834 367414
rect 508834 367392 508862 367414
rect 508828 367380 508862 367392
rect 508928 367380 508962 367414
rect 509028 367380 509062 367414
rect 509128 367392 509160 367414
rect 509160 367392 509162 367414
rect 509228 367392 509250 367414
rect 509250 367392 509262 367414
rect 509328 367392 509340 367414
rect 509340 367392 509362 367414
rect 509128 367380 509162 367392
rect 509228 367380 509262 367392
rect 509328 367380 509362 367392
rect 508828 367302 508834 367314
rect 508834 367302 508862 367314
rect 508828 367280 508862 367302
rect 508928 367280 508962 367314
rect 509028 367280 509062 367314
rect 509128 367302 509160 367314
rect 509160 367302 509162 367314
rect 509228 367302 509250 367314
rect 509250 367302 509262 367314
rect 509328 367302 509340 367314
rect 509340 367302 509362 367314
rect 509128 367280 509162 367302
rect 509228 367280 509262 367302
rect 509328 367280 509362 367302
rect 508828 367212 508834 367214
rect 508834 367212 508862 367214
rect 508828 367180 508862 367212
rect 508928 367180 508962 367214
rect 509028 367180 509062 367214
rect 509128 367212 509160 367214
rect 509160 367212 509162 367214
rect 509228 367212 509250 367214
rect 509250 367212 509262 367214
rect 509328 367212 509340 367214
rect 509340 367212 509362 367214
rect 509128 367180 509162 367212
rect 509228 367180 509262 367212
rect 509328 367180 509362 367212
rect 508828 367080 508862 367114
rect 508928 367080 508962 367114
rect 509028 367080 509062 367114
rect 509128 367080 509162 367114
rect 509228 367080 509262 367114
rect 509328 367080 509362 367114
rect 508828 366980 508862 367014
rect 508928 366980 508962 367014
rect 509028 366980 509062 367014
rect 509128 366980 509162 367014
rect 509228 366980 509262 367014
rect 509328 366980 509362 367014
rect 508828 366886 508862 366914
rect 508828 366880 508834 366886
rect 508834 366880 508862 366886
rect 508928 366880 508962 366914
rect 509028 366880 509062 366914
rect 509128 366886 509162 366914
rect 509228 366886 509262 366914
rect 509328 366886 509362 366914
rect 509128 366880 509160 366886
rect 509160 366880 509162 366886
rect 509228 366880 509250 366886
rect 509250 366880 509262 366886
rect 509328 366880 509340 366886
rect 509340 366880 509362 366886
rect 508624 366770 508658 366790
rect 508624 366756 508626 366770
rect 508626 366756 508658 366770
rect 508624 366666 508658 366700
rect 508464 366560 508498 366594
rect 508464 366390 508498 366424
rect 508464 366314 508498 366334
rect 508464 366300 508479 366314
rect 508479 366300 508498 366314
rect 508464 366224 508498 366244
rect 508464 366210 508479 366224
rect 508479 366210 508498 366224
rect 508464 366134 508498 366154
rect 508464 366120 508479 366134
rect 508479 366120 508498 366134
rect 508464 366044 508498 366064
rect 508464 366030 508479 366044
rect 508479 366030 508498 366044
rect 508464 365954 508498 365974
rect 508464 365940 508479 365954
rect 508479 365940 508498 365954
rect 508464 365864 508498 365884
rect 508464 365850 508479 365864
rect 508479 365850 508498 365864
rect 508464 365774 508498 365794
rect 508464 365760 508479 365774
rect 508479 365760 508498 365774
rect 508464 365684 508498 365704
rect 508464 365670 508479 365684
rect 508479 365670 508498 365684
rect 508464 365594 508498 365614
rect 508464 365580 508479 365594
rect 508479 365580 508498 365594
rect 508464 365504 508498 365524
rect 508464 365490 508479 365504
rect 508479 365490 508498 365504
rect 508464 365414 508498 365434
rect 508464 365400 508479 365414
rect 508479 365400 508498 365414
rect 508464 365324 508498 365344
rect 508464 365310 508479 365324
rect 508479 365310 508498 365324
rect 508624 366226 508658 366260
rect 508624 366150 508658 366170
rect 508624 366136 508626 366150
rect 508626 366136 508658 366150
rect 508624 366060 508658 366080
rect 508624 366046 508626 366060
rect 508626 366046 508658 366060
rect 508624 365970 508658 365990
rect 508624 365956 508626 365970
rect 508626 365956 508658 365970
rect 508624 365880 508658 365900
rect 508624 365866 508626 365880
rect 508626 365866 508658 365880
rect 508624 365790 508658 365810
rect 508624 365776 508626 365790
rect 508626 365776 508658 365790
rect 508624 365700 508658 365720
rect 508624 365686 508626 365700
rect 508626 365686 508658 365700
rect 508624 365610 508658 365630
rect 508624 365596 508626 365610
rect 508626 365596 508658 365610
rect 508624 365520 508658 365540
rect 508624 365506 508626 365520
rect 508626 365506 508658 365520
rect 508828 366052 508834 366074
rect 508834 366052 508862 366074
rect 508828 366040 508862 366052
rect 508928 366040 508962 366074
rect 509028 366040 509062 366074
rect 509128 366052 509160 366074
rect 509160 366052 509162 366074
rect 509228 366052 509250 366074
rect 509250 366052 509262 366074
rect 509328 366052 509340 366074
rect 509340 366052 509362 366074
rect 509128 366040 509162 366052
rect 509228 366040 509262 366052
rect 509328 366040 509362 366052
rect 508828 365962 508834 365974
rect 508834 365962 508862 365974
rect 508828 365940 508862 365962
rect 508928 365940 508962 365974
rect 509028 365940 509062 365974
rect 509128 365962 509160 365974
rect 509160 365962 509162 365974
rect 509228 365962 509250 365974
rect 509250 365962 509262 365974
rect 509328 365962 509340 365974
rect 509340 365962 509362 365974
rect 509128 365940 509162 365962
rect 509228 365940 509262 365962
rect 509328 365940 509362 365962
rect 508828 365872 508834 365874
rect 508834 365872 508862 365874
rect 508828 365840 508862 365872
rect 508928 365840 508962 365874
rect 509028 365840 509062 365874
rect 509128 365872 509160 365874
rect 509160 365872 509162 365874
rect 509228 365872 509250 365874
rect 509250 365872 509262 365874
rect 509328 365872 509340 365874
rect 509340 365872 509362 365874
rect 509128 365840 509162 365872
rect 509228 365840 509262 365872
rect 509328 365840 509362 365872
rect 508828 365740 508862 365774
rect 508928 365740 508962 365774
rect 509028 365740 509062 365774
rect 509128 365740 509162 365774
rect 509228 365740 509262 365774
rect 509328 365740 509362 365774
rect 508828 365640 508862 365674
rect 508928 365640 508962 365674
rect 509028 365640 509062 365674
rect 509128 365640 509162 365674
rect 509228 365640 509262 365674
rect 509328 365640 509362 365674
rect 508828 365546 508862 365574
rect 508828 365540 508834 365546
rect 508834 365540 508862 365546
rect 508928 365540 508962 365574
rect 509028 365540 509062 365574
rect 509128 365546 509162 365574
rect 509228 365546 509262 365574
rect 509328 365546 509362 365574
rect 509128 365540 509160 365546
rect 509160 365540 509162 365546
rect 509228 365540 509250 365546
rect 509250 365540 509262 365546
rect 509328 365540 509340 365546
rect 509340 365540 509362 365546
rect 508624 365430 508658 365450
rect 508624 365416 508626 365430
rect 508626 365416 508658 365430
rect 508624 365326 508658 365360
rect 508464 365220 508498 365254
rect 508464 365050 508498 365084
rect 508464 364974 508498 364994
rect 508464 364960 508479 364974
rect 508479 364960 508498 364974
rect 508464 364884 508498 364904
rect 508464 364870 508479 364884
rect 508479 364870 508498 364884
rect 508464 364794 508498 364814
rect 508464 364780 508479 364794
rect 508479 364780 508498 364794
rect 508464 364704 508498 364724
rect 508464 364690 508479 364704
rect 508479 364690 508498 364704
rect 508464 364614 508498 364634
rect 508464 364600 508479 364614
rect 508479 364600 508498 364614
rect 508464 364524 508498 364544
rect 508464 364510 508479 364524
rect 508479 364510 508498 364524
rect 508464 364434 508498 364454
rect 508464 364420 508479 364434
rect 508479 364420 508498 364434
rect 508464 364344 508498 364364
rect 508464 364330 508479 364344
rect 508479 364330 508498 364344
rect 508464 364254 508498 364274
rect 508464 364240 508479 364254
rect 508479 364240 508498 364254
rect 508464 364164 508498 364184
rect 508464 364150 508479 364164
rect 508479 364150 508498 364164
rect 508464 364074 508498 364094
rect 508464 364060 508479 364074
rect 508479 364060 508498 364074
rect 508464 363984 508498 364004
rect 508464 363970 508479 363984
rect 508479 363970 508498 363984
rect 508624 364886 508658 364920
rect 508624 364810 508658 364830
rect 508624 364796 508626 364810
rect 508626 364796 508658 364810
rect 508624 364720 508658 364740
rect 508624 364706 508626 364720
rect 508626 364706 508658 364720
rect 508624 364630 508658 364650
rect 508624 364616 508626 364630
rect 508626 364616 508658 364630
rect 508624 364540 508658 364560
rect 508624 364526 508626 364540
rect 508626 364526 508658 364540
rect 508624 364450 508658 364470
rect 508624 364436 508626 364450
rect 508626 364436 508658 364450
rect 508624 364360 508658 364380
rect 508624 364346 508626 364360
rect 508626 364346 508658 364360
rect 508624 364270 508658 364290
rect 508624 364256 508626 364270
rect 508626 364256 508658 364270
rect 508624 364180 508658 364200
rect 508624 364166 508626 364180
rect 508626 364166 508658 364180
rect 508828 364712 508834 364734
rect 508834 364712 508862 364734
rect 508828 364700 508862 364712
rect 508928 364700 508962 364734
rect 509028 364700 509062 364734
rect 509128 364712 509160 364734
rect 509160 364712 509162 364734
rect 509228 364712 509250 364734
rect 509250 364712 509262 364734
rect 509328 364712 509340 364734
rect 509340 364712 509362 364734
rect 509128 364700 509162 364712
rect 509228 364700 509262 364712
rect 509328 364700 509362 364712
rect 508828 364622 508834 364634
rect 508834 364622 508862 364634
rect 508828 364600 508862 364622
rect 508928 364600 508962 364634
rect 509028 364600 509062 364634
rect 509128 364622 509160 364634
rect 509160 364622 509162 364634
rect 509228 364622 509250 364634
rect 509250 364622 509262 364634
rect 509328 364622 509340 364634
rect 509340 364622 509362 364634
rect 509128 364600 509162 364622
rect 509228 364600 509262 364622
rect 509328 364600 509362 364622
rect 508828 364532 508834 364534
rect 508834 364532 508862 364534
rect 508828 364500 508862 364532
rect 508928 364500 508962 364534
rect 509028 364500 509062 364534
rect 509128 364532 509160 364534
rect 509160 364532 509162 364534
rect 509228 364532 509250 364534
rect 509250 364532 509262 364534
rect 509328 364532 509340 364534
rect 509340 364532 509362 364534
rect 509128 364500 509162 364532
rect 509228 364500 509262 364532
rect 509328 364500 509362 364532
rect 508828 364400 508862 364434
rect 508928 364400 508962 364434
rect 509028 364400 509062 364434
rect 509128 364400 509162 364434
rect 509228 364400 509262 364434
rect 509328 364400 509362 364434
rect 508828 364300 508862 364334
rect 508928 364300 508962 364334
rect 509028 364300 509062 364334
rect 509128 364300 509162 364334
rect 509228 364300 509262 364334
rect 509328 364300 509362 364334
rect 508828 364206 508862 364234
rect 508828 364200 508834 364206
rect 508834 364200 508862 364206
rect 508928 364200 508962 364234
rect 509028 364200 509062 364234
rect 509128 364206 509162 364234
rect 509228 364206 509262 364234
rect 509328 364206 509362 364234
rect 509128 364200 509160 364206
rect 509160 364200 509162 364206
rect 509228 364200 509250 364206
rect 509250 364200 509262 364206
rect 509328 364200 509340 364206
rect 509340 364200 509362 364206
rect 508624 364090 508658 364110
rect 508624 364076 508626 364090
rect 508626 364076 508658 364090
rect 508624 363986 508658 364020
rect 508464 363880 508498 363914
rect 508464 363710 508498 363744
rect 508464 363634 508498 363654
rect 508464 363620 508479 363634
rect 508479 363620 508498 363634
rect 508464 363544 508498 363564
rect 508464 363530 508479 363544
rect 508479 363530 508498 363544
rect 508464 363454 508498 363474
rect 508464 363440 508479 363454
rect 508479 363440 508498 363454
rect 508464 363364 508498 363384
rect 508464 363350 508479 363364
rect 508479 363350 508498 363364
rect 508464 363274 508498 363294
rect 508464 363260 508479 363274
rect 508479 363260 508498 363274
rect 508464 363184 508498 363204
rect 508464 363170 508479 363184
rect 508479 363170 508498 363184
rect 508464 363094 508498 363114
rect 508464 363080 508479 363094
rect 508479 363080 508498 363094
rect 508464 363004 508498 363024
rect 508464 362990 508479 363004
rect 508479 362990 508498 363004
rect 508464 362914 508498 362934
rect 508464 362900 508479 362914
rect 508479 362900 508498 362914
rect 508464 362824 508498 362844
rect 508464 362810 508479 362824
rect 508479 362810 508498 362824
rect 508464 362734 508498 362754
rect 508464 362720 508479 362734
rect 508479 362720 508498 362734
rect 508464 362644 508498 362664
rect 508464 362630 508479 362644
rect 508479 362630 508498 362644
rect 508624 363546 508658 363580
rect 508624 363470 508658 363490
rect 508624 363456 508626 363470
rect 508626 363456 508658 363470
rect 508624 363380 508658 363400
rect 508624 363366 508626 363380
rect 508626 363366 508658 363380
rect 508624 363290 508658 363310
rect 508624 363276 508626 363290
rect 508626 363276 508658 363290
rect 508624 363200 508658 363220
rect 508624 363186 508626 363200
rect 508626 363186 508658 363200
rect 508624 363110 508658 363130
rect 508624 363096 508626 363110
rect 508626 363096 508658 363110
rect 508624 363020 508658 363040
rect 508624 363006 508626 363020
rect 508626 363006 508658 363020
rect 508624 362930 508658 362950
rect 508624 362916 508626 362930
rect 508626 362916 508658 362930
rect 508624 362840 508658 362860
rect 508624 362826 508626 362840
rect 508626 362826 508658 362840
rect 508828 363372 508834 363394
rect 508834 363372 508862 363394
rect 508828 363360 508862 363372
rect 508928 363360 508962 363394
rect 509028 363360 509062 363394
rect 509128 363372 509160 363394
rect 509160 363372 509162 363394
rect 509228 363372 509250 363394
rect 509250 363372 509262 363394
rect 509328 363372 509340 363394
rect 509340 363372 509362 363394
rect 509128 363360 509162 363372
rect 509228 363360 509262 363372
rect 509328 363360 509362 363372
rect 508828 363282 508834 363294
rect 508834 363282 508862 363294
rect 508828 363260 508862 363282
rect 508928 363260 508962 363294
rect 509028 363260 509062 363294
rect 509128 363282 509160 363294
rect 509160 363282 509162 363294
rect 509228 363282 509250 363294
rect 509250 363282 509262 363294
rect 509328 363282 509340 363294
rect 509340 363282 509362 363294
rect 509128 363260 509162 363282
rect 509228 363260 509262 363282
rect 509328 363260 509362 363282
rect 508828 363192 508834 363194
rect 508834 363192 508862 363194
rect 508828 363160 508862 363192
rect 508928 363160 508962 363194
rect 509028 363160 509062 363194
rect 509128 363192 509160 363194
rect 509160 363192 509162 363194
rect 509228 363192 509250 363194
rect 509250 363192 509262 363194
rect 509328 363192 509340 363194
rect 509340 363192 509362 363194
rect 509128 363160 509162 363192
rect 509228 363160 509262 363192
rect 509328 363160 509362 363192
rect 508828 363060 508862 363094
rect 508928 363060 508962 363094
rect 509028 363060 509062 363094
rect 509128 363060 509162 363094
rect 509228 363060 509262 363094
rect 509328 363060 509362 363094
rect 508828 362960 508862 362994
rect 508928 362960 508962 362994
rect 509028 362960 509062 362994
rect 509128 362960 509162 362994
rect 509228 362960 509262 362994
rect 509328 362960 509362 362994
rect 508828 362866 508862 362894
rect 508828 362860 508834 362866
rect 508834 362860 508862 362866
rect 508928 362860 508962 362894
rect 509028 362860 509062 362894
rect 509128 362866 509162 362894
rect 509228 362866 509262 362894
rect 509328 362866 509362 362894
rect 509128 362860 509160 362866
rect 509160 362860 509162 362866
rect 509228 362860 509250 362866
rect 509250 362860 509262 362866
rect 509328 362860 509340 362866
rect 509340 362860 509362 362866
rect 508624 362750 508658 362770
rect 508624 362736 508626 362750
rect 508626 362736 508658 362750
rect 508624 362646 508658 362680
rect 508464 362540 508498 362574
rect 510011 372953 510045 372987
rect 510011 372753 510045 372787
rect 510011 372553 510045 372587
rect 510011 372353 510045 372387
rect 510011 372153 510045 372187
rect 510011 371953 510045 371987
rect 510011 371753 510045 371787
rect 510011 371553 510045 371587
rect 510011 371353 510045 371387
rect 510011 371153 510045 371187
rect 510011 370953 510045 370987
rect 510011 370753 510045 370787
rect 510011 370553 510045 370587
rect 510011 370353 510045 370387
rect 510011 370153 510045 370187
rect 510011 369953 510045 369987
rect 510011 369753 510045 369787
rect 510011 369553 510045 369587
rect 510011 369353 510045 369387
rect 510011 369153 510045 369187
rect 510011 368953 510045 368987
rect 510011 368753 510045 368787
rect 510011 368553 510045 368587
rect 510011 368353 510045 368387
rect 510011 368153 510045 368187
rect 510011 367953 510045 367987
rect 510011 367753 510045 367787
rect 510011 367553 510045 367587
rect 510011 367353 510045 367387
rect 510011 367153 510045 367187
rect 510011 366953 510045 366987
rect 510011 366753 510045 366787
rect 510011 366553 510045 366587
rect 510011 366353 510045 366387
rect 510011 366153 510045 366187
rect 510011 365953 510045 365987
rect 510011 365753 510045 365787
rect 510011 365553 510045 365587
rect 510011 365353 510045 365387
rect 510011 365153 510045 365187
rect 510011 364953 510045 364987
rect 510011 364753 510045 364787
rect 510011 364553 510045 364587
rect 510011 364353 510045 364387
rect 510011 364153 510045 364187
rect 510011 363953 510045 363987
rect 510011 363753 510045 363787
rect 510011 363553 510045 363587
rect 510011 363353 510045 363387
rect 510011 363153 510045 363187
rect 510011 362953 510045 362987
rect 510011 362753 510045 362787
rect 510011 362553 510045 362587
rect 511891 372953 511925 372987
rect 511891 372753 511925 372787
rect 511891 372553 511925 372587
rect 511891 372353 511925 372387
rect 511891 372153 511925 372187
rect 511891 371953 511925 371987
rect 511891 371753 511925 371787
rect 511891 371553 511925 371587
rect 511891 371353 511925 371387
rect 511891 371153 511925 371187
rect 511891 370953 511925 370987
rect 511891 370753 511925 370787
rect 511891 370553 511925 370587
rect 511891 370353 511925 370387
rect 511891 370153 511925 370187
rect 511891 369953 511925 369987
rect 511891 369753 511925 369787
rect 511891 369553 511925 369587
rect 511891 369353 511925 369387
rect 511891 369153 511925 369187
rect 511891 368953 511925 368987
rect 511891 368753 511925 368787
rect 511891 368553 511925 368587
rect 511891 368353 511925 368387
rect 511891 368153 511925 368187
rect 511891 367953 511925 367987
rect 511891 367753 511925 367787
rect 511891 367553 511925 367587
rect 511891 367353 511925 367387
rect 511891 367153 511925 367187
rect 511891 366953 511925 366987
rect 511891 366753 511925 366787
rect 511891 366553 511925 366587
rect 511891 366353 511925 366387
rect 511891 366153 511925 366187
rect 511891 365953 511925 365987
rect 511891 365753 511925 365787
rect 511891 365553 511925 365587
rect 511891 365353 511925 365387
rect 511891 365153 511925 365187
rect 511891 364953 511925 364987
rect 511891 364753 511925 364787
rect 511891 364553 511925 364587
rect 511891 364353 511925 364387
rect 511891 364153 511925 364187
rect 511891 363953 511925 363987
rect 511891 363753 511925 363787
rect 511891 363553 511925 363587
rect 511891 363353 511925 363387
rect 511891 363153 511925 363187
rect 511891 362953 511925 362987
rect 511891 362753 511925 362787
rect 511891 362553 511925 362587
rect 512224 373090 512258 373124
rect 512224 373014 512258 373034
rect 512224 373000 512239 373014
rect 512239 373000 512258 373014
rect 512224 372924 512258 372944
rect 512224 372910 512239 372924
rect 512239 372910 512258 372924
rect 512224 372834 512258 372854
rect 512224 372820 512239 372834
rect 512239 372820 512258 372834
rect 512224 372744 512258 372764
rect 512224 372730 512239 372744
rect 512239 372730 512258 372744
rect 512224 372654 512258 372674
rect 512224 372640 512239 372654
rect 512239 372640 512258 372654
rect 512224 372564 512258 372584
rect 512224 372550 512239 372564
rect 512239 372550 512258 372564
rect 512224 372474 512258 372494
rect 512224 372460 512239 372474
rect 512239 372460 512258 372474
rect 512224 372384 512258 372404
rect 512224 372370 512239 372384
rect 512239 372370 512258 372384
rect 512224 372294 512258 372314
rect 512224 372280 512239 372294
rect 512239 372280 512258 372294
rect 512224 372204 512258 372224
rect 512224 372190 512239 372204
rect 512239 372190 512258 372204
rect 512224 372114 512258 372134
rect 512224 372100 512239 372114
rect 512239 372100 512258 372114
rect 512224 372024 512258 372044
rect 512224 372010 512239 372024
rect 512239 372010 512258 372024
rect 512384 372926 512418 372960
rect 512384 372850 512418 372870
rect 512384 372836 512386 372850
rect 512386 372836 512418 372850
rect 512384 372760 512418 372780
rect 512384 372746 512386 372760
rect 512386 372746 512418 372760
rect 512384 372670 512418 372690
rect 512384 372656 512386 372670
rect 512386 372656 512418 372670
rect 512384 372580 512418 372600
rect 512384 372566 512386 372580
rect 512386 372566 512418 372580
rect 512384 372490 512418 372510
rect 512384 372476 512386 372490
rect 512386 372476 512418 372490
rect 512384 372400 512418 372420
rect 512384 372386 512386 372400
rect 512386 372386 512418 372400
rect 512384 372310 512418 372330
rect 512384 372296 512386 372310
rect 512386 372296 512418 372310
rect 512384 372220 512418 372240
rect 512384 372206 512386 372220
rect 512386 372206 512418 372220
rect 512588 372752 512594 372774
rect 512594 372752 512622 372774
rect 512588 372740 512622 372752
rect 512688 372740 512722 372774
rect 512788 372740 512822 372774
rect 512888 372752 512920 372774
rect 512920 372752 512922 372774
rect 512988 372752 513010 372774
rect 513010 372752 513022 372774
rect 513088 372752 513100 372774
rect 513100 372752 513122 372774
rect 512888 372740 512922 372752
rect 512988 372740 513022 372752
rect 513088 372740 513122 372752
rect 512588 372662 512594 372674
rect 512594 372662 512622 372674
rect 512588 372640 512622 372662
rect 512688 372640 512722 372674
rect 512788 372640 512822 372674
rect 512888 372662 512920 372674
rect 512920 372662 512922 372674
rect 512988 372662 513010 372674
rect 513010 372662 513022 372674
rect 513088 372662 513100 372674
rect 513100 372662 513122 372674
rect 512888 372640 512922 372662
rect 512988 372640 513022 372662
rect 513088 372640 513122 372662
rect 512588 372572 512594 372574
rect 512594 372572 512622 372574
rect 512588 372540 512622 372572
rect 512688 372540 512722 372574
rect 512788 372540 512822 372574
rect 512888 372572 512920 372574
rect 512920 372572 512922 372574
rect 512988 372572 513010 372574
rect 513010 372572 513022 372574
rect 513088 372572 513100 372574
rect 513100 372572 513122 372574
rect 512888 372540 512922 372572
rect 512988 372540 513022 372572
rect 513088 372540 513122 372572
rect 512588 372440 512622 372474
rect 512688 372440 512722 372474
rect 512788 372440 512822 372474
rect 512888 372440 512922 372474
rect 512988 372440 513022 372474
rect 513088 372440 513122 372474
rect 512588 372340 512622 372374
rect 512688 372340 512722 372374
rect 512788 372340 512822 372374
rect 512888 372340 512922 372374
rect 512988 372340 513022 372374
rect 513088 372340 513122 372374
rect 512588 372246 512622 372274
rect 512588 372240 512594 372246
rect 512594 372240 512622 372246
rect 512688 372240 512722 372274
rect 512788 372240 512822 372274
rect 512888 372246 512922 372274
rect 512988 372246 513022 372274
rect 513088 372246 513122 372274
rect 512888 372240 512920 372246
rect 512920 372240 512922 372246
rect 512988 372240 513010 372246
rect 513010 372240 513022 372246
rect 513088 372240 513100 372246
rect 513100 372240 513122 372246
rect 512384 372130 512418 372150
rect 512384 372116 512386 372130
rect 512386 372116 512418 372130
rect 512384 372026 512418 372060
rect 512224 371920 512258 371954
rect 512224 371750 512258 371784
rect 512224 371674 512258 371694
rect 512224 371660 512239 371674
rect 512239 371660 512258 371674
rect 512224 371584 512258 371604
rect 512224 371570 512239 371584
rect 512239 371570 512258 371584
rect 512224 371494 512258 371514
rect 512224 371480 512239 371494
rect 512239 371480 512258 371494
rect 512224 371404 512258 371424
rect 512224 371390 512239 371404
rect 512239 371390 512258 371404
rect 512224 371314 512258 371334
rect 512224 371300 512239 371314
rect 512239 371300 512258 371314
rect 512224 371224 512258 371244
rect 512224 371210 512239 371224
rect 512239 371210 512258 371224
rect 512224 371134 512258 371154
rect 512224 371120 512239 371134
rect 512239 371120 512258 371134
rect 512224 371044 512258 371064
rect 512224 371030 512239 371044
rect 512239 371030 512258 371044
rect 512224 370954 512258 370974
rect 512224 370940 512239 370954
rect 512239 370940 512258 370954
rect 512224 370864 512258 370884
rect 512224 370850 512239 370864
rect 512239 370850 512258 370864
rect 512224 370774 512258 370794
rect 512224 370760 512239 370774
rect 512239 370760 512258 370774
rect 512224 370684 512258 370704
rect 512224 370670 512239 370684
rect 512239 370670 512258 370684
rect 512384 371586 512418 371620
rect 512384 371510 512418 371530
rect 512384 371496 512386 371510
rect 512386 371496 512418 371510
rect 512384 371420 512418 371440
rect 512384 371406 512386 371420
rect 512386 371406 512418 371420
rect 512384 371330 512418 371350
rect 512384 371316 512386 371330
rect 512386 371316 512418 371330
rect 512384 371240 512418 371260
rect 512384 371226 512386 371240
rect 512386 371226 512418 371240
rect 512384 371150 512418 371170
rect 512384 371136 512386 371150
rect 512386 371136 512418 371150
rect 512384 371060 512418 371080
rect 512384 371046 512386 371060
rect 512386 371046 512418 371060
rect 512384 370970 512418 370990
rect 512384 370956 512386 370970
rect 512386 370956 512418 370970
rect 512384 370880 512418 370900
rect 512384 370866 512386 370880
rect 512386 370866 512418 370880
rect 512588 371412 512594 371434
rect 512594 371412 512622 371434
rect 512588 371400 512622 371412
rect 512688 371400 512722 371434
rect 512788 371400 512822 371434
rect 512888 371412 512920 371434
rect 512920 371412 512922 371434
rect 512988 371412 513010 371434
rect 513010 371412 513022 371434
rect 513088 371412 513100 371434
rect 513100 371412 513122 371434
rect 512888 371400 512922 371412
rect 512988 371400 513022 371412
rect 513088 371400 513122 371412
rect 512588 371322 512594 371334
rect 512594 371322 512622 371334
rect 512588 371300 512622 371322
rect 512688 371300 512722 371334
rect 512788 371300 512822 371334
rect 512888 371322 512920 371334
rect 512920 371322 512922 371334
rect 512988 371322 513010 371334
rect 513010 371322 513022 371334
rect 513088 371322 513100 371334
rect 513100 371322 513122 371334
rect 512888 371300 512922 371322
rect 512988 371300 513022 371322
rect 513088 371300 513122 371322
rect 512588 371232 512594 371234
rect 512594 371232 512622 371234
rect 512588 371200 512622 371232
rect 512688 371200 512722 371234
rect 512788 371200 512822 371234
rect 512888 371232 512920 371234
rect 512920 371232 512922 371234
rect 512988 371232 513010 371234
rect 513010 371232 513022 371234
rect 513088 371232 513100 371234
rect 513100 371232 513122 371234
rect 512888 371200 512922 371232
rect 512988 371200 513022 371232
rect 513088 371200 513122 371232
rect 512588 371100 512622 371134
rect 512688 371100 512722 371134
rect 512788 371100 512822 371134
rect 512888 371100 512922 371134
rect 512988 371100 513022 371134
rect 513088 371100 513122 371134
rect 512588 371000 512622 371034
rect 512688 371000 512722 371034
rect 512788 371000 512822 371034
rect 512888 371000 512922 371034
rect 512988 371000 513022 371034
rect 513088 371000 513122 371034
rect 512588 370906 512622 370934
rect 512588 370900 512594 370906
rect 512594 370900 512622 370906
rect 512688 370900 512722 370934
rect 512788 370900 512822 370934
rect 512888 370906 512922 370934
rect 512988 370906 513022 370934
rect 513088 370906 513122 370934
rect 512888 370900 512920 370906
rect 512920 370900 512922 370906
rect 512988 370900 513010 370906
rect 513010 370900 513022 370906
rect 513088 370900 513100 370906
rect 513100 370900 513122 370906
rect 512384 370790 512418 370810
rect 512384 370776 512386 370790
rect 512386 370776 512418 370790
rect 512384 370686 512418 370720
rect 512224 370580 512258 370614
rect 512224 370410 512258 370444
rect 512224 370334 512258 370354
rect 512224 370320 512239 370334
rect 512239 370320 512258 370334
rect 512224 370244 512258 370264
rect 512224 370230 512239 370244
rect 512239 370230 512258 370244
rect 512224 370154 512258 370174
rect 512224 370140 512239 370154
rect 512239 370140 512258 370154
rect 512224 370064 512258 370084
rect 512224 370050 512239 370064
rect 512239 370050 512258 370064
rect 512224 369974 512258 369994
rect 512224 369960 512239 369974
rect 512239 369960 512258 369974
rect 512224 369884 512258 369904
rect 512224 369870 512239 369884
rect 512239 369870 512258 369884
rect 512224 369794 512258 369814
rect 512224 369780 512239 369794
rect 512239 369780 512258 369794
rect 512224 369704 512258 369724
rect 512224 369690 512239 369704
rect 512239 369690 512258 369704
rect 512224 369614 512258 369634
rect 512224 369600 512239 369614
rect 512239 369600 512258 369614
rect 512224 369524 512258 369544
rect 512224 369510 512239 369524
rect 512239 369510 512258 369524
rect 512224 369434 512258 369454
rect 512224 369420 512239 369434
rect 512239 369420 512258 369434
rect 512224 369344 512258 369364
rect 512224 369330 512239 369344
rect 512239 369330 512258 369344
rect 512384 370246 512418 370280
rect 512384 370170 512418 370190
rect 512384 370156 512386 370170
rect 512386 370156 512418 370170
rect 512384 370080 512418 370100
rect 512384 370066 512386 370080
rect 512386 370066 512418 370080
rect 512384 369990 512418 370010
rect 512384 369976 512386 369990
rect 512386 369976 512418 369990
rect 512384 369900 512418 369920
rect 512384 369886 512386 369900
rect 512386 369886 512418 369900
rect 512384 369810 512418 369830
rect 512384 369796 512386 369810
rect 512386 369796 512418 369810
rect 512384 369720 512418 369740
rect 512384 369706 512386 369720
rect 512386 369706 512418 369720
rect 512384 369630 512418 369650
rect 512384 369616 512386 369630
rect 512386 369616 512418 369630
rect 512384 369540 512418 369560
rect 512384 369526 512386 369540
rect 512386 369526 512418 369540
rect 512588 370072 512594 370094
rect 512594 370072 512622 370094
rect 512588 370060 512622 370072
rect 512688 370060 512722 370094
rect 512788 370060 512822 370094
rect 512888 370072 512920 370094
rect 512920 370072 512922 370094
rect 512988 370072 513010 370094
rect 513010 370072 513022 370094
rect 513088 370072 513100 370094
rect 513100 370072 513122 370094
rect 512888 370060 512922 370072
rect 512988 370060 513022 370072
rect 513088 370060 513122 370072
rect 512588 369982 512594 369994
rect 512594 369982 512622 369994
rect 512588 369960 512622 369982
rect 512688 369960 512722 369994
rect 512788 369960 512822 369994
rect 512888 369982 512920 369994
rect 512920 369982 512922 369994
rect 512988 369982 513010 369994
rect 513010 369982 513022 369994
rect 513088 369982 513100 369994
rect 513100 369982 513122 369994
rect 512888 369960 512922 369982
rect 512988 369960 513022 369982
rect 513088 369960 513122 369982
rect 512588 369892 512594 369894
rect 512594 369892 512622 369894
rect 512588 369860 512622 369892
rect 512688 369860 512722 369894
rect 512788 369860 512822 369894
rect 512888 369892 512920 369894
rect 512920 369892 512922 369894
rect 512988 369892 513010 369894
rect 513010 369892 513022 369894
rect 513088 369892 513100 369894
rect 513100 369892 513122 369894
rect 512888 369860 512922 369892
rect 512988 369860 513022 369892
rect 513088 369860 513122 369892
rect 512588 369760 512622 369794
rect 512688 369760 512722 369794
rect 512788 369760 512822 369794
rect 512888 369760 512922 369794
rect 512988 369760 513022 369794
rect 513088 369760 513122 369794
rect 512588 369660 512622 369694
rect 512688 369660 512722 369694
rect 512788 369660 512822 369694
rect 512888 369660 512922 369694
rect 512988 369660 513022 369694
rect 513088 369660 513122 369694
rect 512588 369566 512622 369594
rect 512588 369560 512594 369566
rect 512594 369560 512622 369566
rect 512688 369560 512722 369594
rect 512788 369560 512822 369594
rect 512888 369566 512922 369594
rect 512988 369566 513022 369594
rect 513088 369566 513122 369594
rect 512888 369560 512920 369566
rect 512920 369560 512922 369566
rect 512988 369560 513010 369566
rect 513010 369560 513022 369566
rect 513088 369560 513100 369566
rect 513100 369560 513122 369566
rect 512384 369450 512418 369470
rect 512384 369436 512386 369450
rect 512386 369436 512418 369450
rect 512384 369346 512418 369380
rect 512224 369240 512258 369274
rect 512224 369070 512258 369104
rect 512224 368994 512258 369014
rect 512224 368980 512239 368994
rect 512239 368980 512258 368994
rect 512224 368904 512258 368924
rect 512224 368890 512239 368904
rect 512239 368890 512258 368904
rect 512224 368814 512258 368834
rect 512224 368800 512239 368814
rect 512239 368800 512258 368814
rect 512224 368724 512258 368744
rect 512224 368710 512239 368724
rect 512239 368710 512258 368724
rect 512224 368634 512258 368654
rect 512224 368620 512239 368634
rect 512239 368620 512258 368634
rect 512224 368544 512258 368564
rect 512224 368530 512239 368544
rect 512239 368530 512258 368544
rect 512224 368454 512258 368474
rect 512224 368440 512239 368454
rect 512239 368440 512258 368454
rect 512224 368364 512258 368384
rect 512224 368350 512239 368364
rect 512239 368350 512258 368364
rect 512224 368274 512258 368294
rect 512224 368260 512239 368274
rect 512239 368260 512258 368274
rect 512224 368184 512258 368204
rect 512224 368170 512239 368184
rect 512239 368170 512258 368184
rect 512224 368094 512258 368114
rect 512224 368080 512239 368094
rect 512239 368080 512258 368094
rect 512224 368004 512258 368024
rect 512224 367990 512239 368004
rect 512239 367990 512258 368004
rect 512384 368906 512418 368940
rect 512384 368830 512418 368850
rect 512384 368816 512386 368830
rect 512386 368816 512418 368830
rect 512384 368740 512418 368760
rect 512384 368726 512386 368740
rect 512386 368726 512418 368740
rect 512384 368650 512418 368670
rect 512384 368636 512386 368650
rect 512386 368636 512418 368650
rect 512384 368560 512418 368580
rect 512384 368546 512386 368560
rect 512386 368546 512418 368560
rect 512384 368470 512418 368490
rect 512384 368456 512386 368470
rect 512386 368456 512418 368470
rect 512384 368380 512418 368400
rect 512384 368366 512386 368380
rect 512386 368366 512418 368380
rect 512384 368290 512418 368310
rect 512384 368276 512386 368290
rect 512386 368276 512418 368290
rect 512384 368200 512418 368220
rect 512384 368186 512386 368200
rect 512386 368186 512418 368200
rect 512588 368732 512594 368754
rect 512594 368732 512622 368754
rect 512588 368720 512622 368732
rect 512688 368720 512722 368754
rect 512788 368720 512822 368754
rect 512888 368732 512920 368754
rect 512920 368732 512922 368754
rect 512988 368732 513010 368754
rect 513010 368732 513022 368754
rect 513088 368732 513100 368754
rect 513100 368732 513122 368754
rect 512888 368720 512922 368732
rect 512988 368720 513022 368732
rect 513088 368720 513122 368732
rect 512588 368642 512594 368654
rect 512594 368642 512622 368654
rect 512588 368620 512622 368642
rect 512688 368620 512722 368654
rect 512788 368620 512822 368654
rect 512888 368642 512920 368654
rect 512920 368642 512922 368654
rect 512988 368642 513010 368654
rect 513010 368642 513022 368654
rect 513088 368642 513100 368654
rect 513100 368642 513122 368654
rect 512888 368620 512922 368642
rect 512988 368620 513022 368642
rect 513088 368620 513122 368642
rect 512588 368552 512594 368554
rect 512594 368552 512622 368554
rect 512588 368520 512622 368552
rect 512688 368520 512722 368554
rect 512788 368520 512822 368554
rect 512888 368552 512920 368554
rect 512920 368552 512922 368554
rect 512988 368552 513010 368554
rect 513010 368552 513022 368554
rect 513088 368552 513100 368554
rect 513100 368552 513122 368554
rect 512888 368520 512922 368552
rect 512988 368520 513022 368552
rect 513088 368520 513122 368552
rect 512588 368420 512622 368454
rect 512688 368420 512722 368454
rect 512788 368420 512822 368454
rect 512888 368420 512922 368454
rect 512988 368420 513022 368454
rect 513088 368420 513122 368454
rect 512588 368320 512622 368354
rect 512688 368320 512722 368354
rect 512788 368320 512822 368354
rect 512888 368320 512922 368354
rect 512988 368320 513022 368354
rect 513088 368320 513122 368354
rect 512588 368226 512622 368254
rect 512588 368220 512594 368226
rect 512594 368220 512622 368226
rect 512688 368220 512722 368254
rect 512788 368220 512822 368254
rect 512888 368226 512922 368254
rect 512988 368226 513022 368254
rect 513088 368226 513122 368254
rect 512888 368220 512920 368226
rect 512920 368220 512922 368226
rect 512988 368220 513010 368226
rect 513010 368220 513022 368226
rect 513088 368220 513100 368226
rect 513100 368220 513122 368226
rect 512384 368110 512418 368130
rect 512384 368096 512386 368110
rect 512386 368096 512418 368110
rect 512384 368006 512418 368040
rect 512224 367900 512258 367934
rect 512224 367730 512258 367764
rect 512224 367654 512258 367674
rect 512224 367640 512239 367654
rect 512239 367640 512258 367654
rect 512224 367564 512258 367584
rect 512224 367550 512239 367564
rect 512239 367550 512258 367564
rect 512224 367474 512258 367494
rect 512224 367460 512239 367474
rect 512239 367460 512258 367474
rect 512224 367384 512258 367404
rect 512224 367370 512239 367384
rect 512239 367370 512258 367384
rect 512224 367294 512258 367314
rect 512224 367280 512239 367294
rect 512239 367280 512258 367294
rect 512224 367204 512258 367224
rect 512224 367190 512239 367204
rect 512239 367190 512258 367204
rect 512224 367114 512258 367134
rect 512224 367100 512239 367114
rect 512239 367100 512258 367114
rect 512224 367024 512258 367044
rect 512224 367010 512239 367024
rect 512239 367010 512258 367024
rect 512224 366934 512258 366954
rect 512224 366920 512239 366934
rect 512239 366920 512258 366934
rect 512224 366844 512258 366864
rect 512224 366830 512239 366844
rect 512239 366830 512258 366844
rect 512224 366754 512258 366774
rect 512224 366740 512239 366754
rect 512239 366740 512258 366754
rect 512224 366664 512258 366684
rect 512224 366650 512239 366664
rect 512239 366650 512258 366664
rect 512384 367566 512418 367600
rect 512384 367490 512418 367510
rect 512384 367476 512386 367490
rect 512386 367476 512418 367490
rect 512384 367400 512418 367420
rect 512384 367386 512386 367400
rect 512386 367386 512418 367400
rect 512384 367310 512418 367330
rect 512384 367296 512386 367310
rect 512386 367296 512418 367310
rect 512384 367220 512418 367240
rect 512384 367206 512386 367220
rect 512386 367206 512418 367220
rect 512384 367130 512418 367150
rect 512384 367116 512386 367130
rect 512386 367116 512418 367130
rect 512384 367040 512418 367060
rect 512384 367026 512386 367040
rect 512386 367026 512418 367040
rect 512384 366950 512418 366970
rect 512384 366936 512386 366950
rect 512386 366936 512418 366950
rect 512384 366860 512418 366880
rect 512384 366846 512386 366860
rect 512386 366846 512418 366860
rect 512588 367392 512594 367414
rect 512594 367392 512622 367414
rect 512588 367380 512622 367392
rect 512688 367380 512722 367414
rect 512788 367380 512822 367414
rect 512888 367392 512920 367414
rect 512920 367392 512922 367414
rect 512988 367392 513010 367414
rect 513010 367392 513022 367414
rect 513088 367392 513100 367414
rect 513100 367392 513122 367414
rect 512888 367380 512922 367392
rect 512988 367380 513022 367392
rect 513088 367380 513122 367392
rect 512588 367302 512594 367314
rect 512594 367302 512622 367314
rect 512588 367280 512622 367302
rect 512688 367280 512722 367314
rect 512788 367280 512822 367314
rect 512888 367302 512920 367314
rect 512920 367302 512922 367314
rect 512988 367302 513010 367314
rect 513010 367302 513022 367314
rect 513088 367302 513100 367314
rect 513100 367302 513122 367314
rect 512888 367280 512922 367302
rect 512988 367280 513022 367302
rect 513088 367280 513122 367302
rect 512588 367212 512594 367214
rect 512594 367212 512622 367214
rect 512588 367180 512622 367212
rect 512688 367180 512722 367214
rect 512788 367180 512822 367214
rect 512888 367212 512920 367214
rect 512920 367212 512922 367214
rect 512988 367212 513010 367214
rect 513010 367212 513022 367214
rect 513088 367212 513100 367214
rect 513100 367212 513122 367214
rect 512888 367180 512922 367212
rect 512988 367180 513022 367212
rect 513088 367180 513122 367212
rect 512588 367080 512622 367114
rect 512688 367080 512722 367114
rect 512788 367080 512822 367114
rect 512888 367080 512922 367114
rect 512988 367080 513022 367114
rect 513088 367080 513122 367114
rect 512588 366980 512622 367014
rect 512688 366980 512722 367014
rect 512788 366980 512822 367014
rect 512888 366980 512922 367014
rect 512988 366980 513022 367014
rect 513088 366980 513122 367014
rect 512588 366886 512622 366914
rect 512588 366880 512594 366886
rect 512594 366880 512622 366886
rect 512688 366880 512722 366914
rect 512788 366880 512822 366914
rect 512888 366886 512922 366914
rect 512988 366886 513022 366914
rect 513088 366886 513122 366914
rect 512888 366880 512920 366886
rect 512920 366880 512922 366886
rect 512988 366880 513010 366886
rect 513010 366880 513022 366886
rect 513088 366880 513100 366886
rect 513100 366880 513122 366886
rect 512384 366770 512418 366790
rect 512384 366756 512386 366770
rect 512386 366756 512418 366770
rect 512384 366666 512418 366700
rect 512224 366560 512258 366594
rect 512224 366390 512258 366424
rect 512224 366314 512258 366334
rect 512224 366300 512239 366314
rect 512239 366300 512258 366314
rect 512224 366224 512258 366244
rect 512224 366210 512239 366224
rect 512239 366210 512258 366224
rect 512224 366134 512258 366154
rect 512224 366120 512239 366134
rect 512239 366120 512258 366134
rect 512224 366044 512258 366064
rect 512224 366030 512239 366044
rect 512239 366030 512258 366044
rect 512224 365954 512258 365974
rect 512224 365940 512239 365954
rect 512239 365940 512258 365954
rect 512224 365864 512258 365884
rect 512224 365850 512239 365864
rect 512239 365850 512258 365864
rect 512224 365774 512258 365794
rect 512224 365760 512239 365774
rect 512239 365760 512258 365774
rect 512224 365684 512258 365704
rect 512224 365670 512239 365684
rect 512239 365670 512258 365684
rect 512224 365594 512258 365614
rect 512224 365580 512239 365594
rect 512239 365580 512258 365594
rect 512224 365504 512258 365524
rect 512224 365490 512239 365504
rect 512239 365490 512258 365504
rect 512224 365414 512258 365434
rect 512224 365400 512239 365414
rect 512239 365400 512258 365414
rect 512224 365324 512258 365344
rect 512224 365310 512239 365324
rect 512239 365310 512258 365324
rect 512384 366226 512418 366260
rect 512384 366150 512418 366170
rect 512384 366136 512386 366150
rect 512386 366136 512418 366150
rect 512384 366060 512418 366080
rect 512384 366046 512386 366060
rect 512386 366046 512418 366060
rect 512384 365970 512418 365990
rect 512384 365956 512386 365970
rect 512386 365956 512418 365970
rect 512384 365880 512418 365900
rect 512384 365866 512386 365880
rect 512386 365866 512418 365880
rect 512384 365790 512418 365810
rect 512384 365776 512386 365790
rect 512386 365776 512418 365790
rect 512384 365700 512418 365720
rect 512384 365686 512386 365700
rect 512386 365686 512418 365700
rect 512384 365610 512418 365630
rect 512384 365596 512386 365610
rect 512386 365596 512418 365610
rect 512384 365520 512418 365540
rect 512384 365506 512386 365520
rect 512386 365506 512418 365520
rect 512588 366052 512594 366074
rect 512594 366052 512622 366074
rect 512588 366040 512622 366052
rect 512688 366040 512722 366074
rect 512788 366040 512822 366074
rect 512888 366052 512920 366074
rect 512920 366052 512922 366074
rect 512988 366052 513010 366074
rect 513010 366052 513022 366074
rect 513088 366052 513100 366074
rect 513100 366052 513122 366074
rect 512888 366040 512922 366052
rect 512988 366040 513022 366052
rect 513088 366040 513122 366052
rect 512588 365962 512594 365974
rect 512594 365962 512622 365974
rect 512588 365940 512622 365962
rect 512688 365940 512722 365974
rect 512788 365940 512822 365974
rect 512888 365962 512920 365974
rect 512920 365962 512922 365974
rect 512988 365962 513010 365974
rect 513010 365962 513022 365974
rect 513088 365962 513100 365974
rect 513100 365962 513122 365974
rect 512888 365940 512922 365962
rect 512988 365940 513022 365962
rect 513088 365940 513122 365962
rect 512588 365872 512594 365874
rect 512594 365872 512622 365874
rect 512588 365840 512622 365872
rect 512688 365840 512722 365874
rect 512788 365840 512822 365874
rect 512888 365872 512920 365874
rect 512920 365872 512922 365874
rect 512988 365872 513010 365874
rect 513010 365872 513022 365874
rect 513088 365872 513100 365874
rect 513100 365872 513122 365874
rect 512888 365840 512922 365872
rect 512988 365840 513022 365872
rect 513088 365840 513122 365872
rect 512588 365740 512622 365774
rect 512688 365740 512722 365774
rect 512788 365740 512822 365774
rect 512888 365740 512922 365774
rect 512988 365740 513022 365774
rect 513088 365740 513122 365774
rect 512588 365640 512622 365674
rect 512688 365640 512722 365674
rect 512788 365640 512822 365674
rect 512888 365640 512922 365674
rect 512988 365640 513022 365674
rect 513088 365640 513122 365674
rect 512588 365546 512622 365574
rect 512588 365540 512594 365546
rect 512594 365540 512622 365546
rect 512688 365540 512722 365574
rect 512788 365540 512822 365574
rect 512888 365546 512922 365574
rect 512988 365546 513022 365574
rect 513088 365546 513122 365574
rect 512888 365540 512920 365546
rect 512920 365540 512922 365546
rect 512988 365540 513010 365546
rect 513010 365540 513022 365546
rect 513088 365540 513100 365546
rect 513100 365540 513122 365546
rect 512384 365430 512418 365450
rect 512384 365416 512386 365430
rect 512386 365416 512418 365430
rect 512384 365326 512418 365360
rect 512224 365220 512258 365254
rect 512224 365050 512258 365084
rect 512224 364974 512258 364994
rect 512224 364960 512239 364974
rect 512239 364960 512258 364974
rect 512224 364884 512258 364904
rect 512224 364870 512239 364884
rect 512239 364870 512258 364884
rect 512224 364794 512258 364814
rect 512224 364780 512239 364794
rect 512239 364780 512258 364794
rect 512224 364704 512258 364724
rect 512224 364690 512239 364704
rect 512239 364690 512258 364704
rect 512224 364614 512258 364634
rect 512224 364600 512239 364614
rect 512239 364600 512258 364614
rect 512224 364524 512258 364544
rect 512224 364510 512239 364524
rect 512239 364510 512258 364524
rect 512224 364434 512258 364454
rect 512224 364420 512239 364434
rect 512239 364420 512258 364434
rect 512224 364344 512258 364364
rect 512224 364330 512239 364344
rect 512239 364330 512258 364344
rect 512224 364254 512258 364274
rect 512224 364240 512239 364254
rect 512239 364240 512258 364254
rect 512224 364164 512258 364184
rect 512224 364150 512239 364164
rect 512239 364150 512258 364164
rect 512224 364074 512258 364094
rect 512224 364060 512239 364074
rect 512239 364060 512258 364074
rect 512224 363984 512258 364004
rect 512224 363970 512239 363984
rect 512239 363970 512258 363984
rect 512384 364886 512418 364920
rect 512384 364810 512418 364830
rect 512384 364796 512386 364810
rect 512386 364796 512418 364810
rect 512384 364720 512418 364740
rect 512384 364706 512386 364720
rect 512386 364706 512418 364720
rect 512384 364630 512418 364650
rect 512384 364616 512386 364630
rect 512386 364616 512418 364630
rect 512384 364540 512418 364560
rect 512384 364526 512386 364540
rect 512386 364526 512418 364540
rect 512384 364450 512418 364470
rect 512384 364436 512386 364450
rect 512386 364436 512418 364450
rect 512384 364360 512418 364380
rect 512384 364346 512386 364360
rect 512386 364346 512418 364360
rect 512384 364270 512418 364290
rect 512384 364256 512386 364270
rect 512386 364256 512418 364270
rect 512384 364180 512418 364200
rect 512384 364166 512386 364180
rect 512386 364166 512418 364180
rect 512588 364712 512594 364734
rect 512594 364712 512622 364734
rect 512588 364700 512622 364712
rect 512688 364700 512722 364734
rect 512788 364700 512822 364734
rect 512888 364712 512920 364734
rect 512920 364712 512922 364734
rect 512988 364712 513010 364734
rect 513010 364712 513022 364734
rect 513088 364712 513100 364734
rect 513100 364712 513122 364734
rect 512888 364700 512922 364712
rect 512988 364700 513022 364712
rect 513088 364700 513122 364712
rect 512588 364622 512594 364634
rect 512594 364622 512622 364634
rect 512588 364600 512622 364622
rect 512688 364600 512722 364634
rect 512788 364600 512822 364634
rect 512888 364622 512920 364634
rect 512920 364622 512922 364634
rect 512988 364622 513010 364634
rect 513010 364622 513022 364634
rect 513088 364622 513100 364634
rect 513100 364622 513122 364634
rect 512888 364600 512922 364622
rect 512988 364600 513022 364622
rect 513088 364600 513122 364622
rect 512588 364532 512594 364534
rect 512594 364532 512622 364534
rect 512588 364500 512622 364532
rect 512688 364500 512722 364534
rect 512788 364500 512822 364534
rect 512888 364532 512920 364534
rect 512920 364532 512922 364534
rect 512988 364532 513010 364534
rect 513010 364532 513022 364534
rect 513088 364532 513100 364534
rect 513100 364532 513122 364534
rect 512888 364500 512922 364532
rect 512988 364500 513022 364532
rect 513088 364500 513122 364532
rect 512588 364400 512622 364434
rect 512688 364400 512722 364434
rect 512788 364400 512822 364434
rect 512888 364400 512922 364434
rect 512988 364400 513022 364434
rect 513088 364400 513122 364434
rect 512588 364300 512622 364334
rect 512688 364300 512722 364334
rect 512788 364300 512822 364334
rect 512888 364300 512922 364334
rect 512988 364300 513022 364334
rect 513088 364300 513122 364334
rect 512588 364206 512622 364234
rect 512588 364200 512594 364206
rect 512594 364200 512622 364206
rect 512688 364200 512722 364234
rect 512788 364200 512822 364234
rect 512888 364206 512922 364234
rect 512988 364206 513022 364234
rect 513088 364206 513122 364234
rect 512888 364200 512920 364206
rect 512920 364200 512922 364206
rect 512988 364200 513010 364206
rect 513010 364200 513022 364206
rect 513088 364200 513100 364206
rect 513100 364200 513122 364206
rect 512384 364090 512418 364110
rect 512384 364076 512386 364090
rect 512386 364076 512418 364090
rect 512384 363986 512418 364020
rect 512224 363880 512258 363914
rect 512224 363710 512258 363744
rect 512224 363634 512258 363654
rect 512224 363620 512239 363634
rect 512239 363620 512258 363634
rect 512224 363544 512258 363564
rect 512224 363530 512239 363544
rect 512239 363530 512258 363544
rect 512224 363454 512258 363474
rect 512224 363440 512239 363454
rect 512239 363440 512258 363454
rect 512224 363364 512258 363384
rect 512224 363350 512239 363364
rect 512239 363350 512258 363364
rect 512224 363274 512258 363294
rect 512224 363260 512239 363274
rect 512239 363260 512258 363274
rect 512224 363184 512258 363204
rect 512224 363170 512239 363184
rect 512239 363170 512258 363184
rect 512224 363094 512258 363114
rect 512224 363080 512239 363094
rect 512239 363080 512258 363094
rect 512224 363004 512258 363024
rect 512224 362990 512239 363004
rect 512239 362990 512258 363004
rect 512224 362914 512258 362934
rect 512224 362900 512239 362914
rect 512239 362900 512258 362914
rect 512224 362824 512258 362844
rect 512224 362810 512239 362824
rect 512239 362810 512258 362824
rect 512224 362734 512258 362754
rect 512224 362720 512239 362734
rect 512239 362720 512258 362734
rect 512224 362644 512258 362664
rect 512224 362630 512239 362644
rect 512239 362630 512258 362644
rect 512384 363546 512418 363580
rect 512384 363470 512418 363490
rect 512384 363456 512386 363470
rect 512386 363456 512418 363470
rect 512384 363380 512418 363400
rect 512384 363366 512386 363380
rect 512386 363366 512418 363380
rect 512384 363290 512418 363310
rect 512384 363276 512386 363290
rect 512386 363276 512418 363290
rect 512384 363200 512418 363220
rect 512384 363186 512386 363200
rect 512386 363186 512418 363200
rect 512384 363110 512418 363130
rect 512384 363096 512386 363110
rect 512386 363096 512418 363110
rect 512384 363020 512418 363040
rect 512384 363006 512386 363020
rect 512386 363006 512418 363020
rect 512384 362930 512418 362950
rect 512384 362916 512386 362930
rect 512386 362916 512418 362930
rect 512384 362840 512418 362860
rect 512384 362826 512386 362840
rect 512386 362826 512418 362840
rect 512588 363372 512594 363394
rect 512594 363372 512622 363394
rect 512588 363360 512622 363372
rect 512688 363360 512722 363394
rect 512788 363360 512822 363394
rect 512888 363372 512920 363394
rect 512920 363372 512922 363394
rect 512988 363372 513010 363394
rect 513010 363372 513022 363394
rect 513088 363372 513100 363394
rect 513100 363372 513122 363394
rect 512888 363360 512922 363372
rect 512988 363360 513022 363372
rect 513088 363360 513122 363372
rect 512588 363282 512594 363294
rect 512594 363282 512622 363294
rect 512588 363260 512622 363282
rect 512688 363260 512722 363294
rect 512788 363260 512822 363294
rect 512888 363282 512920 363294
rect 512920 363282 512922 363294
rect 512988 363282 513010 363294
rect 513010 363282 513022 363294
rect 513088 363282 513100 363294
rect 513100 363282 513122 363294
rect 512888 363260 512922 363282
rect 512988 363260 513022 363282
rect 513088 363260 513122 363282
rect 512588 363192 512594 363194
rect 512594 363192 512622 363194
rect 512588 363160 512622 363192
rect 512688 363160 512722 363194
rect 512788 363160 512822 363194
rect 512888 363192 512920 363194
rect 512920 363192 512922 363194
rect 512988 363192 513010 363194
rect 513010 363192 513022 363194
rect 513088 363192 513100 363194
rect 513100 363192 513122 363194
rect 512888 363160 512922 363192
rect 512988 363160 513022 363192
rect 513088 363160 513122 363192
rect 512588 363060 512622 363094
rect 512688 363060 512722 363094
rect 512788 363060 512822 363094
rect 512888 363060 512922 363094
rect 512988 363060 513022 363094
rect 513088 363060 513122 363094
rect 512588 362960 512622 362994
rect 512688 362960 512722 362994
rect 512788 362960 512822 362994
rect 512888 362960 512922 362994
rect 512988 362960 513022 362994
rect 513088 362960 513122 362994
rect 512588 362866 512622 362894
rect 512588 362860 512594 362866
rect 512594 362860 512622 362866
rect 512688 362860 512722 362894
rect 512788 362860 512822 362894
rect 512888 362866 512922 362894
rect 512988 362866 513022 362894
rect 513088 362866 513122 362894
rect 512888 362860 512920 362866
rect 512920 362860 512922 362866
rect 512988 362860 513010 362866
rect 513010 362860 513022 362866
rect 513088 362860 513100 362866
rect 513100 362860 513122 362866
rect 512384 362750 512418 362770
rect 512384 362736 512386 362750
rect 512386 362736 512418 362750
rect 512384 362646 512418 362680
rect 512224 362540 512258 362574
rect 513771 372953 513805 372987
rect 513771 372753 513805 372787
rect 513771 372553 513805 372587
rect 513771 372353 513805 372387
rect 515651 372999 515685 373033
rect 515651 372799 515685 372833
rect 517531 373199 517565 373233
rect 517531 372999 517565 373033
rect 515651 372599 515685 372633
rect 515919 372396 516457 372790
rect 516879 372396 517417 372790
rect 517531 372799 517565 372833
rect 517531 372599 517565 372633
rect 519411 374599 519445 374633
rect 519411 374399 519445 374433
rect 519679 374403 520217 374797
rect 520639 374403 521177 374797
rect 521291 374599 521325 374633
rect 521291 374399 521325 374433
rect 519411 374199 519445 374233
rect 519411 373999 519445 374033
rect 521291 374199 521325 374233
rect 521291 373999 521325 374033
rect 519411 373799 519445 373833
rect 519411 373599 519445 373633
rect 519411 373399 519445 373433
rect 521291 373799 521325 373833
rect 521291 373599 521325 373633
rect 521291 373399 521325 373433
rect 519411 373199 519445 373233
rect 519411 372999 519445 373033
rect 519411 372799 519445 372833
rect 521291 373199 521325 373233
rect 521291 372999 521325 373033
rect 519411 372599 519445 372633
rect 519679 372396 520217 372790
rect 520639 372396 521177 372790
rect 521291 372799 521325 372833
rect 521291 372599 521325 372633
rect 523171 374707 523205 374741
rect 523171 374307 523205 374341
rect 523171 373907 523205 373941
rect 523439 374471 523473 374505
rect 523511 374471 523541 374505
rect 523541 374471 523545 374505
rect 523583 374471 523609 374505
rect 523609 374471 523617 374505
rect 523655 374471 523677 374505
rect 523677 374471 523689 374505
rect 523727 374471 523745 374505
rect 523745 374471 523761 374505
rect 523799 374471 523813 374505
rect 523813 374471 523833 374505
rect 523871 374471 523881 374505
rect 523881 374471 523905 374505
rect 523943 374471 523949 374505
rect 523949 374471 523977 374505
rect 524015 374471 524017 374505
rect 524017 374471 524049 374505
rect 524087 374471 524119 374505
rect 524119 374471 524121 374505
rect 524159 374471 524187 374505
rect 524187 374471 524193 374505
rect 524231 374471 524255 374505
rect 524255 374471 524265 374505
rect 524303 374471 524323 374505
rect 524323 374471 524337 374505
rect 524375 374471 524391 374505
rect 524391 374471 524409 374505
rect 524447 374471 524459 374505
rect 524459 374471 524481 374505
rect 524519 374471 524527 374505
rect 524527 374471 524553 374505
rect 524591 374471 524595 374505
rect 524595 374471 524625 374505
rect 524663 374471 524697 374505
rect 523439 374013 523473 374047
rect 523511 374013 523541 374047
rect 523541 374013 523545 374047
rect 523583 374013 523609 374047
rect 523609 374013 523617 374047
rect 523655 374013 523677 374047
rect 523677 374013 523689 374047
rect 523727 374013 523745 374047
rect 523745 374013 523761 374047
rect 523799 374013 523813 374047
rect 523813 374013 523833 374047
rect 523871 374013 523881 374047
rect 523881 374013 523905 374047
rect 523943 374013 523949 374047
rect 523949 374013 523977 374047
rect 524015 374013 524017 374047
rect 524017 374013 524049 374047
rect 524087 374013 524119 374047
rect 524119 374013 524121 374047
rect 524159 374013 524187 374047
rect 524187 374013 524193 374047
rect 524231 374013 524255 374047
rect 524255 374013 524265 374047
rect 524303 374013 524323 374047
rect 524323 374013 524337 374047
rect 524375 374013 524391 374047
rect 524391 374013 524409 374047
rect 524447 374013 524459 374047
rect 524459 374013 524481 374047
rect 524519 374013 524527 374047
rect 524527 374013 524553 374047
rect 524591 374013 524595 374047
rect 524595 374013 524625 374047
rect 524663 374013 524697 374047
rect 523171 373507 523205 373541
rect 523171 373107 523205 373141
rect 523171 372707 523205 372741
rect 513771 372153 513805 372187
rect 523171 372307 523205 372341
rect 523439 373555 523473 373589
rect 523511 373555 523541 373589
rect 523541 373555 523545 373589
rect 523583 373555 523609 373589
rect 523609 373555 523617 373589
rect 523655 373555 523677 373589
rect 523677 373555 523689 373589
rect 523727 373555 523745 373589
rect 523745 373555 523761 373589
rect 523799 373555 523813 373589
rect 523813 373555 523833 373589
rect 523871 373555 523881 373589
rect 523881 373555 523905 373589
rect 523943 373555 523949 373589
rect 523949 373555 523977 373589
rect 524015 373555 524017 373589
rect 524017 373555 524049 373589
rect 524087 373555 524119 373589
rect 524119 373555 524121 373589
rect 524159 373555 524187 373589
rect 524187 373555 524193 373589
rect 524231 373555 524255 373589
rect 524255 373555 524265 373589
rect 524303 373555 524323 373589
rect 524323 373555 524337 373589
rect 524375 373555 524391 373589
rect 524391 373555 524409 373589
rect 524447 373555 524459 373589
rect 524459 373555 524481 373589
rect 524519 373555 524527 373589
rect 524527 373555 524553 373589
rect 524591 373555 524595 373589
rect 524595 373555 524625 373589
rect 524663 373555 524697 373589
rect 523439 373097 523473 373131
rect 523511 373097 523541 373131
rect 523541 373097 523545 373131
rect 523583 373097 523609 373131
rect 523609 373097 523617 373131
rect 523655 373097 523677 373131
rect 523677 373097 523689 373131
rect 523727 373097 523745 373131
rect 523745 373097 523761 373131
rect 523799 373097 523813 373131
rect 523813 373097 523833 373131
rect 523871 373097 523881 373131
rect 523881 373097 523905 373131
rect 523943 373097 523949 373131
rect 523949 373097 523977 373131
rect 524015 373097 524017 373131
rect 524017 373097 524049 373131
rect 524087 373097 524119 373131
rect 524119 373097 524121 373131
rect 524159 373097 524187 373131
rect 524187 373097 524193 373131
rect 524231 373097 524255 373131
rect 524255 373097 524265 373131
rect 524303 373097 524323 373131
rect 524323 373097 524337 373131
rect 524375 373097 524391 373131
rect 524391 373097 524409 373131
rect 524447 373097 524459 373131
rect 524459 373097 524481 373131
rect 524519 373097 524527 373131
rect 524527 373097 524553 373131
rect 524591 373097 524595 373131
rect 524595 373097 524625 373131
rect 524663 373097 524697 373131
rect 523439 372639 523473 372673
rect 523511 372639 523541 372673
rect 523541 372639 523545 372673
rect 523583 372639 523609 372673
rect 523609 372639 523617 372673
rect 523655 372639 523677 372673
rect 523677 372639 523689 372673
rect 523727 372639 523745 372673
rect 523745 372639 523761 372673
rect 523799 372639 523813 372673
rect 523813 372639 523833 372673
rect 523871 372639 523881 372673
rect 523881 372639 523905 372673
rect 523943 372639 523949 372673
rect 523949 372639 523977 372673
rect 524015 372639 524017 372673
rect 524017 372639 524049 372673
rect 524087 372639 524119 372673
rect 524119 372639 524121 372673
rect 524159 372639 524187 372673
rect 524187 372639 524193 372673
rect 524231 372639 524255 372673
rect 524255 372639 524265 372673
rect 524303 372639 524323 372673
rect 524323 372639 524337 372673
rect 524375 372639 524391 372673
rect 524391 372639 524409 372673
rect 524447 372639 524459 372673
rect 524459 372639 524481 372673
rect 524519 372639 524527 372673
rect 524527 372639 524553 372673
rect 524591 372639 524595 372673
rect 524595 372639 524625 372673
rect 524663 372639 524697 372673
rect 523439 372181 523473 372215
rect 523511 372181 523541 372215
rect 523541 372181 523545 372215
rect 523583 372181 523609 372215
rect 523609 372181 523617 372215
rect 523655 372181 523677 372215
rect 523677 372181 523689 372215
rect 523727 372181 523745 372215
rect 523745 372181 523761 372215
rect 523799 372181 523813 372215
rect 523813 372181 523833 372215
rect 523871 372181 523881 372215
rect 523881 372181 523905 372215
rect 523943 372181 523949 372215
rect 523949 372181 523977 372215
rect 524015 372181 524017 372215
rect 524017 372181 524049 372215
rect 524087 372181 524119 372215
rect 524119 372181 524121 372215
rect 524159 372181 524187 372215
rect 524187 372181 524193 372215
rect 524231 372181 524255 372215
rect 524255 372181 524265 372215
rect 524303 372181 524323 372215
rect 524323 372181 524337 372215
rect 524375 372181 524391 372215
rect 524391 372181 524409 372215
rect 524447 372181 524459 372215
rect 524459 372181 524481 372215
rect 524519 372181 524527 372215
rect 524527 372181 524553 372215
rect 524591 372181 524595 372215
rect 524595 372181 524625 372215
rect 524663 372181 524697 372215
rect 513771 371953 513805 371987
rect 513771 371753 513805 371787
rect 513771 371553 513805 371587
rect 513771 371353 513805 371387
rect 513771 371153 513805 371187
rect 513771 370953 513805 370987
rect 513771 370753 513805 370787
rect 513771 370553 513805 370587
rect 513771 370353 513805 370387
rect 513771 370153 513805 370187
rect 513771 369953 513805 369987
rect 513771 369753 513805 369787
rect 515651 371855 515685 371889
rect 515651 371655 515685 371689
rect 515919 371659 516457 372053
rect 516879 371659 517417 372053
rect 517531 371855 517565 371889
rect 517531 371655 517565 371689
rect 515651 371455 515685 371489
rect 515651 371255 515685 371289
rect 517531 371455 517565 371489
rect 517531 371255 517565 371289
rect 515651 371055 515685 371089
rect 515651 370855 515685 370889
rect 515651 370655 515685 370689
rect 517531 371055 517565 371089
rect 517531 370855 517565 370889
rect 517531 370655 517565 370689
rect 515651 370455 515685 370489
rect 515651 370255 515685 370289
rect 515651 370055 515685 370089
rect 517531 370455 517565 370489
rect 517531 370255 517565 370289
rect 515651 369855 515685 369889
rect 515919 369652 516457 370046
rect 516879 369652 517417 370046
rect 517531 370055 517565 370089
rect 517531 369855 517565 369889
rect 523171 371907 523205 371941
rect 523171 371507 523205 371541
rect 523171 371107 523205 371141
rect 523439 371723 523473 371757
rect 523511 371723 523541 371757
rect 523541 371723 523545 371757
rect 523583 371723 523609 371757
rect 523609 371723 523617 371757
rect 523655 371723 523677 371757
rect 523677 371723 523689 371757
rect 523727 371723 523745 371757
rect 523745 371723 523761 371757
rect 523799 371723 523813 371757
rect 523813 371723 523833 371757
rect 523871 371723 523881 371757
rect 523881 371723 523905 371757
rect 523943 371723 523949 371757
rect 523949 371723 523977 371757
rect 524015 371723 524017 371757
rect 524017 371723 524049 371757
rect 524087 371723 524119 371757
rect 524119 371723 524121 371757
rect 524159 371723 524187 371757
rect 524187 371723 524193 371757
rect 524231 371723 524255 371757
rect 524255 371723 524265 371757
rect 524303 371723 524323 371757
rect 524323 371723 524337 371757
rect 524375 371723 524391 371757
rect 524391 371723 524409 371757
rect 524447 371723 524459 371757
rect 524459 371723 524481 371757
rect 524519 371723 524527 371757
rect 524527 371723 524553 371757
rect 524591 371723 524595 371757
rect 524595 371723 524625 371757
rect 524663 371723 524697 371757
rect 523439 371265 523473 371299
rect 523511 371265 523541 371299
rect 523541 371265 523545 371299
rect 523583 371265 523609 371299
rect 523609 371265 523617 371299
rect 523655 371265 523677 371299
rect 523677 371265 523689 371299
rect 523727 371265 523745 371299
rect 523745 371265 523761 371299
rect 523799 371265 523813 371299
rect 523813 371265 523833 371299
rect 523871 371265 523881 371299
rect 523881 371265 523905 371299
rect 523943 371265 523949 371299
rect 523949 371265 523977 371299
rect 524015 371265 524017 371299
rect 524017 371265 524049 371299
rect 524087 371265 524119 371299
rect 524119 371265 524121 371299
rect 524159 371265 524187 371299
rect 524187 371265 524193 371299
rect 524231 371265 524255 371299
rect 524255 371265 524265 371299
rect 524303 371265 524323 371299
rect 524323 371265 524337 371299
rect 524375 371265 524391 371299
rect 524391 371265 524409 371299
rect 524447 371265 524459 371299
rect 524459 371265 524481 371299
rect 524519 371265 524527 371299
rect 524527 371265 524553 371299
rect 524591 371265 524595 371299
rect 524595 371265 524625 371299
rect 524663 371265 524697 371299
rect 523171 370707 523205 370741
rect 523171 370307 523205 370341
rect 523171 369907 523205 369941
rect 523439 370807 523473 370841
rect 523511 370807 523541 370841
rect 523541 370807 523545 370841
rect 523583 370807 523609 370841
rect 523609 370807 523617 370841
rect 523655 370807 523677 370841
rect 523677 370807 523689 370841
rect 523727 370807 523745 370841
rect 523745 370807 523761 370841
rect 523799 370807 523813 370841
rect 523813 370807 523833 370841
rect 523871 370807 523881 370841
rect 523881 370807 523905 370841
rect 523943 370807 523949 370841
rect 523949 370807 523977 370841
rect 524015 370807 524017 370841
rect 524017 370807 524049 370841
rect 524087 370807 524119 370841
rect 524119 370807 524121 370841
rect 524159 370807 524187 370841
rect 524187 370807 524193 370841
rect 524231 370807 524255 370841
rect 524255 370807 524265 370841
rect 524303 370807 524323 370841
rect 524323 370807 524337 370841
rect 524375 370807 524391 370841
rect 524391 370807 524409 370841
rect 524447 370807 524459 370841
rect 524459 370807 524481 370841
rect 524519 370807 524527 370841
rect 524527 370807 524553 370841
rect 524591 370807 524595 370841
rect 524595 370807 524625 370841
rect 524663 370807 524697 370841
rect 523439 370349 523473 370383
rect 523511 370349 523541 370383
rect 523541 370349 523545 370383
rect 523583 370349 523609 370383
rect 523609 370349 523617 370383
rect 523655 370349 523677 370383
rect 523677 370349 523689 370383
rect 523727 370349 523745 370383
rect 523745 370349 523761 370383
rect 523799 370349 523813 370383
rect 523813 370349 523833 370383
rect 523871 370349 523881 370383
rect 523881 370349 523905 370383
rect 523943 370349 523949 370383
rect 523949 370349 523977 370383
rect 524015 370349 524017 370383
rect 524017 370349 524049 370383
rect 524087 370349 524119 370383
rect 524119 370349 524121 370383
rect 524159 370349 524187 370383
rect 524187 370349 524193 370383
rect 524231 370349 524255 370383
rect 524255 370349 524265 370383
rect 524303 370349 524323 370383
rect 524323 370349 524337 370383
rect 524375 370349 524391 370383
rect 524391 370349 524409 370383
rect 524447 370349 524459 370383
rect 524459 370349 524481 370383
rect 524519 370349 524527 370383
rect 524527 370349 524553 370383
rect 524591 370349 524595 370383
rect 524595 370349 524625 370383
rect 524663 370349 524697 370383
rect 513771 369553 513805 369587
rect 513771 369353 513805 369387
rect 523171 369507 523205 369541
rect 513771 369153 513805 369187
rect 513771 368953 513805 368987
rect 513771 368753 513805 368787
rect 513771 368553 513805 368587
rect 513771 368353 513805 368387
rect 513771 368153 513805 368187
rect 513771 367953 513805 367987
rect 513771 367753 513805 367787
rect 513771 367553 513805 367587
rect 513771 367353 513805 367387
rect 513771 367153 513805 367187
rect 513771 366953 513805 366987
rect 515651 369111 515685 369145
rect 515651 368911 515685 368945
rect 515919 368915 516457 369309
rect 516879 368915 517417 369309
rect 517531 369111 517565 369145
rect 517531 368911 517565 368945
rect 515651 368711 515685 368745
rect 515651 368511 515685 368545
rect 517531 368711 517565 368745
rect 517531 368511 517565 368545
rect 515651 368311 515685 368345
rect 515651 368111 515685 368145
rect 515651 367911 515685 367945
rect 517531 368311 517565 368345
rect 517531 368111 517565 368145
rect 517531 367911 517565 367945
rect 515651 367711 515685 367745
rect 515651 367511 515685 367545
rect 515651 367311 515685 367345
rect 517531 367711 517565 367745
rect 517531 367511 517565 367545
rect 515651 367111 515685 367145
rect 515919 366908 516457 367302
rect 516879 366908 517417 367302
rect 517531 367311 517565 367345
rect 517531 367111 517565 367145
rect 523171 369107 523205 369141
rect 523171 368707 523205 368741
rect 523439 369891 523473 369925
rect 523511 369891 523541 369925
rect 523541 369891 523545 369925
rect 523583 369891 523609 369925
rect 523609 369891 523617 369925
rect 523655 369891 523677 369925
rect 523677 369891 523689 369925
rect 523727 369891 523745 369925
rect 523745 369891 523761 369925
rect 523799 369891 523813 369925
rect 523813 369891 523833 369925
rect 523871 369891 523881 369925
rect 523881 369891 523905 369925
rect 523943 369891 523949 369925
rect 523949 369891 523977 369925
rect 524015 369891 524017 369925
rect 524017 369891 524049 369925
rect 524087 369891 524119 369925
rect 524119 369891 524121 369925
rect 524159 369891 524187 369925
rect 524187 369891 524193 369925
rect 524231 369891 524255 369925
rect 524255 369891 524265 369925
rect 524303 369891 524323 369925
rect 524323 369891 524337 369925
rect 524375 369891 524391 369925
rect 524391 369891 524409 369925
rect 524447 369891 524459 369925
rect 524459 369891 524481 369925
rect 524519 369891 524527 369925
rect 524527 369891 524553 369925
rect 524591 369891 524595 369925
rect 524595 369891 524625 369925
rect 524663 369891 524697 369925
rect 523439 369433 523473 369467
rect 523511 369433 523541 369467
rect 523541 369433 523545 369467
rect 523583 369433 523609 369467
rect 523609 369433 523617 369467
rect 523655 369433 523677 369467
rect 523677 369433 523689 369467
rect 523727 369433 523745 369467
rect 523745 369433 523761 369467
rect 523799 369433 523813 369467
rect 523813 369433 523833 369467
rect 523871 369433 523881 369467
rect 523881 369433 523905 369467
rect 523943 369433 523949 369467
rect 523949 369433 523977 369467
rect 524015 369433 524017 369467
rect 524017 369433 524049 369467
rect 524087 369433 524119 369467
rect 524119 369433 524121 369467
rect 524159 369433 524187 369467
rect 524187 369433 524193 369467
rect 524231 369433 524255 369467
rect 524255 369433 524265 369467
rect 524303 369433 524323 369467
rect 524323 369433 524337 369467
rect 524375 369433 524391 369467
rect 524391 369433 524409 369467
rect 524447 369433 524459 369467
rect 524459 369433 524481 369467
rect 524519 369433 524527 369467
rect 524527 369433 524553 369467
rect 524591 369433 524595 369467
rect 524595 369433 524625 369467
rect 524663 369433 524697 369467
rect 523439 368975 523473 369009
rect 523511 368975 523541 369009
rect 523541 368975 523545 369009
rect 523583 368975 523609 369009
rect 523609 368975 523617 369009
rect 523655 368975 523677 369009
rect 523677 368975 523689 369009
rect 523727 368975 523745 369009
rect 523745 368975 523761 369009
rect 523799 368975 523813 369009
rect 523813 368975 523833 369009
rect 523871 368975 523881 369009
rect 523881 368975 523905 369009
rect 523943 368975 523949 369009
rect 523949 368975 523977 369009
rect 524015 368975 524017 369009
rect 524017 368975 524049 369009
rect 524087 368975 524119 369009
rect 524119 368975 524121 369009
rect 524159 368975 524187 369009
rect 524187 368975 524193 369009
rect 524231 368975 524255 369009
rect 524255 368975 524265 369009
rect 524303 368975 524323 369009
rect 524323 368975 524337 369009
rect 524375 368975 524391 369009
rect 524391 368975 524409 369009
rect 524447 368975 524459 369009
rect 524459 368975 524481 369009
rect 524519 368975 524527 369009
rect 524527 368975 524553 369009
rect 524591 368975 524595 369009
rect 524595 368975 524625 369009
rect 524663 368975 524697 369009
rect 523439 368517 523473 368551
rect 523511 368517 523541 368551
rect 523541 368517 523545 368551
rect 523583 368517 523609 368551
rect 523609 368517 523617 368551
rect 523655 368517 523677 368551
rect 523677 368517 523689 368551
rect 523727 368517 523745 368551
rect 523745 368517 523761 368551
rect 523799 368517 523813 368551
rect 523813 368517 523833 368551
rect 523871 368517 523881 368551
rect 523881 368517 523905 368551
rect 523943 368517 523949 368551
rect 523949 368517 523977 368551
rect 524015 368517 524017 368551
rect 524017 368517 524049 368551
rect 524087 368517 524119 368551
rect 524119 368517 524121 368551
rect 524159 368517 524187 368551
rect 524187 368517 524193 368551
rect 524231 368517 524255 368551
rect 524255 368517 524265 368551
rect 524303 368517 524323 368551
rect 524323 368517 524337 368551
rect 524375 368517 524391 368551
rect 524391 368517 524409 368551
rect 524447 368517 524459 368551
rect 524459 368517 524481 368551
rect 524519 368517 524527 368551
rect 524527 368517 524553 368551
rect 524591 368517 524595 368551
rect 524595 368517 524625 368551
rect 524663 368517 524697 368551
rect 523171 368307 523205 368341
rect 523171 367907 523205 367941
rect 523171 367507 523205 367541
rect 523171 367107 523205 367141
rect 523439 368059 523473 368093
rect 523511 368059 523541 368093
rect 523541 368059 523545 368093
rect 523583 368059 523609 368093
rect 523609 368059 523617 368093
rect 523655 368059 523677 368093
rect 523677 368059 523689 368093
rect 523727 368059 523745 368093
rect 523745 368059 523761 368093
rect 523799 368059 523813 368093
rect 523813 368059 523833 368093
rect 523871 368059 523881 368093
rect 523881 368059 523905 368093
rect 523943 368059 523949 368093
rect 523949 368059 523977 368093
rect 524015 368059 524017 368093
rect 524017 368059 524049 368093
rect 524087 368059 524119 368093
rect 524119 368059 524121 368093
rect 524159 368059 524187 368093
rect 524187 368059 524193 368093
rect 524231 368059 524255 368093
rect 524255 368059 524265 368093
rect 524303 368059 524323 368093
rect 524323 368059 524337 368093
rect 524375 368059 524391 368093
rect 524391 368059 524409 368093
rect 524447 368059 524459 368093
rect 524459 368059 524481 368093
rect 524519 368059 524527 368093
rect 524527 368059 524553 368093
rect 524591 368059 524595 368093
rect 524595 368059 524625 368093
rect 524663 368059 524697 368093
rect 523439 367601 523473 367635
rect 523511 367601 523541 367635
rect 523541 367601 523545 367635
rect 523583 367601 523609 367635
rect 523609 367601 523617 367635
rect 523655 367601 523677 367635
rect 523677 367601 523689 367635
rect 523727 367601 523745 367635
rect 523745 367601 523761 367635
rect 523799 367601 523813 367635
rect 523813 367601 523833 367635
rect 523871 367601 523881 367635
rect 523881 367601 523905 367635
rect 523943 367601 523949 367635
rect 523949 367601 523977 367635
rect 524015 367601 524017 367635
rect 524017 367601 524049 367635
rect 524087 367601 524119 367635
rect 524119 367601 524121 367635
rect 524159 367601 524187 367635
rect 524187 367601 524193 367635
rect 524231 367601 524255 367635
rect 524255 367601 524265 367635
rect 524303 367601 524323 367635
rect 524323 367601 524337 367635
rect 524375 367601 524391 367635
rect 524391 367601 524409 367635
rect 524447 367601 524459 367635
rect 524459 367601 524481 367635
rect 524519 367601 524527 367635
rect 524527 367601 524553 367635
rect 524591 367601 524595 367635
rect 524595 367601 524625 367635
rect 524663 367601 524697 367635
rect 513771 366753 513805 366787
rect 513771 366553 513805 366587
rect 523171 366707 523205 366741
rect 513771 366353 513805 366387
rect 513771 366153 513805 366187
rect 513771 365953 513805 365987
rect 513771 365753 513805 365787
rect 513771 365553 513805 365587
rect 513771 365353 513805 365387
rect 513771 365153 513805 365187
rect 513771 364953 513805 364987
rect 513771 364753 513805 364787
rect 513771 364553 513805 364587
rect 513771 364353 513805 364387
rect 513771 364153 513805 364187
rect 515651 366367 515685 366401
rect 515651 366167 515685 366201
rect 515919 366171 516457 366565
rect 516879 366171 517417 366565
rect 517531 366367 517565 366401
rect 517531 366167 517565 366201
rect 515651 365967 515685 366001
rect 515651 365767 515685 365801
rect 517531 365967 517565 366001
rect 517531 365767 517565 365801
rect 515651 365567 515685 365601
rect 515651 365367 515685 365401
rect 515651 365167 515685 365201
rect 517531 365567 517565 365601
rect 517531 365367 517565 365401
rect 517531 365167 517565 365201
rect 515651 364967 515685 365001
rect 515651 364767 515685 364801
rect 515651 364567 515685 364601
rect 517531 364967 517565 365001
rect 517531 364767 517565 364801
rect 515651 364367 515685 364401
rect 515919 364164 516457 364558
rect 516879 364164 517417 364558
rect 517531 364567 517565 364601
rect 517531 364367 517565 364401
rect 519411 366367 519445 366401
rect 519411 366167 519445 366201
rect 519679 366171 520217 366565
rect 520639 366171 521177 366565
rect 521291 366367 521325 366401
rect 521291 366167 521325 366201
rect 519411 365967 519445 366001
rect 519411 365767 519445 365801
rect 521291 365967 521325 366001
rect 521291 365767 521325 365801
rect 519411 365567 519445 365601
rect 519411 365367 519445 365401
rect 519411 365167 519445 365201
rect 521291 365567 521325 365601
rect 521291 365367 521325 365401
rect 521291 365167 521325 365201
rect 519411 364967 519445 365001
rect 519411 364767 519445 364801
rect 519411 364567 519445 364601
rect 521291 364967 521325 365001
rect 521291 364767 521325 364801
rect 519411 364367 519445 364401
rect 519679 364164 520217 364558
rect 520639 364164 521177 364558
rect 521291 364567 521325 364601
rect 521291 364367 521325 364401
rect 523171 366307 523205 366341
rect 523171 365907 523205 365941
rect 523439 367143 523473 367177
rect 523511 367143 523541 367177
rect 523541 367143 523545 367177
rect 523583 367143 523609 367177
rect 523609 367143 523617 367177
rect 523655 367143 523677 367177
rect 523677 367143 523689 367177
rect 523727 367143 523745 367177
rect 523745 367143 523761 367177
rect 523799 367143 523813 367177
rect 523813 367143 523833 367177
rect 523871 367143 523881 367177
rect 523881 367143 523905 367177
rect 523943 367143 523949 367177
rect 523949 367143 523977 367177
rect 524015 367143 524017 367177
rect 524017 367143 524049 367177
rect 524087 367143 524119 367177
rect 524119 367143 524121 367177
rect 524159 367143 524187 367177
rect 524187 367143 524193 367177
rect 524231 367143 524255 367177
rect 524255 367143 524265 367177
rect 524303 367143 524323 367177
rect 524323 367143 524337 367177
rect 524375 367143 524391 367177
rect 524391 367143 524409 367177
rect 524447 367143 524459 367177
rect 524459 367143 524481 367177
rect 524519 367143 524527 367177
rect 524527 367143 524553 367177
rect 524591 367143 524595 367177
rect 524595 367143 524625 367177
rect 524663 367143 524697 367177
rect 523439 366685 523473 366719
rect 523511 366685 523541 366719
rect 523541 366685 523545 366719
rect 523583 366685 523609 366719
rect 523609 366685 523617 366719
rect 523655 366685 523677 366719
rect 523677 366685 523689 366719
rect 523727 366685 523745 366719
rect 523745 366685 523761 366719
rect 523799 366685 523813 366719
rect 523813 366685 523833 366719
rect 523871 366685 523881 366719
rect 523881 366685 523905 366719
rect 523943 366685 523949 366719
rect 523949 366685 523977 366719
rect 524015 366685 524017 366719
rect 524017 366685 524049 366719
rect 524087 366685 524119 366719
rect 524119 366685 524121 366719
rect 524159 366685 524187 366719
rect 524187 366685 524193 366719
rect 524231 366685 524255 366719
rect 524255 366685 524265 366719
rect 524303 366685 524323 366719
rect 524323 366685 524337 366719
rect 524375 366685 524391 366719
rect 524391 366685 524409 366719
rect 524447 366685 524459 366719
rect 524459 366685 524481 366719
rect 524519 366685 524527 366719
rect 524527 366685 524553 366719
rect 524591 366685 524595 366719
rect 524595 366685 524625 366719
rect 524663 366685 524697 366719
rect 523439 366227 523473 366261
rect 523511 366227 523541 366261
rect 523541 366227 523545 366261
rect 523583 366227 523609 366261
rect 523609 366227 523617 366261
rect 523655 366227 523677 366261
rect 523677 366227 523689 366261
rect 523727 366227 523745 366261
rect 523745 366227 523761 366261
rect 523799 366227 523813 366261
rect 523813 366227 523833 366261
rect 523871 366227 523881 366261
rect 523881 366227 523905 366261
rect 523943 366227 523949 366261
rect 523949 366227 523977 366261
rect 524015 366227 524017 366261
rect 524017 366227 524049 366261
rect 524087 366227 524119 366261
rect 524119 366227 524121 366261
rect 524159 366227 524187 366261
rect 524187 366227 524193 366261
rect 524231 366227 524255 366261
rect 524255 366227 524265 366261
rect 524303 366227 524323 366261
rect 524323 366227 524337 366261
rect 524375 366227 524391 366261
rect 524391 366227 524409 366261
rect 524447 366227 524459 366261
rect 524459 366227 524481 366261
rect 524519 366227 524527 366261
rect 524527 366227 524553 366261
rect 524591 366227 524595 366261
rect 524595 366227 524625 366261
rect 524663 366227 524697 366261
rect 523439 365769 523473 365803
rect 523511 365769 523541 365803
rect 523541 365769 523545 365803
rect 523583 365769 523609 365803
rect 523609 365769 523617 365803
rect 523655 365769 523677 365803
rect 523677 365769 523689 365803
rect 523727 365769 523745 365803
rect 523745 365769 523761 365803
rect 523799 365769 523813 365803
rect 523813 365769 523833 365803
rect 523871 365769 523881 365803
rect 523881 365769 523905 365803
rect 523943 365769 523949 365803
rect 523949 365769 523977 365803
rect 524015 365769 524017 365803
rect 524017 365769 524049 365803
rect 524087 365769 524119 365803
rect 524119 365769 524121 365803
rect 524159 365769 524187 365803
rect 524187 365769 524193 365803
rect 524231 365769 524255 365803
rect 524255 365769 524265 365803
rect 524303 365769 524323 365803
rect 524323 365769 524337 365803
rect 524375 365769 524391 365803
rect 524391 365769 524409 365803
rect 524447 365769 524459 365803
rect 524459 365769 524481 365803
rect 524519 365769 524527 365803
rect 524527 365769 524553 365803
rect 524591 365769 524595 365803
rect 524595 365769 524625 365803
rect 524663 365769 524697 365803
rect 523171 365507 523205 365541
rect 523171 365107 523205 365141
rect 523171 364707 523205 364741
rect 523439 365311 523473 365345
rect 523511 365311 523541 365345
rect 523541 365311 523545 365345
rect 523583 365311 523609 365345
rect 523609 365311 523617 365345
rect 523655 365311 523677 365345
rect 523677 365311 523689 365345
rect 523727 365311 523745 365345
rect 523745 365311 523761 365345
rect 523799 365311 523813 365345
rect 523813 365311 523833 365345
rect 523871 365311 523881 365345
rect 523881 365311 523905 365345
rect 523943 365311 523949 365345
rect 523949 365311 523977 365345
rect 524015 365311 524017 365345
rect 524017 365311 524049 365345
rect 524087 365311 524119 365345
rect 524119 365311 524121 365345
rect 524159 365311 524187 365345
rect 524187 365311 524193 365345
rect 524231 365311 524255 365345
rect 524255 365311 524265 365345
rect 524303 365311 524323 365345
rect 524323 365311 524337 365345
rect 524375 365311 524391 365345
rect 524391 365311 524409 365345
rect 524447 365311 524459 365345
rect 524459 365311 524481 365345
rect 524519 365311 524527 365345
rect 524527 365311 524553 365345
rect 524591 365311 524595 365345
rect 524595 365311 524625 365345
rect 524663 365311 524697 365345
rect 523439 364853 523473 364887
rect 523511 364853 523541 364887
rect 523541 364853 523545 364887
rect 523583 364853 523609 364887
rect 523609 364853 523617 364887
rect 523655 364853 523677 364887
rect 523677 364853 523689 364887
rect 523727 364853 523745 364887
rect 523745 364853 523761 364887
rect 523799 364853 523813 364887
rect 523813 364853 523833 364887
rect 523871 364853 523881 364887
rect 523881 364853 523905 364887
rect 523943 364853 523949 364887
rect 523949 364853 523977 364887
rect 524015 364853 524017 364887
rect 524017 364853 524049 364887
rect 524087 364853 524119 364887
rect 524119 364853 524121 364887
rect 524159 364853 524187 364887
rect 524187 364853 524193 364887
rect 524231 364853 524255 364887
rect 524255 364853 524265 364887
rect 524303 364853 524323 364887
rect 524323 364853 524337 364887
rect 524375 364853 524391 364887
rect 524391 364853 524409 364887
rect 524447 364853 524459 364887
rect 524459 364853 524481 364887
rect 524519 364853 524527 364887
rect 524527 364853 524553 364887
rect 524591 364853 524595 364887
rect 524595 364853 524625 364887
rect 524663 364853 524697 364887
rect 523171 364307 523205 364341
rect 513771 363953 513805 363987
rect 513771 363753 513805 363787
rect 513771 363553 513805 363587
rect 513771 363353 513805 363387
rect 513771 363153 513805 363187
rect 513771 362953 513805 362987
rect 513771 362753 513805 362787
rect 513771 362553 513805 362587
rect 523171 363907 523205 363941
rect 523171 363507 523205 363541
rect 523171 363107 523205 363141
rect 523171 362707 523205 362741
rect 523439 364395 523473 364429
rect 523511 364395 523541 364429
rect 523541 364395 523545 364429
rect 523583 364395 523609 364429
rect 523609 364395 523617 364429
rect 523655 364395 523677 364429
rect 523677 364395 523689 364429
rect 523727 364395 523745 364429
rect 523745 364395 523761 364429
rect 523799 364395 523813 364429
rect 523813 364395 523833 364429
rect 523871 364395 523881 364429
rect 523881 364395 523905 364429
rect 523943 364395 523949 364429
rect 523949 364395 523977 364429
rect 524015 364395 524017 364429
rect 524017 364395 524049 364429
rect 524087 364395 524119 364429
rect 524119 364395 524121 364429
rect 524159 364395 524187 364429
rect 524187 364395 524193 364429
rect 524231 364395 524255 364429
rect 524255 364395 524265 364429
rect 524303 364395 524323 364429
rect 524323 364395 524337 364429
rect 524375 364395 524391 364429
rect 524391 364395 524409 364429
rect 524447 364395 524459 364429
rect 524459 364395 524481 364429
rect 524519 364395 524527 364429
rect 524527 364395 524553 364429
rect 524591 364395 524595 364429
rect 524595 364395 524625 364429
rect 524663 364395 524697 364429
rect 523439 363937 523473 363971
rect 523511 363937 523541 363971
rect 523541 363937 523545 363971
rect 523583 363937 523609 363971
rect 523609 363937 523617 363971
rect 523655 363937 523677 363971
rect 523677 363937 523689 363971
rect 523727 363937 523745 363971
rect 523745 363937 523761 363971
rect 523799 363937 523813 363971
rect 523813 363937 523833 363971
rect 523871 363937 523881 363971
rect 523881 363937 523905 363971
rect 523943 363937 523949 363971
rect 523949 363937 523977 363971
rect 524015 363937 524017 363971
rect 524017 363937 524049 363971
rect 524087 363937 524119 363971
rect 524119 363937 524121 363971
rect 524159 363937 524187 363971
rect 524187 363937 524193 363971
rect 524231 363937 524255 363971
rect 524255 363937 524265 363971
rect 524303 363937 524323 363971
rect 524323 363937 524337 363971
rect 524375 363937 524391 363971
rect 524391 363937 524409 363971
rect 524447 363937 524459 363971
rect 524459 363937 524481 363971
rect 524519 363937 524527 363971
rect 524527 363937 524553 363971
rect 524591 363937 524595 363971
rect 524595 363937 524625 363971
rect 524663 363937 524697 363971
rect 523439 363479 523473 363513
rect 523511 363479 523541 363513
rect 523541 363479 523545 363513
rect 523583 363479 523609 363513
rect 523609 363479 523617 363513
rect 523655 363479 523677 363513
rect 523677 363479 523689 363513
rect 523727 363479 523745 363513
rect 523745 363479 523761 363513
rect 523799 363479 523813 363513
rect 523813 363479 523833 363513
rect 523871 363479 523881 363513
rect 523881 363479 523905 363513
rect 523943 363479 523949 363513
rect 523949 363479 523977 363513
rect 524015 363479 524017 363513
rect 524017 363479 524049 363513
rect 524087 363479 524119 363513
rect 524119 363479 524121 363513
rect 524159 363479 524187 363513
rect 524187 363479 524193 363513
rect 524231 363479 524255 363513
rect 524255 363479 524265 363513
rect 524303 363479 524323 363513
rect 524323 363479 524337 363513
rect 524375 363479 524391 363513
rect 524391 363479 524409 363513
rect 524447 363479 524459 363513
rect 524459 363479 524481 363513
rect 524519 363479 524527 363513
rect 524527 363479 524553 363513
rect 524591 363479 524595 363513
rect 524595 363479 524625 363513
rect 524663 363479 524697 363513
rect 523439 363021 523473 363055
rect 523511 363021 523541 363055
rect 523541 363021 523545 363055
rect 523583 363021 523609 363055
rect 523609 363021 523617 363055
rect 523655 363021 523677 363055
rect 523677 363021 523689 363055
rect 523727 363021 523745 363055
rect 523745 363021 523761 363055
rect 523799 363021 523813 363055
rect 523813 363021 523833 363055
rect 523871 363021 523881 363055
rect 523881 363021 523905 363055
rect 523943 363021 523949 363055
rect 523949 363021 523977 363055
rect 524015 363021 524017 363055
rect 524017 363021 524049 363055
rect 524087 363021 524119 363055
rect 524119 363021 524121 363055
rect 524159 363021 524187 363055
rect 524187 363021 524193 363055
rect 524231 363021 524255 363055
rect 524255 363021 524265 363055
rect 524303 363021 524323 363055
rect 524323 363021 524337 363055
rect 524375 363021 524391 363055
rect 524391 363021 524409 363055
rect 524447 363021 524459 363055
rect 524459 363021 524481 363055
rect 524519 363021 524527 363055
rect 524527 363021 524553 363055
rect 524591 363021 524595 363055
rect 524595 363021 524625 363055
rect 524663 363021 524697 363055
rect 523439 362563 523473 362597
rect 523511 362563 523541 362597
rect 523541 362563 523545 362597
rect 523583 362563 523609 362597
rect 523609 362563 523617 362597
rect 523655 362563 523677 362597
rect 523677 362563 523689 362597
rect 523727 362563 523745 362597
rect 523745 362563 523761 362597
rect 523799 362563 523813 362597
rect 523813 362563 523833 362597
rect 523871 362563 523881 362597
rect 523881 362563 523905 362597
rect 523943 362563 523949 362597
rect 523949 362563 523977 362597
rect 524015 362563 524017 362597
rect 524017 362563 524049 362597
rect 524087 362563 524119 362597
rect 524119 362563 524121 362597
rect 524159 362563 524187 362597
rect 524187 362563 524193 362597
rect 524231 362563 524255 362597
rect 524255 362563 524265 362597
rect 524303 362563 524323 362597
rect 524323 362563 524337 362597
rect 524375 362563 524391 362597
rect 524391 362563 524409 362597
rect 524447 362563 524459 362597
rect 524459 362563 524481 362597
rect 524519 362563 524527 362597
rect 524527 362563 524553 362597
rect 524591 362563 524595 362597
rect 524595 362563 524625 362597
rect 524663 362563 524697 362597
rect 524907 389507 524917 389533
rect 524917 389507 524941 389533
rect 524907 389499 524941 389507
rect 525051 389907 525085 389941
rect 525051 389507 525085 389541
rect 525051 389107 525085 389141
rect 525051 388707 525085 388741
rect 525051 388307 525085 388341
rect 525051 387907 525085 387941
rect 525051 387507 525085 387541
rect 525051 387107 525085 387141
rect 525051 386707 525085 386741
rect 525051 386307 525085 386341
rect 525051 385907 525085 385941
rect 525051 385507 525085 385541
rect 525051 385107 525085 385141
rect 525051 384707 525085 384741
rect 525051 384307 525085 384341
rect 525051 383907 525085 383941
rect 525051 383507 525085 383541
rect 525051 383107 525085 383141
rect 525051 382707 525085 382741
rect 525051 382307 525085 382341
rect 525051 381907 525085 381941
rect 525051 381507 525085 381541
rect 525051 381107 525085 381141
rect 525051 380707 525085 380741
rect 525051 380307 525085 380341
rect 525051 379907 525085 379941
rect 525051 379507 525085 379541
rect 525051 379107 525085 379141
rect 525051 378707 525085 378741
rect 525051 378307 525085 378341
rect 525051 377907 525085 377941
rect 525051 377507 525085 377541
rect 525051 377107 525085 377141
rect 525051 376707 525085 376741
rect 525051 376307 525085 376341
rect 525051 375907 525085 375941
rect 525051 375507 525085 375541
rect 525051 375107 525085 375141
rect 525051 374707 525085 374741
rect 525051 374307 525085 374341
rect 525051 373907 525085 373941
rect 525051 373507 525085 373541
rect 525051 373107 525085 373141
rect 525051 372707 525085 372741
rect 525051 372307 525085 372341
rect 525051 371907 525085 371941
rect 525051 371507 525085 371541
rect 525051 371107 525085 371141
rect 525051 370707 525085 370741
rect 525051 370307 525085 370341
rect 525051 369907 525085 369941
rect 525051 369507 525085 369541
rect 525051 369107 525085 369141
rect 525051 368707 525085 368741
rect 526931 370875 526965 370909
rect 526931 370675 526965 370709
rect 527199 370679 527737 371073
rect 528159 370679 528697 371073
rect 528811 370875 528845 370909
rect 528811 370675 528845 370709
rect 526931 370475 526965 370509
rect 526931 370275 526965 370309
rect 528811 370475 528845 370509
rect 528811 370275 528845 370309
rect 526931 370075 526965 370109
rect 526931 369875 526965 369909
rect 526931 369675 526965 369709
rect 528811 370075 528845 370109
rect 528811 369875 528845 369909
rect 528811 369675 528845 369709
rect 526931 369475 526965 369509
rect 526931 369275 526965 369309
rect 526931 369075 526965 369109
rect 528811 369475 528845 369509
rect 528811 369275 528845 369309
rect 526931 368875 526965 368909
rect 527199 368672 527737 369066
rect 528159 368672 528697 369066
rect 528811 369075 528845 369109
rect 528811 368875 528845 368909
rect 530691 370973 530725 371007
rect 530691 370773 530725 370807
rect 530959 370777 531497 371171
rect 531919 370777 532457 371171
rect 532571 370973 532605 371007
rect 532571 370773 532605 370807
rect 530691 370573 530725 370607
rect 530691 370373 530725 370407
rect 532571 370573 532605 370607
rect 532571 370373 532605 370407
rect 530691 370173 530725 370207
rect 530691 369973 530725 370007
rect 530691 369773 530725 369807
rect 532571 370173 532605 370207
rect 532571 369973 532605 370007
rect 532571 369773 532605 369807
rect 530691 369573 530725 369607
rect 530691 369373 530725 369407
rect 530691 369173 530725 369207
rect 532571 369573 532605 369607
rect 532571 369373 532605 369407
rect 530691 368973 530725 369007
rect 530959 368770 531497 369164
rect 531919 368770 532457 369164
rect 532571 369173 532605 369207
rect 532571 368973 532605 369007
rect 534451 370189 534485 370223
rect 534451 369989 534485 370023
rect 534719 369993 535257 370387
rect 535679 369993 536217 370387
rect 536331 370189 536365 370223
rect 536331 369989 536365 370023
rect 534451 369789 534485 369823
rect 534451 369589 534485 369623
rect 536331 369789 536365 369823
rect 536331 369589 536365 369623
rect 534451 369389 534485 369423
rect 534451 369189 534485 369223
rect 534451 368989 534485 369023
rect 536331 369389 536365 369423
rect 536331 369189 536365 369223
rect 536331 368989 536365 369023
rect 534451 368789 534485 368823
rect 534451 368589 534485 368623
rect 525051 368307 525085 368341
rect 525051 367907 525085 367941
rect 525051 367507 525085 367541
rect 525051 367107 525085 367141
rect 525051 366707 525085 366741
rect 525051 366307 525085 366341
rect 525051 365907 525085 365941
rect 526931 368131 526965 368165
rect 526931 367931 526965 367965
rect 527199 367935 527737 368329
rect 528159 367935 528697 368329
rect 528811 368131 528845 368165
rect 528811 367931 528845 367965
rect 526931 367731 526965 367765
rect 526931 367531 526965 367565
rect 528811 367731 528845 367765
rect 528811 367531 528845 367565
rect 526931 367331 526965 367365
rect 526931 367131 526965 367165
rect 526931 366931 526965 366965
rect 528811 367331 528845 367365
rect 528811 367131 528845 367165
rect 528811 366931 528845 366965
rect 526931 366731 526965 366765
rect 526931 366531 526965 366565
rect 526931 366331 526965 366365
rect 528811 366731 528845 366765
rect 528811 366531 528845 366565
rect 526931 366131 526965 366165
rect 527199 365928 527737 366322
rect 528159 365928 528697 366322
rect 528811 366331 528845 366365
rect 528811 366131 528845 366165
rect 530691 368229 530725 368263
rect 530691 368029 530725 368063
rect 530959 368033 531497 368427
rect 531919 368033 532457 368427
rect 532571 368229 532605 368263
rect 532571 368029 532605 368063
rect 530691 367829 530725 367863
rect 530691 367629 530725 367663
rect 534451 368389 534485 368423
rect 536331 368789 536365 368823
rect 536331 368589 536365 368623
rect 534451 368189 534485 368223
rect 534719 367986 535257 368380
rect 535679 367986 536217 368380
rect 536331 368389 536365 368423
rect 536331 368189 536365 368223
rect 532571 367829 532605 367863
rect 532571 367629 532605 367663
rect 530691 367429 530725 367463
rect 530691 367229 530725 367263
rect 530691 367029 530725 367063
rect 532571 367429 532605 367463
rect 532571 367229 532605 367263
rect 532571 367029 532605 367063
rect 530691 366829 530725 366863
rect 530691 366629 530725 366663
rect 530691 366429 530725 366463
rect 532571 366829 532605 366863
rect 532571 366629 532605 366663
rect 530691 366229 530725 366263
rect 530959 366026 531497 366420
rect 531919 366026 532457 366420
rect 532571 366429 532605 366463
rect 532571 366229 532605 366263
rect 534451 367445 534485 367479
rect 534451 367245 534485 367279
rect 534719 367249 535257 367643
rect 535679 367249 536217 367643
rect 536331 367445 536365 367479
rect 536331 367245 536365 367279
rect 534451 367045 534485 367079
rect 534451 366845 534485 366879
rect 536331 367045 536365 367079
rect 536331 366845 536365 366879
rect 534451 366645 534485 366679
rect 534451 366445 534485 366479
rect 534451 366245 534485 366279
rect 536331 366645 536365 366679
rect 536331 366445 536365 366479
rect 536331 366245 536365 366279
rect 534451 366045 534485 366079
rect 534451 365845 534485 365879
rect 525051 365507 525085 365541
rect 525051 365107 525085 365141
rect 525051 364707 525085 364741
rect 525051 364307 525085 364341
rect 525051 363907 525085 363941
rect 525051 363507 525085 363541
rect 526931 365387 526965 365421
rect 526931 365187 526965 365221
rect 527199 365191 527737 365585
rect 528159 365191 528697 365585
rect 528811 365387 528845 365421
rect 528811 365187 528845 365221
rect 526931 364987 526965 365021
rect 526931 364787 526965 364821
rect 528811 364987 528845 365021
rect 528811 364787 528845 364821
rect 526931 364587 526965 364621
rect 526931 364387 526965 364421
rect 526931 364187 526965 364221
rect 528811 364587 528845 364621
rect 528811 364387 528845 364421
rect 528811 364187 528845 364221
rect 526931 363987 526965 364021
rect 526931 363787 526965 363821
rect 526931 363587 526965 363621
rect 528811 363987 528845 364021
rect 528811 363787 528845 363821
rect 526931 363387 526965 363421
rect 527199 363184 527737 363578
rect 528159 363184 528697 363578
rect 528811 363587 528845 363621
rect 528811 363387 528845 363421
rect 530691 365485 530725 365519
rect 530691 365285 530725 365319
rect 530959 365289 531497 365683
rect 531919 365289 532457 365683
rect 532571 365485 532605 365519
rect 532571 365285 532605 365319
rect 530691 365085 530725 365119
rect 530691 364885 530725 364919
rect 534451 365645 534485 365679
rect 536331 366045 536365 366079
rect 536331 365845 536365 365879
rect 534451 365445 534485 365479
rect 534719 365242 535257 365636
rect 535679 365242 536217 365636
rect 536331 365645 536365 365679
rect 536331 365445 536365 365479
rect 532571 365085 532605 365119
rect 532571 364885 532605 364919
rect 530691 364685 530725 364719
rect 530691 364485 530725 364519
rect 530691 364285 530725 364319
rect 532571 364685 532605 364719
rect 532571 364485 532605 364519
rect 532571 364285 532605 364319
rect 530691 364085 530725 364119
rect 530691 363885 530725 363919
rect 530691 363685 530725 363719
rect 532571 364085 532605 364119
rect 532571 363885 532605 363919
rect 530691 363485 530725 363519
rect 530959 363282 531497 363676
rect 531919 363282 532457 363676
rect 532571 363685 532605 363719
rect 532571 363485 532605 363519
rect 534451 364701 534485 364735
rect 534451 364501 534485 364535
rect 534719 364505 535257 364899
rect 535679 364505 536217 364899
rect 536331 364701 536365 364735
rect 536331 364501 536365 364535
rect 534451 364301 534485 364335
rect 534451 364101 534485 364135
rect 536331 364301 536365 364335
rect 536331 364101 536365 364135
rect 534451 363901 534485 363935
rect 534451 363701 534485 363735
rect 534451 363501 534485 363535
rect 536331 363901 536365 363935
rect 536331 363701 536365 363735
rect 536331 363501 536365 363535
rect 534451 363301 534485 363335
rect 525051 363107 525085 363141
rect 525051 362707 525085 362741
rect 534451 363101 534485 363135
rect 534451 362901 534485 362935
rect 536331 363301 536365 363335
rect 536331 363101 536365 363135
rect 534451 362701 534485 362735
rect 534719 362498 535257 362892
rect 535679 362498 536217 362892
rect 536331 362901 536365 362935
rect 536331 362701 536365 362735
rect 560728 359330 560788 359390
rect 560928 359330 560988 359390
rect 561128 359330 561188 359390
rect 561328 359330 561388 359390
rect 561528 359330 561588 359390
rect 561728 359330 561788 359390
rect 561928 359330 561988 359390
rect 562128 359330 562188 359390
rect 562328 359330 562388 359390
rect 562528 359330 562588 359390
rect 562728 359330 562788 359390
rect 562928 359330 562988 359390
rect 563128 359330 563188 359390
rect 563328 359330 563388 359390
rect 563528 359330 563588 359390
rect 563728 359330 563788 359390
rect 563928 359330 563988 359390
rect 564128 359330 564188 359390
rect 564328 359330 564388 359390
rect 564528 359330 564588 359390
rect 564728 359330 564788 359390
rect 564928 359330 564988 359390
rect 565128 359330 565188 359390
rect 565328 359330 565388 359390
rect 565528 359330 565588 359390
rect 574702 359260 574762 359320
rect 574902 359260 574962 359320
rect 575102 359260 575162 359320
rect 575302 359260 575362 359320
rect 575502 359260 575562 359320
rect 575702 359260 575762 359320
rect 575902 359260 575962 359320
rect 576102 359260 576162 359320
rect 576302 359260 576362 359320
rect 576502 359260 576562 359320
rect 576702 359260 576762 359320
rect 576902 359260 576962 359320
rect 577102 359260 577162 359320
rect 577302 359260 577362 359320
rect 577502 359260 577562 359320
rect 577702 359260 577762 359320
rect 577902 359260 577962 359320
rect 578102 359260 578162 359320
rect 578302 359260 578362 359320
rect 578502 359260 578562 359320
rect 578702 359260 578762 359320
rect 578902 359260 578962 359320
rect 579102 359260 579162 359320
rect 579302 359260 579362 359320
rect 579502 359260 579562 359320
rect 579702 359260 579762 359320
rect 560232 357872 560364 358022
rect 560553 357992 560587 358968
rect 560811 357992 560845 358968
rect 561069 357992 561103 358968
rect 561327 357992 561361 358968
rect 561585 357992 561619 358968
rect 561843 357992 561877 358968
rect 562101 357992 562135 358968
rect 562359 357992 562393 358968
rect 562617 357992 562651 358968
rect 562875 357992 562909 358968
rect 563133 357992 563167 358968
rect 563391 357992 563425 358968
rect 563649 357992 563683 358968
rect 563907 357992 563941 358968
rect 564165 357992 564199 358968
rect 564423 357992 564457 358968
rect 564681 357992 564715 358968
rect 564939 357992 564973 358968
rect 565197 357992 565231 358968
rect 565455 357992 565489 358968
rect 565713 357992 565747 358968
rect 565966 357860 566126 357968
rect 574691 357922 574725 358898
rect 574949 357922 574983 358898
rect 575207 357922 575241 358898
rect 575465 357922 575499 358898
rect 575723 357922 575757 358898
rect 575981 357922 576015 358898
rect 576239 357922 576273 358898
rect 576497 357922 576531 358898
rect 576755 357922 576789 358898
rect 577013 357922 577047 358898
rect 577271 357922 577305 358898
rect 577529 357922 577563 358898
rect 577787 357922 577821 358898
rect 578045 357922 578079 358898
rect 578303 357922 578337 358898
rect 578561 357922 578595 358898
rect 578819 357922 578853 358898
rect 579077 357922 579111 358898
rect 579335 357922 579369 358898
rect 579593 357922 579627 358898
rect 579851 357922 579885 358898
rect 580016 357726 580106 357814
rect 574408 357576 574500 357680
rect 560728 357450 560788 357510
rect 560928 357450 560988 357510
rect 561128 357450 561188 357510
rect 561328 357450 561388 357510
rect 561528 357450 561588 357510
rect 561728 357450 561788 357510
rect 561928 357450 561988 357510
rect 562128 357450 562188 357510
rect 562328 357450 562388 357510
rect 562528 357450 562588 357510
rect 562728 357450 562788 357510
rect 562928 357450 562988 357510
rect 563128 357450 563188 357510
rect 563328 357450 563388 357510
rect 563528 357450 563588 357510
rect 563728 357450 563788 357510
rect 563928 357450 563988 357510
rect 564128 357450 564188 357510
rect 564328 357450 564388 357510
rect 564528 357450 564588 357510
rect 564728 357450 564788 357510
rect 564928 357450 564988 357510
rect 565128 357450 565188 357510
rect 565328 357450 565388 357510
rect 565528 357450 565588 357510
rect 574702 357380 574762 357440
rect 574902 357380 574962 357440
rect 575102 357380 575162 357440
rect 575302 357380 575362 357440
rect 575502 357380 575562 357440
rect 575702 357380 575762 357440
rect 575902 357380 575962 357440
rect 576102 357380 576162 357440
rect 576302 357380 576362 357440
rect 576502 357380 576562 357440
rect 576702 357380 576762 357440
rect 576902 357380 576962 357440
rect 577102 357380 577162 357440
rect 577302 357380 577362 357440
rect 577502 357380 577562 357440
rect 577702 357380 577762 357440
rect 577902 357380 577962 357440
rect 578102 357380 578162 357440
rect 578302 357380 578362 357440
rect 578502 357380 578562 357440
rect 578702 357380 578762 357440
rect 578902 357380 578962 357440
rect 579102 357380 579162 357440
rect 579302 357380 579362 357440
rect 579502 357380 579562 357440
rect 579702 357380 579762 357440
rect 575150 313092 575210 313152
rect 575350 313092 575410 313152
rect 575550 313092 575610 313152
rect 575750 313092 575810 313152
rect 575950 313092 576010 313152
rect 576150 313092 576210 313152
rect 576350 313092 576410 313152
rect 576550 313092 576610 313152
rect 576750 313092 576810 313152
rect 576950 313092 577010 313152
rect 577150 313092 577210 313152
rect 577350 313092 577410 313152
rect 577550 313092 577610 313152
rect 577750 313092 577810 313152
rect 577950 313092 578010 313152
rect 578150 313092 578210 313152
rect 578350 313092 578410 313152
rect 578550 313092 578610 313152
rect 578750 313092 578810 313152
rect 578950 313092 579010 313152
rect 579150 313092 579210 313152
rect 579350 313092 579410 313152
rect 579550 313092 579610 313152
rect 579750 313092 579810 313152
rect 579950 313092 580010 313152
rect 580150 313092 580210 313152
rect 560590 313022 560650 313082
rect 560790 313022 560850 313082
rect 560990 313022 561050 313082
rect 561190 313022 561250 313082
rect 561390 313022 561450 313082
rect 561590 313022 561650 313082
rect 561790 313022 561850 313082
rect 561990 313022 562050 313082
rect 562190 313022 562250 313082
rect 562390 313022 562450 313082
rect 562590 313022 562650 313082
rect 562790 313022 562850 313082
rect 562990 313022 563050 313082
rect 563190 313022 563250 313082
rect 563390 313022 563450 313082
rect 563590 313022 563650 313082
rect 563790 313022 563850 313082
rect 563990 313022 564050 313082
rect 564190 313022 564250 313082
rect 564390 313022 564450 313082
rect 564590 313022 564650 313082
rect 564790 313022 564850 313082
rect 564990 313022 565050 313082
rect 565190 313022 565250 313082
rect 565390 313022 565450 313082
rect 560094 311564 560226 311714
rect 560415 311684 560449 312660
rect 560673 311684 560707 312660
rect 560931 311684 560965 312660
rect 561189 311684 561223 312660
rect 561447 311684 561481 312660
rect 561705 311684 561739 312660
rect 561963 311684 561997 312660
rect 562221 311684 562255 312660
rect 562479 311684 562513 312660
rect 562737 311684 562771 312660
rect 562995 311684 563029 312660
rect 563253 311684 563287 312660
rect 563511 311684 563545 312660
rect 563769 311684 563803 312660
rect 564027 311684 564061 312660
rect 564285 311684 564319 312660
rect 564543 311684 564577 312660
rect 564801 311684 564835 312660
rect 565059 311684 565093 312660
rect 565317 311684 565351 312660
rect 565575 311684 565609 312660
rect 565828 311552 565988 311660
rect 575139 311754 575173 312730
rect 575397 311754 575431 312730
rect 575655 311754 575689 312730
rect 575913 311754 575947 312730
rect 576171 311754 576205 312730
rect 576429 311754 576463 312730
rect 576687 311754 576721 312730
rect 576945 311754 576979 312730
rect 577203 311754 577237 312730
rect 577461 311754 577495 312730
rect 577719 311754 577753 312730
rect 577977 311754 578011 312730
rect 578235 311754 578269 312730
rect 578493 311754 578527 312730
rect 578751 311754 578785 312730
rect 579009 311754 579043 312730
rect 579267 311754 579301 312730
rect 579525 311754 579559 312730
rect 579783 311754 579817 312730
rect 580041 311754 580075 312730
rect 580299 311754 580333 312730
rect 580464 311558 580554 311646
rect 574856 311408 574948 311512
rect 575150 311212 575210 311272
rect 575350 311212 575410 311272
rect 575550 311212 575610 311272
rect 575750 311212 575810 311272
rect 575950 311212 576010 311272
rect 576150 311212 576210 311272
rect 576350 311212 576410 311272
rect 576550 311212 576610 311272
rect 576750 311212 576810 311272
rect 576950 311212 577010 311272
rect 577150 311212 577210 311272
rect 577350 311212 577410 311272
rect 577550 311212 577610 311272
rect 577750 311212 577810 311272
rect 577950 311212 578010 311272
rect 578150 311212 578210 311272
rect 578350 311212 578410 311272
rect 578550 311212 578610 311272
rect 578750 311212 578810 311272
rect 578950 311212 579010 311272
rect 579150 311212 579210 311272
rect 579350 311212 579410 311272
rect 579550 311212 579610 311272
rect 579750 311212 579810 311272
rect 579950 311212 580010 311272
rect 580150 311212 580210 311272
rect 560590 311142 560650 311202
rect 560790 311142 560850 311202
rect 560990 311142 561050 311202
rect 561190 311142 561250 311202
rect 561390 311142 561450 311202
rect 561590 311142 561650 311202
rect 561790 311142 561850 311202
rect 561990 311142 562050 311202
rect 562190 311142 562250 311202
rect 562390 311142 562450 311202
rect 562590 311142 562650 311202
rect 562790 311142 562850 311202
rect 562990 311142 563050 311202
rect 563190 311142 563250 311202
rect 563390 311142 563450 311202
rect 563590 311142 563650 311202
rect 563790 311142 563850 311202
rect 563990 311142 564050 311202
rect 564190 311142 564250 311202
rect 564390 311142 564450 311202
rect 564590 311142 564650 311202
rect 564790 311142 564850 311202
rect 564990 311142 565050 311202
rect 565190 311142 565250 311202
rect 565390 311142 565450 311202
<< metal1 >>
rect 566176 494126 566186 494310
rect 566408 494126 566418 494310
rect 580846 494136 580856 494348
rect 581040 494136 581050 494348
rect 560650 493850 565964 493880
rect 560650 493790 560836 493850
rect 560896 493790 561036 493850
rect 561096 493790 561236 493850
rect 561296 493790 561436 493850
rect 561496 493790 561636 493850
rect 561696 493790 561836 493850
rect 561896 493790 562036 493850
rect 562096 493790 562236 493850
rect 562296 493790 562436 493850
rect 562496 493790 562636 493850
rect 562696 493790 562836 493850
rect 562896 493790 563036 493850
rect 563096 493790 563236 493850
rect 563296 493790 563436 493850
rect 563496 493790 563636 493850
rect 563696 493790 563836 493850
rect 563896 493790 564036 493850
rect 564096 493790 564236 493850
rect 564296 493790 564436 493850
rect 564496 493790 564636 493850
rect 564696 493790 564836 493850
rect 564896 493790 565036 493850
rect 565096 493790 565236 493850
rect 565296 493790 565436 493850
rect 565496 493790 565636 493850
rect 565696 493790 565964 493850
rect 560650 493760 565964 493790
rect 560655 493428 560701 493440
rect 559792 492536 560110 492554
rect 559792 492324 559802 492536
rect 560012 492512 560110 492536
rect 560012 492482 560486 492512
rect 560012 492332 560340 492482
rect 560472 492332 560486 492482
rect 560655 492452 560661 493428
rect 560695 492452 560701 493428
rect 560655 492440 560701 492452
rect 560913 493428 560959 493440
rect 560913 492452 560919 493428
rect 560953 492452 560959 493428
rect 560913 492440 560959 492452
rect 561171 493428 561217 493440
rect 561171 492452 561177 493428
rect 561211 492452 561217 493428
rect 561171 492440 561217 492452
rect 561429 493428 561475 493440
rect 561429 492452 561435 493428
rect 561469 492452 561475 493428
rect 561429 492440 561475 492452
rect 561687 493428 561733 493440
rect 561687 492452 561693 493428
rect 561727 492452 561733 493428
rect 561687 492440 561733 492452
rect 561945 493428 561991 493440
rect 561945 492452 561951 493428
rect 561985 492452 561991 493428
rect 561945 492440 561991 492452
rect 562203 493428 562249 493440
rect 562203 492452 562209 493428
rect 562243 492452 562249 493428
rect 562203 492440 562249 492452
rect 562461 493428 562507 493440
rect 562461 492452 562467 493428
rect 562501 492452 562507 493428
rect 562461 492440 562507 492452
rect 562719 493428 562765 493440
rect 562719 492452 562725 493428
rect 562759 492452 562765 493428
rect 562719 492440 562765 492452
rect 562977 493428 563023 493440
rect 562977 492452 562983 493428
rect 563017 492452 563023 493428
rect 562977 492440 563023 492452
rect 563235 493428 563281 493440
rect 563235 492452 563241 493428
rect 563275 492452 563281 493428
rect 563235 492440 563281 492452
rect 563493 493428 563539 493440
rect 563493 492452 563499 493428
rect 563533 492452 563539 493428
rect 563493 492440 563539 492452
rect 563751 493428 563797 493440
rect 563751 492452 563757 493428
rect 563791 492452 563797 493428
rect 563751 492440 563797 492452
rect 564009 493428 564055 493440
rect 564009 492452 564015 493428
rect 564049 492452 564055 493428
rect 564009 492440 564055 492452
rect 564267 493428 564313 493440
rect 564267 492452 564273 493428
rect 564307 492452 564313 493428
rect 564267 492440 564313 492452
rect 564525 493428 564571 493440
rect 564525 492452 564531 493428
rect 564565 492452 564571 493428
rect 564525 492440 564571 492452
rect 564783 493428 564829 493440
rect 564783 492452 564789 493428
rect 564823 492452 564829 493428
rect 564783 492440 564829 492452
rect 565041 493428 565087 493440
rect 565041 492452 565047 493428
rect 565081 492452 565087 493428
rect 565041 492440 565087 492452
rect 565299 493428 565345 493440
rect 565299 492452 565305 493428
rect 565339 492452 565345 493428
rect 565299 492440 565345 492452
rect 565557 493428 565603 493440
rect 565557 492452 565563 493428
rect 565597 492452 565603 493428
rect 565557 492440 565603 492452
rect 565815 493428 565861 493440
rect 565815 492452 565821 493428
rect 565855 492452 565861 493428
rect 566196 492512 566404 494126
rect 575170 493624 580556 493654
rect 575170 493564 575228 493624
rect 575288 493564 575428 493624
rect 575488 493564 575628 493624
rect 575688 493564 575828 493624
rect 575888 493564 576028 493624
rect 576088 493564 576228 493624
rect 576288 493564 576428 493624
rect 576488 493564 576628 493624
rect 576688 493564 576828 493624
rect 576888 493564 577028 493624
rect 577088 493564 577228 493624
rect 577288 493564 577428 493624
rect 577488 493564 577628 493624
rect 577688 493564 577828 493624
rect 577888 493564 578028 493624
rect 578088 493564 578228 493624
rect 578288 493564 578428 493624
rect 578488 493564 578628 493624
rect 578688 493564 578828 493624
rect 578888 493564 579028 493624
rect 579088 493564 579228 493624
rect 579288 493564 579428 493624
rect 579488 493564 579628 493624
rect 579688 493564 579828 493624
rect 579888 493564 580028 493624
rect 580088 493564 580228 493624
rect 580288 493564 580556 493624
rect 575170 493534 580556 493564
rect 565815 492440 565861 492452
rect 566034 492452 566404 492512
rect 575211 493202 575257 493214
rect 560012 492324 560486 492332
rect 559792 492304 560486 492324
rect 566034 492428 566526 492452
rect 566034 492320 566074 492428
rect 566234 492320 566526 492428
rect 566034 492304 566526 492320
rect 575211 492226 575217 493202
rect 575251 492226 575257 493202
rect 575211 492214 575257 492226
rect 575469 493202 575515 493214
rect 575469 492226 575475 493202
rect 575509 492226 575515 493202
rect 575469 492214 575515 492226
rect 575727 493202 575773 493214
rect 575727 492226 575733 493202
rect 575767 492226 575773 493202
rect 575727 492214 575773 492226
rect 575985 493202 576031 493214
rect 575985 492226 575991 493202
rect 576025 492226 576031 493202
rect 575985 492214 576031 492226
rect 576243 493202 576289 493214
rect 576243 492226 576249 493202
rect 576283 492226 576289 493202
rect 576243 492214 576289 492226
rect 576501 493202 576547 493214
rect 576501 492226 576507 493202
rect 576541 492226 576547 493202
rect 576501 492214 576547 492226
rect 576759 493202 576805 493214
rect 576759 492226 576765 493202
rect 576799 492226 576805 493202
rect 576759 492214 576805 492226
rect 577017 493202 577063 493214
rect 577017 492226 577023 493202
rect 577057 492226 577063 493202
rect 577017 492214 577063 492226
rect 577275 493202 577321 493214
rect 577275 492226 577281 493202
rect 577315 492226 577321 493202
rect 577275 492214 577321 492226
rect 577533 493202 577579 493214
rect 577533 492226 577539 493202
rect 577573 492226 577579 493202
rect 577533 492214 577579 492226
rect 577791 493202 577837 493214
rect 577791 492226 577797 493202
rect 577831 492226 577837 493202
rect 577791 492214 577837 492226
rect 578049 493202 578095 493214
rect 578049 492226 578055 493202
rect 578089 492226 578095 493202
rect 578049 492214 578095 492226
rect 578307 493202 578353 493214
rect 578307 492226 578313 493202
rect 578347 492226 578353 493202
rect 578307 492214 578353 492226
rect 578565 493202 578611 493214
rect 578565 492226 578571 493202
rect 578605 492226 578611 493202
rect 578565 492214 578611 492226
rect 578823 493202 578869 493214
rect 578823 492226 578829 493202
rect 578863 492226 578869 493202
rect 578823 492214 578869 492226
rect 579081 493202 579127 493214
rect 579081 492226 579087 493202
rect 579121 492226 579127 493202
rect 579081 492214 579127 492226
rect 579339 493202 579385 493214
rect 579339 492226 579345 493202
rect 579379 492226 579385 493202
rect 579339 492214 579385 492226
rect 579597 493202 579643 493214
rect 579597 492226 579603 493202
rect 579637 492226 579643 493202
rect 579597 492214 579643 492226
rect 579855 493202 579901 493214
rect 579855 492226 579861 493202
rect 579895 492226 579901 493202
rect 579855 492214 579901 492226
rect 580113 493202 580159 493214
rect 580113 492226 580119 493202
rect 580153 492226 580159 493202
rect 580113 492214 580159 492226
rect 580371 493202 580417 493214
rect 580371 492226 580377 493202
rect 580411 492226 580417 493202
rect 580371 492214 580417 492226
rect 573506 492160 573954 492196
rect 560650 491970 565964 492000
rect 560650 491910 560836 491970
rect 560896 491910 561036 491970
rect 561096 491910 561236 491970
rect 561296 491910 561436 491970
rect 561496 491910 561636 491970
rect 561696 491910 561836 491970
rect 561896 491910 562036 491970
rect 562096 491910 562236 491970
rect 562296 491910 562436 491970
rect 562496 491910 562636 491970
rect 562696 491910 562836 491970
rect 562896 491910 563036 491970
rect 563096 491910 563236 491970
rect 563296 491910 563436 491970
rect 563496 491910 563636 491970
rect 563696 491910 563836 491970
rect 563896 491910 564036 491970
rect 564096 491910 564236 491970
rect 564296 491910 564436 491970
rect 564496 491910 564636 491970
rect 564696 491910 564836 491970
rect 564896 491910 565036 491970
rect 565096 491910 565236 491970
rect 565296 491910 565436 491970
rect 565496 491910 565636 491970
rect 565696 491910 565964 491970
rect 560650 491880 565964 491910
rect 573506 491888 573564 492160
rect 573874 492076 573954 492160
rect 580852 492130 581040 494136
rect 580530 492118 581040 492130
rect 573874 491984 575038 492076
rect 580530 492030 580542 492118
rect 580632 492030 581040 492118
rect 580530 492026 581040 492030
rect 580530 492024 580644 492026
rect 573874 491888 574934 491984
rect 573506 491880 574934 491888
rect 575026 491948 575038 491984
rect 575026 491880 575034 491948
rect 573506 491868 575034 491880
rect 575170 491744 580556 491774
rect 575170 491684 575228 491744
rect 575288 491684 575428 491744
rect 575488 491684 575628 491744
rect 575688 491684 575828 491744
rect 575888 491684 576028 491744
rect 576088 491684 576228 491744
rect 576288 491684 576428 491744
rect 576488 491684 576628 491744
rect 576688 491684 576828 491744
rect 576888 491684 577028 491744
rect 577088 491684 577228 491744
rect 577288 491684 577428 491744
rect 577488 491684 577628 491744
rect 577688 491684 577828 491744
rect 577888 491684 578028 491744
rect 578088 491684 578228 491744
rect 578288 491684 578428 491744
rect 578488 491684 578628 491744
rect 578688 491684 578828 491744
rect 578888 491684 579028 491744
rect 579088 491684 579228 491744
rect 579288 491684 579428 491744
rect 579488 491684 579628 491744
rect 579688 491684 579828 491744
rect 579888 491684 580028 491744
rect 580088 491684 580228 491744
rect 580288 491684 580556 491744
rect 575170 491654 580556 491684
rect 491168 414032 491288 414054
rect 491168 412444 491170 414032
rect 491286 412444 491288 414032
rect 491168 359028 491288 412444
rect 494928 414032 495048 414054
rect 494928 412444 494930 414032
rect 495046 412444 495048 414032
rect 493048 411584 493168 411606
rect 493048 409996 493050 411584
rect 493166 409996 493168 411584
rect 493048 408853 493168 409996
rect 493048 408819 493091 408853
rect 493125 408819 493168 408853
rect 493048 408453 493168 408819
rect 493048 408419 493091 408453
rect 493125 408419 493168 408453
rect 493048 408053 493168 408419
rect 493048 408019 493091 408053
rect 493125 408019 493168 408053
rect 493048 407653 493168 408019
rect 493048 407619 493091 407653
rect 493125 407619 493168 407653
rect 493048 407253 493168 407619
rect 493048 407219 493091 407253
rect 493125 407219 493168 407253
rect 493048 406853 493168 407219
rect 493048 406819 493091 406853
rect 493125 406819 493168 406853
rect 493048 406453 493168 406819
rect 493048 406419 493091 406453
rect 493125 406419 493168 406453
rect 493048 406053 493168 406419
rect 493048 406019 493091 406053
rect 493125 406019 493168 406053
rect 493048 405653 493168 406019
rect 493048 405619 493091 405653
rect 493125 405619 493168 405653
rect 493048 405253 493168 405619
rect 493048 405219 493091 405253
rect 493125 405219 493168 405253
rect 493048 404853 493168 405219
rect 493048 404819 493091 404853
rect 493125 404819 493168 404853
rect 493048 404453 493168 404819
rect 493048 404419 493091 404453
rect 493125 404419 493168 404453
rect 493048 404053 493168 404419
rect 493048 404019 493091 404053
rect 493125 404019 493168 404053
rect 493048 403653 493168 404019
rect 493048 403619 493091 403653
rect 493125 403619 493168 403653
rect 493048 403253 493168 403619
rect 493048 403219 493091 403253
rect 493125 403219 493168 403253
rect 493048 402853 493168 403219
rect 493048 402819 493091 402853
rect 493125 402819 493168 402853
rect 493048 402453 493168 402819
rect 493048 402419 493091 402453
rect 493125 402419 493168 402453
rect 493048 402053 493168 402419
rect 493048 402019 493091 402053
rect 493125 402019 493168 402053
rect 493048 401405 493168 402019
rect 493048 401371 493091 401405
rect 493125 401371 493168 401405
rect 493048 401005 493168 401371
rect 493048 400971 493091 401005
rect 493125 400971 493168 401005
rect 493048 400605 493168 400971
rect 493048 400571 493091 400605
rect 493125 400571 493168 400605
rect 493048 400205 493168 400571
rect 493048 400171 493091 400205
rect 493125 400171 493168 400205
rect 493048 399805 493168 400171
rect 493048 399771 493091 399805
rect 493125 399771 493168 399805
rect 493048 399405 493168 399771
rect 493048 399371 493091 399405
rect 493125 399371 493168 399405
rect 493048 399005 493168 399371
rect 493048 398971 493091 399005
rect 493125 398971 493168 399005
rect 493048 398605 493168 398971
rect 493048 398571 493091 398605
rect 493125 398571 493168 398605
rect 493048 398205 493168 398571
rect 493048 398171 493091 398205
rect 493125 398171 493168 398205
rect 493048 397805 493168 398171
rect 493048 397771 493091 397805
rect 493125 397771 493168 397805
rect 493048 397405 493168 397771
rect 493048 397371 493091 397405
rect 493125 397371 493168 397405
rect 493048 397005 493168 397371
rect 493048 396971 493091 397005
rect 493125 396971 493168 397005
rect 493048 396605 493168 396971
rect 493048 396571 493091 396605
rect 493125 396571 493168 396605
rect 493048 396205 493168 396571
rect 493048 396171 493091 396205
rect 493125 396171 493168 396205
rect 493048 395805 493168 396171
rect 493048 395771 493091 395805
rect 493125 395771 493168 395805
rect 493048 395405 493168 395771
rect 494928 408853 495048 412444
rect 498688 414032 498808 414054
rect 498688 412444 498690 414032
rect 498806 412444 498808 414032
rect 494928 408819 494971 408853
rect 495005 408819 495048 408853
rect 494928 408453 495048 408819
rect 494928 408419 494971 408453
rect 495005 408419 495048 408453
rect 494928 408053 495048 408419
rect 494928 408019 494971 408053
rect 495005 408019 495048 408053
rect 494928 407653 495048 408019
rect 494928 407619 494971 407653
rect 495005 407619 495048 407653
rect 494928 407253 495048 407619
rect 494928 407219 494971 407253
rect 495005 407219 495048 407253
rect 494928 406853 495048 407219
rect 494928 406819 494971 406853
rect 495005 406819 495048 406853
rect 494928 406453 495048 406819
rect 494928 406419 494971 406453
rect 495005 406419 495048 406453
rect 494928 406053 495048 406419
rect 494928 406019 494971 406053
rect 495005 406019 495048 406053
rect 494928 405653 495048 406019
rect 494928 405619 494971 405653
rect 495005 405619 495048 405653
rect 494928 405253 495048 405619
rect 494928 405219 494971 405253
rect 495005 405219 495048 405253
rect 494928 404853 495048 405219
rect 494928 404819 494971 404853
rect 495005 404819 495048 404853
rect 494928 404453 495048 404819
rect 494928 404419 494971 404453
rect 495005 404419 495048 404453
rect 494928 404053 495048 404419
rect 494928 404019 494971 404053
rect 495005 404019 495048 404053
rect 494928 403653 495048 404019
rect 494928 403619 494971 403653
rect 495005 403619 495048 403653
rect 494928 403253 495048 403619
rect 494928 403219 494971 403253
rect 495005 403219 495048 403253
rect 494928 402853 495048 403219
rect 494928 402819 494971 402853
rect 495005 402819 495048 402853
rect 494928 402453 495048 402819
rect 494928 402419 494971 402453
rect 495005 402419 495048 402453
rect 494928 402053 495048 402419
rect 494928 402019 494971 402053
rect 495005 402019 495048 402053
rect 494928 401405 495048 402019
rect 494928 401371 494971 401405
rect 495005 401371 495048 401405
rect 494928 401005 495048 401371
rect 494928 400971 494971 401005
rect 495005 400971 495048 401005
rect 494928 400605 495048 400971
rect 494928 400571 494971 400605
rect 495005 400571 495048 400605
rect 494928 400205 495048 400571
rect 494928 400171 494971 400205
rect 495005 400171 495048 400205
rect 494928 399805 495048 400171
rect 494928 399771 494971 399805
rect 495005 399771 495048 399805
rect 494928 399405 495048 399771
rect 494928 399371 494971 399405
rect 495005 399371 495048 399405
rect 494928 399005 495048 399371
rect 494928 398971 494971 399005
rect 495005 398971 495048 399005
rect 494928 398605 495048 398971
rect 494928 398571 494971 398605
rect 495005 398571 495048 398605
rect 494928 398205 495048 398571
rect 494928 398171 494971 398205
rect 495005 398171 495048 398205
rect 494928 397805 495048 398171
rect 494928 397771 494971 397805
rect 495005 397771 495048 397805
rect 494928 397405 495048 397771
rect 494928 397371 494971 397405
rect 495005 397371 495048 397405
rect 494928 397270 495048 397371
rect 494928 397218 494944 397270
rect 494996 397218 495048 397270
rect 494928 397005 495048 397218
rect 494928 396971 494971 397005
rect 495005 396971 495048 397005
rect 494928 396605 495048 396971
rect 494928 396571 494971 396605
rect 495005 396571 495048 396605
rect 494928 396205 495048 396571
rect 494928 396171 494971 396205
rect 495005 396171 495048 396205
rect 494928 395805 495048 396171
rect 494928 395771 494971 395805
rect 495005 395771 495048 395805
rect 494740 395522 494792 395528
rect 494740 395464 494792 395470
rect 493048 395371 493091 395405
rect 493125 395371 493168 395405
rect 493048 395005 493168 395371
rect 493048 394971 493091 395005
rect 493125 394971 493168 395005
rect 493048 394605 493168 394971
rect 493048 394571 493091 394605
rect 493125 394571 493168 394605
rect 493048 393939 493168 394571
rect 494752 394111 494780 395464
rect 494928 395405 495048 395771
rect 494928 395371 494971 395405
rect 495005 395371 495048 395405
rect 494928 395005 495048 395371
rect 494928 394971 494971 395005
rect 495005 394971 495048 395005
rect 494928 394605 495048 394971
rect 494928 394571 494971 394605
rect 495005 394571 495048 394605
rect 493048 393905 493091 393939
rect 493125 393905 493168 393939
rect 493048 393739 493168 393905
rect 493048 393705 493091 393739
rect 493125 393705 493168 393739
rect 493048 393539 493168 393705
rect 493347 394103 493909 394111
rect 493347 393709 493359 394103
rect 493897 393946 493909 394103
rect 494307 394103 494869 394111
rect 493992 393958 494044 393964
rect 493897 393918 493992 393946
rect 493897 393709 493909 393918
rect 493992 393900 494044 393906
rect 493347 393701 493909 393709
rect 494307 393709 494319 394103
rect 494857 393709 494869 394103
rect 494307 393701 494869 393709
rect 494928 393939 495048 394571
rect 494928 393905 494971 393939
rect 495005 393905 495048 393939
rect 494928 393739 495048 393905
rect 494928 393705 494971 393739
rect 495005 393705 495048 393739
rect 493048 393505 493091 393539
rect 493125 393505 493168 393539
rect 493048 393339 493168 393505
rect 493048 393305 493091 393339
rect 493125 393305 493168 393339
rect 493048 393139 493168 393305
rect 493048 393105 493091 393139
rect 493125 393105 493168 393139
rect 493048 392939 493168 393105
rect 493048 392905 493091 392939
rect 493125 392905 493168 392939
rect 493048 392739 493168 392905
rect 493048 392705 493091 392739
rect 493125 392705 493168 392739
rect 493048 392539 493168 392705
rect 493048 392505 493091 392539
rect 493125 392505 493168 392539
rect 493048 392339 493168 392505
rect 493048 392305 493091 392339
rect 493125 392305 493168 392339
rect 493048 392139 493168 392305
rect 493048 392105 493091 392139
rect 493125 392105 493168 392139
rect 494928 393539 495048 393705
rect 494928 393505 494971 393539
rect 495005 393505 495048 393539
rect 494928 393339 495048 393505
rect 494928 393305 494971 393339
rect 495005 393305 495048 393339
rect 494928 393139 495048 393305
rect 494928 393105 494971 393139
rect 495005 393105 495048 393139
rect 494928 392939 495048 393105
rect 494928 392905 494971 392939
rect 495005 392905 495048 392939
rect 494928 392739 495048 392905
rect 494928 392705 494971 392739
rect 495005 392705 495048 392739
rect 494928 392539 495048 392705
rect 494928 392505 494971 392539
rect 495005 392505 495048 392539
rect 494928 392339 495048 392505
rect 494928 392305 494971 392339
rect 495005 392305 495048 392339
rect 494928 392139 495048 392305
rect 493048 391939 493168 392105
rect 493909 392103 494873 392114
rect 493048 391905 493091 391939
rect 493125 391905 493168 391939
rect 493048 390853 493168 391905
rect 493347 392096 494873 392103
rect 493347 391702 493359 392096
rect 493897 391702 494319 392096
rect 494857 391702 494873 392096
rect 493347 391693 494873 391702
rect 493909 391682 494873 391693
rect 494928 392105 494971 392139
rect 495005 392105 495048 392139
rect 494928 391939 495048 392105
rect 494928 391905 494971 391939
rect 495005 391905 495048 391939
rect 494808 391198 494860 391204
rect 494808 391140 494860 391146
rect 493588 391024 494388 391030
rect 493588 390990 493611 391024
rect 493645 390990 493683 391024
rect 493717 390990 493755 391024
rect 493789 390990 493827 391024
rect 493861 390990 493899 391024
rect 493933 390990 493971 391024
rect 494005 390990 494043 391024
rect 494077 390990 494115 391024
rect 494149 390990 494187 391024
rect 494221 390990 494259 391024
rect 494293 390990 494331 391024
rect 494365 390990 494388 391024
rect 493588 390984 494388 390990
rect 494344 390910 494372 390984
rect 494820 390925 494848 391140
rect 494811 390913 494857 390925
rect 494811 390910 494817 390913
rect 494344 390882 494817 390910
rect 494811 390879 494817 390882
rect 494851 390879 494857 390913
rect 494811 390867 494857 390879
rect 493048 390819 493091 390853
rect 493125 390819 493168 390853
rect 493048 389941 493168 390819
rect 494928 390853 495048 391905
rect 494928 390819 494971 390853
rect 495005 390819 495048 390853
rect 494928 390634 495048 390819
rect 494344 390606 495048 390634
rect 494344 390572 494372 390606
rect 493588 390566 494388 390572
rect 493588 390532 493611 390566
rect 493645 390532 493683 390566
rect 493717 390532 493755 390566
rect 493789 390532 493827 390566
rect 493861 390532 493899 390566
rect 493933 390532 493971 390566
rect 494005 390532 494043 390566
rect 494077 390532 494115 390566
rect 494149 390532 494187 390566
rect 494221 390532 494259 390566
rect 494293 390532 494331 390566
rect 494365 390532 494388 390566
rect 493588 390526 494388 390532
rect 493343 390077 494633 390083
rect 493343 390043 493359 390077
rect 493393 390043 493431 390077
rect 493465 390043 493503 390077
rect 493537 390043 493575 390077
rect 493609 390043 493647 390077
rect 493681 390043 493719 390077
rect 493753 390043 493791 390077
rect 493825 390043 493863 390077
rect 493897 390043 493935 390077
rect 493969 390043 494007 390077
rect 494041 390043 494079 390077
rect 494113 390043 494151 390077
rect 494185 390043 494223 390077
rect 494257 390043 494295 390077
rect 494329 390043 494367 390077
rect 494401 390043 494439 390077
rect 494473 390043 494511 390077
rect 494545 390043 494583 390077
rect 494617 390043 494633 390077
rect 493343 390037 494633 390043
rect 493048 389907 493091 389941
rect 493125 389907 493168 389941
rect 493048 389622 493168 389907
rect 494928 389941 495048 390606
rect 494928 389907 494971 389941
rect 495005 389907 495048 389941
rect 493343 389622 494633 389625
rect 493048 389619 494633 389622
rect 493048 389594 493359 389619
rect 493048 389541 493168 389594
rect 493343 389585 493359 389594
rect 493393 389585 493431 389619
rect 493465 389585 493503 389619
rect 493537 389585 493575 389619
rect 493609 389585 493647 389619
rect 493681 389585 493719 389619
rect 493753 389585 493791 389619
rect 493825 389585 493863 389619
rect 493897 389585 493935 389619
rect 493969 389585 494007 389619
rect 494041 389585 494079 389619
rect 494113 389585 494151 389619
rect 494185 389585 494223 389619
rect 494257 389585 494295 389619
rect 494329 389585 494367 389619
rect 494401 389585 494439 389619
rect 494473 389585 494511 389619
rect 494545 389585 494583 389619
rect 494617 389585 494633 389619
rect 493343 389579 494633 389585
rect 493048 389507 493091 389541
rect 493125 389507 493168 389541
rect 493048 389141 493168 389507
rect 494928 389541 495048 389907
rect 494928 389507 494971 389541
rect 495005 389507 495048 389541
rect 493048 389107 493091 389141
rect 493125 389107 493168 389141
rect 493343 389161 494633 389167
rect 493343 389127 493359 389161
rect 493393 389127 493431 389161
rect 493465 389127 493503 389161
rect 493537 389127 493575 389161
rect 493609 389127 493647 389161
rect 493681 389127 493719 389161
rect 493753 389127 493791 389161
rect 493825 389127 493863 389161
rect 493897 389127 493935 389161
rect 493969 389127 494007 389161
rect 494041 389127 494079 389161
rect 494113 389127 494151 389161
rect 494185 389127 494223 389161
rect 494257 389127 494295 389161
rect 494329 389127 494367 389161
rect 494401 389127 494439 389161
rect 494473 389127 494511 389161
rect 494545 389127 494583 389161
rect 494617 389127 494633 389161
rect 493343 389121 494633 389127
rect 494928 389141 495048 389507
rect 493048 388741 493168 389107
rect 493048 388707 493091 388741
rect 493125 388707 493168 388741
rect 494928 389107 494971 389141
rect 495005 389107 495048 389141
rect 494928 388741 495048 389107
rect 493048 388341 493168 388707
rect 493343 388703 494633 388709
rect 493343 388669 493359 388703
rect 493393 388669 493431 388703
rect 493465 388669 493503 388703
rect 493537 388669 493575 388703
rect 493609 388669 493647 388703
rect 493681 388669 493719 388703
rect 493753 388669 493791 388703
rect 493825 388669 493863 388703
rect 493897 388669 493935 388703
rect 493969 388669 494007 388703
rect 494041 388669 494079 388703
rect 494113 388669 494151 388703
rect 494185 388669 494223 388703
rect 494257 388669 494295 388703
rect 494329 388669 494367 388703
rect 494401 388669 494439 388703
rect 494473 388669 494511 388703
rect 494545 388669 494583 388703
rect 494617 388669 494633 388703
rect 493343 388663 494633 388669
rect 494928 388707 494971 388741
rect 495005 388707 495048 388741
rect 493048 388307 493091 388341
rect 493125 388307 493168 388341
rect 493048 387941 493168 388307
rect 494928 388341 495048 388707
rect 494928 388307 494971 388341
rect 495005 388307 495048 388341
rect 493343 388245 494633 388251
rect 493343 388211 493359 388245
rect 493393 388211 493431 388245
rect 493465 388211 493503 388245
rect 493537 388211 493575 388245
rect 493609 388211 493647 388245
rect 493681 388211 493719 388245
rect 493753 388211 493791 388245
rect 493825 388211 493863 388245
rect 493897 388211 493935 388245
rect 493969 388211 494007 388245
rect 494041 388211 494079 388245
rect 494113 388211 494151 388245
rect 494185 388211 494223 388245
rect 494257 388211 494295 388245
rect 494329 388211 494367 388245
rect 494401 388211 494439 388245
rect 494473 388211 494511 388245
rect 494545 388211 494583 388245
rect 494617 388211 494633 388245
rect 493343 388205 494633 388211
rect 493048 387907 493091 387941
rect 493125 387907 493168 387941
rect 493048 387541 493168 387907
rect 494928 387941 495048 388307
rect 494928 387907 494971 387941
rect 495005 387907 495048 387941
rect 493343 387787 494633 387793
rect 493343 387753 493359 387787
rect 493393 387753 493431 387787
rect 493465 387753 493503 387787
rect 493537 387753 493575 387787
rect 493609 387753 493647 387787
rect 493681 387753 493719 387787
rect 493753 387753 493791 387787
rect 493825 387753 493863 387787
rect 493897 387753 493935 387787
rect 493969 387753 494007 387787
rect 494041 387753 494079 387787
rect 494113 387753 494151 387787
rect 494185 387753 494223 387787
rect 494257 387753 494295 387787
rect 494329 387753 494367 387787
rect 494401 387753 494439 387787
rect 494473 387753 494511 387787
rect 494545 387753 494583 387787
rect 494617 387753 494633 387787
rect 493343 387747 494633 387753
rect 493048 387507 493091 387541
rect 493125 387507 493168 387541
rect 493048 387141 493168 387507
rect 494928 387541 495048 387907
rect 494928 387507 494971 387541
rect 495005 387507 495048 387541
rect 493343 387329 494633 387335
rect 493343 387295 493359 387329
rect 493393 387295 493431 387329
rect 493465 387295 493503 387329
rect 493537 387295 493575 387329
rect 493609 387295 493647 387329
rect 493681 387295 493719 387329
rect 493753 387295 493791 387329
rect 493825 387295 493863 387329
rect 493897 387295 493935 387329
rect 493969 387295 494007 387329
rect 494041 387295 494079 387329
rect 494113 387295 494151 387329
rect 494185 387295 494223 387329
rect 494257 387295 494295 387329
rect 494329 387295 494367 387329
rect 494401 387295 494439 387329
rect 494473 387295 494511 387329
rect 494545 387295 494583 387329
rect 494617 387295 494633 387329
rect 493343 387289 494633 387295
rect 493048 387107 493091 387141
rect 493125 387107 493168 387141
rect 493048 386741 493168 387107
rect 494928 387141 495048 387507
rect 494928 387107 494971 387141
rect 495005 387107 495048 387141
rect 493343 386871 494633 386877
rect 493343 386837 493359 386871
rect 493393 386837 493431 386871
rect 493465 386837 493503 386871
rect 493537 386837 493575 386871
rect 493609 386837 493647 386871
rect 493681 386837 493719 386871
rect 493753 386837 493791 386871
rect 493825 386837 493863 386871
rect 493897 386837 493935 386871
rect 493969 386837 494007 386871
rect 494041 386837 494079 386871
rect 494113 386837 494151 386871
rect 494185 386837 494223 386871
rect 494257 386837 494295 386871
rect 494329 386837 494367 386871
rect 494401 386837 494439 386871
rect 494473 386837 494511 386871
rect 494545 386837 494583 386871
rect 494617 386837 494633 386871
rect 493343 386831 494633 386837
rect 493048 386707 493091 386741
rect 493125 386707 493168 386741
rect 493048 386341 493168 386707
rect 494928 386741 495048 387107
rect 494928 386707 494971 386741
rect 495005 386707 495048 386741
rect 493343 386413 494633 386419
rect 493343 386379 493359 386413
rect 493393 386379 493431 386413
rect 493465 386379 493503 386413
rect 493537 386379 493575 386413
rect 493609 386379 493647 386413
rect 493681 386379 493719 386413
rect 493753 386379 493791 386413
rect 493825 386379 493863 386413
rect 493897 386379 493935 386413
rect 493969 386379 494007 386413
rect 494041 386379 494079 386413
rect 494113 386379 494151 386413
rect 494185 386379 494223 386413
rect 494257 386379 494295 386413
rect 494329 386379 494367 386413
rect 494401 386379 494439 386413
rect 494473 386379 494511 386413
rect 494545 386379 494583 386413
rect 494617 386379 494633 386413
rect 493343 386373 494633 386379
rect 493048 386307 493091 386341
rect 493125 386307 493168 386341
rect 493048 385941 493168 386307
rect 494928 386341 495048 386707
rect 494928 386307 494971 386341
rect 495005 386307 495048 386341
rect 493048 385907 493091 385941
rect 493125 385907 493168 385941
rect 493343 385955 494633 385961
rect 493343 385921 493359 385955
rect 493393 385921 493431 385955
rect 493465 385921 493503 385955
rect 493537 385921 493575 385955
rect 493609 385921 493647 385955
rect 493681 385921 493719 385955
rect 493753 385921 493791 385955
rect 493825 385921 493863 385955
rect 493897 385921 493935 385955
rect 493969 385921 494007 385955
rect 494041 385921 494079 385955
rect 494113 385921 494151 385955
rect 494185 385921 494223 385955
rect 494257 385921 494295 385955
rect 494329 385921 494367 385955
rect 494401 385921 494439 385955
rect 494473 385921 494511 385955
rect 494545 385921 494583 385955
rect 494617 385921 494633 385955
rect 493343 385915 494633 385921
rect 494928 385941 495048 386307
rect 493048 385541 493168 385907
rect 494928 385907 494971 385941
rect 495005 385907 495048 385941
rect 493048 385507 493091 385541
rect 493125 385507 493168 385541
rect 493048 385141 493168 385507
rect 493343 385497 494633 385503
rect 494820 385500 494848 385555
rect 494928 385541 495048 385907
rect 494928 385507 494971 385541
rect 495005 385507 495048 385541
rect 493343 385463 493359 385497
rect 493393 385463 493431 385497
rect 493465 385463 493503 385497
rect 493537 385463 493575 385497
rect 493609 385463 493647 385497
rect 493681 385463 493719 385497
rect 493753 385463 493791 385497
rect 493825 385463 493863 385497
rect 493897 385463 493935 385497
rect 493969 385463 494007 385497
rect 494041 385463 494079 385497
rect 494113 385463 494151 385497
rect 494185 385463 494223 385497
rect 494257 385463 494295 385497
rect 494329 385463 494367 385497
rect 494401 385463 494439 385497
rect 494473 385463 494511 385497
rect 494545 385463 494583 385497
rect 494617 385463 494633 385497
rect 493343 385457 494633 385463
rect 494808 385494 494860 385500
rect 494808 385436 494860 385442
rect 493048 385107 493091 385141
rect 493125 385107 493168 385141
rect 493048 384741 493168 385107
rect 494928 385141 495048 385507
rect 494928 385107 494971 385141
rect 495005 385107 495048 385141
rect 493343 385039 494633 385045
rect 493343 385005 493359 385039
rect 493393 385005 493431 385039
rect 493465 385005 493503 385039
rect 493537 385005 493575 385039
rect 493609 385005 493647 385039
rect 493681 385005 493719 385039
rect 493753 385005 493791 385039
rect 493825 385005 493863 385039
rect 493897 385005 493935 385039
rect 493969 385005 494007 385039
rect 494041 385005 494079 385039
rect 494113 385005 494151 385039
rect 494185 385005 494223 385039
rect 494257 385005 494295 385039
rect 494329 385005 494367 385039
rect 494401 385005 494439 385039
rect 494473 385005 494511 385039
rect 494545 385005 494583 385039
rect 494617 385005 494633 385039
rect 493343 384999 494633 385005
rect 493048 384707 493091 384741
rect 493125 384707 493168 384741
rect 493048 384341 493168 384707
rect 494928 384741 495048 385107
rect 494928 384707 494971 384741
rect 495005 384707 495048 384741
rect 493343 384581 494633 384587
rect 493343 384547 493359 384581
rect 493393 384547 493431 384581
rect 493465 384547 493503 384581
rect 493537 384547 493575 384581
rect 493609 384547 493647 384581
rect 493681 384547 493719 384581
rect 493753 384547 493791 384581
rect 493825 384547 493863 384581
rect 493897 384547 493935 384581
rect 493969 384547 494007 384581
rect 494041 384547 494079 384581
rect 494113 384547 494151 384581
rect 494185 384547 494223 384581
rect 494257 384547 494295 384581
rect 494329 384547 494367 384581
rect 494401 384547 494439 384581
rect 494473 384547 494511 384581
rect 494545 384547 494583 384581
rect 494617 384547 494633 384581
rect 493343 384541 494633 384547
rect 493048 384307 493091 384341
rect 493125 384307 493168 384341
rect 493048 383941 493168 384307
rect 494928 384341 495048 384707
rect 494928 384307 494971 384341
rect 495005 384307 495048 384341
rect 493343 384123 494633 384129
rect 493343 384089 493359 384123
rect 493393 384089 493431 384123
rect 493465 384089 493503 384123
rect 493537 384089 493575 384123
rect 493609 384089 493647 384123
rect 493681 384089 493719 384123
rect 493753 384089 493791 384123
rect 493825 384089 493863 384123
rect 493897 384089 493935 384123
rect 493969 384089 494007 384123
rect 494041 384089 494079 384123
rect 494113 384089 494151 384123
rect 494185 384089 494223 384123
rect 494257 384089 494295 384123
rect 494329 384089 494367 384123
rect 494401 384089 494439 384123
rect 494473 384089 494511 384123
rect 494545 384089 494583 384123
rect 494617 384089 494633 384123
rect 493343 384083 494633 384089
rect 493048 383907 493091 383941
rect 493125 383907 493168 383941
rect 493048 383541 493168 383907
rect 494928 383941 495048 384307
rect 494928 383907 494971 383941
rect 495005 383907 495048 383941
rect 493343 383665 494633 383671
rect 493343 383631 493359 383665
rect 493393 383631 493431 383665
rect 493465 383631 493503 383665
rect 493537 383631 493575 383665
rect 493609 383631 493647 383665
rect 493681 383631 493719 383665
rect 493753 383631 493791 383665
rect 493825 383631 493863 383665
rect 493897 383631 493935 383665
rect 493969 383631 494007 383665
rect 494041 383631 494079 383665
rect 494113 383631 494151 383665
rect 494185 383631 494223 383665
rect 494257 383631 494295 383665
rect 494329 383631 494367 383665
rect 494401 383631 494439 383665
rect 494473 383631 494511 383665
rect 494545 383631 494583 383665
rect 494617 383631 494633 383665
rect 493343 383625 494633 383631
rect 493048 383507 493091 383541
rect 493125 383507 493168 383541
rect 493048 383141 493168 383507
rect 494928 383541 495048 383907
rect 494928 383507 494971 383541
rect 495005 383507 495048 383541
rect 493343 383207 494633 383213
rect 493343 383173 493359 383207
rect 493393 383173 493431 383207
rect 493465 383173 493503 383207
rect 493537 383173 493575 383207
rect 493609 383173 493647 383207
rect 493681 383173 493719 383207
rect 493753 383173 493791 383207
rect 493825 383173 493863 383207
rect 493897 383173 493935 383207
rect 493969 383173 494007 383207
rect 494041 383173 494079 383207
rect 494113 383173 494151 383207
rect 494185 383173 494223 383207
rect 494257 383173 494295 383207
rect 494329 383173 494367 383207
rect 494401 383173 494439 383207
rect 494473 383173 494511 383207
rect 494545 383173 494583 383207
rect 494617 383173 494633 383207
rect 493343 383167 494633 383173
rect 493048 383107 493091 383141
rect 493125 383107 493168 383141
rect 493048 382741 493168 383107
rect 494928 383141 495048 383507
rect 494928 383107 494971 383141
rect 495005 383107 495048 383141
rect 493048 382707 493091 382741
rect 493125 382707 493168 382741
rect 493343 382749 494633 382755
rect 493343 382715 493359 382749
rect 493393 382715 493431 382749
rect 493465 382715 493503 382749
rect 493537 382715 493575 382749
rect 493609 382715 493647 382749
rect 493681 382715 493719 382749
rect 493753 382715 493791 382749
rect 493825 382715 493863 382749
rect 493897 382715 493935 382749
rect 493969 382715 494007 382749
rect 494041 382715 494079 382749
rect 494113 382715 494151 382749
rect 494185 382715 494223 382749
rect 494257 382715 494295 382749
rect 494329 382715 494367 382749
rect 494401 382715 494439 382749
rect 494473 382715 494511 382749
rect 494545 382715 494583 382749
rect 494617 382715 494633 382749
rect 493343 382709 494633 382715
rect 494928 382741 495048 383107
rect 493048 382341 493168 382707
rect 493048 382307 493091 382341
rect 493125 382307 493168 382341
rect 493048 381941 493168 382307
rect 494928 382707 494971 382741
rect 495005 382707 495048 382741
rect 494928 382341 495048 382707
rect 494928 382307 494971 382341
rect 495005 382307 495048 382341
rect 493343 382291 494633 382297
rect 493343 382257 493359 382291
rect 493393 382257 493431 382291
rect 493465 382257 493503 382291
rect 493537 382257 493575 382291
rect 493609 382257 493647 382291
rect 493681 382257 493719 382291
rect 493753 382257 493791 382291
rect 493825 382257 493863 382291
rect 493897 382257 493935 382291
rect 493969 382257 494007 382291
rect 494041 382257 494079 382291
rect 494113 382257 494151 382291
rect 494185 382257 494223 382291
rect 494257 382257 494295 382291
rect 494329 382257 494367 382291
rect 494401 382257 494439 382291
rect 494473 382257 494511 382291
rect 494545 382257 494583 382291
rect 494617 382257 494633 382291
rect 493343 382251 494633 382257
rect 493048 381907 493091 381941
rect 493125 381907 493168 381941
rect 493048 381541 493168 381907
rect 494928 381941 495048 382307
rect 494928 381907 494971 381941
rect 495005 381907 495048 381941
rect 493343 381833 494633 381839
rect 493343 381799 493359 381833
rect 493393 381799 493431 381833
rect 493465 381799 493503 381833
rect 493537 381799 493575 381833
rect 493609 381799 493647 381833
rect 493681 381799 493719 381833
rect 493753 381799 493791 381833
rect 493825 381799 493863 381833
rect 493897 381799 493935 381833
rect 493969 381799 494007 381833
rect 494041 381799 494079 381833
rect 494113 381799 494151 381833
rect 494185 381799 494223 381833
rect 494257 381799 494295 381833
rect 494329 381799 494367 381833
rect 494401 381799 494439 381833
rect 494473 381799 494511 381833
rect 494545 381799 494583 381833
rect 494617 381799 494633 381833
rect 493343 381793 494633 381799
rect 493048 381507 493091 381541
rect 493125 381507 493168 381541
rect 493048 381141 493168 381507
rect 494928 381541 495048 381907
rect 494928 381507 494971 381541
rect 495005 381507 495048 381541
rect 493343 381375 494633 381381
rect 493343 381341 493359 381375
rect 493393 381341 493431 381375
rect 493465 381341 493503 381375
rect 493537 381341 493575 381375
rect 493609 381341 493647 381375
rect 493681 381341 493719 381375
rect 493753 381341 493791 381375
rect 493825 381341 493863 381375
rect 493897 381341 493935 381375
rect 493969 381341 494007 381375
rect 494041 381341 494079 381375
rect 494113 381341 494151 381375
rect 494185 381341 494223 381375
rect 494257 381341 494295 381375
rect 494329 381341 494367 381375
rect 494401 381341 494439 381375
rect 494473 381341 494511 381375
rect 494545 381341 494583 381375
rect 494617 381341 494633 381375
rect 493343 381335 494633 381341
rect 493048 381107 493091 381141
rect 493125 381107 493168 381141
rect 493048 380741 493168 381107
rect 494928 381141 495048 381507
rect 494928 381107 494971 381141
rect 495005 381107 495048 381141
rect 493343 380917 494633 380923
rect 493343 380883 493359 380917
rect 493393 380883 493431 380917
rect 493465 380883 493503 380917
rect 493537 380883 493575 380917
rect 493609 380883 493647 380917
rect 493681 380883 493719 380917
rect 493753 380883 493791 380917
rect 493825 380883 493863 380917
rect 493897 380883 493935 380917
rect 493969 380883 494007 380917
rect 494041 380883 494079 380917
rect 494113 380883 494151 380917
rect 494185 380883 494223 380917
rect 494257 380883 494295 380917
rect 494329 380883 494367 380917
rect 494401 380883 494439 380917
rect 494473 380883 494511 380917
rect 494545 380883 494583 380917
rect 494617 380883 494633 380917
rect 493343 380877 494633 380883
rect 493048 380707 493091 380741
rect 493125 380707 493168 380741
rect 493048 380341 493168 380707
rect 494928 380741 495048 381107
rect 494928 380707 494971 380741
rect 495005 380707 495048 380741
rect 493343 380459 494633 380465
rect 493343 380425 493359 380459
rect 493393 380425 493431 380459
rect 493465 380425 493503 380459
rect 493537 380425 493575 380459
rect 493609 380425 493647 380459
rect 493681 380425 493719 380459
rect 493753 380425 493791 380459
rect 493825 380425 493863 380459
rect 493897 380425 493935 380459
rect 493969 380425 494007 380459
rect 494041 380425 494079 380459
rect 494113 380425 494151 380459
rect 494185 380425 494223 380459
rect 494257 380425 494295 380459
rect 494329 380425 494367 380459
rect 494401 380425 494439 380459
rect 494473 380425 494511 380459
rect 494545 380425 494583 380459
rect 494617 380425 494633 380459
rect 493343 380419 494633 380425
rect 493048 380307 493091 380341
rect 493125 380307 493168 380341
rect 493048 379941 493168 380307
rect 494928 380341 495048 380707
rect 494928 380307 494971 380341
rect 495005 380307 495048 380341
rect 493343 380001 494633 380007
rect 493343 379967 493359 380001
rect 493393 379967 493431 380001
rect 493465 379967 493503 380001
rect 493537 379967 493575 380001
rect 493609 379967 493647 380001
rect 493681 379967 493719 380001
rect 493753 379967 493791 380001
rect 493825 379967 493863 380001
rect 493897 379967 493935 380001
rect 493969 379967 494007 380001
rect 494041 379967 494079 380001
rect 494113 379967 494151 380001
rect 494185 379967 494223 380001
rect 494257 379967 494295 380001
rect 494329 379967 494367 380001
rect 494401 379967 494439 380001
rect 494473 379967 494511 380001
rect 494545 379967 494583 380001
rect 494617 379967 494633 380001
rect 493343 379961 494633 379967
rect 493048 379907 493091 379941
rect 493125 379907 493168 379941
rect 493048 379541 493168 379907
rect 494928 379941 495048 380307
rect 494928 379907 494971 379941
rect 495005 379907 495048 379941
rect 493048 379507 493091 379541
rect 493125 379507 493168 379541
rect 493048 379141 493168 379507
rect 493343 379543 494633 379549
rect 493343 379509 493359 379543
rect 493393 379509 493431 379543
rect 493465 379509 493503 379543
rect 493537 379509 493575 379543
rect 493609 379509 493647 379543
rect 493681 379509 493719 379543
rect 493753 379509 493791 379543
rect 493825 379509 493863 379543
rect 493897 379509 493935 379543
rect 493969 379509 494007 379543
rect 494041 379509 494079 379543
rect 494113 379509 494151 379543
rect 494185 379509 494223 379543
rect 494257 379509 494295 379543
rect 494329 379509 494367 379543
rect 494401 379509 494439 379543
rect 494473 379509 494511 379543
rect 494545 379509 494583 379543
rect 494617 379509 494633 379543
rect 493343 379503 494633 379509
rect 494928 379541 495048 379907
rect 494928 379507 494971 379541
rect 495005 379507 495048 379541
rect 493048 379107 493091 379141
rect 493125 379107 493168 379141
rect 493048 378741 493168 379107
rect 494928 379141 495048 379507
rect 494928 379107 494971 379141
rect 495005 379107 495048 379141
rect 493343 379085 494633 379091
rect 493343 379051 493359 379085
rect 493393 379051 493431 379085
rect 493465 379051 493503 379085
rect 493537 379051 493575 379085
rect 493609 379051 493647 379085
rect 493681 379051 493719 379085
rect 493753 379051 493791 379085
rect 493825 379051 493863 379085
rect 493897 379051 493935 379085
rect 493969 379051 494007 379085
rect 494041 379051 494079 379085
rect 494113 379051 494151 379085
rect 494185 379051 494223 379085
rect 494257 379051 494295 379085
rect 494329 379051 494367 379085
rect 494401 379051 494439 379085
rect 494473 379051 494511 379085
rect 494545 379051 494583 379085
rect 494617 379051 494633 379085
rect 493343 379045 494633 379051
rect 493048 378707 493091 378741
rect 493125 378707 493168 378741
rect 493048 378341 493168 378707
rect 494928 378741 495048 379107
rect 494928 378707 494971 378741
rect 495005 378707 495048 378741
rect 493343 378627 494633 378633
rect 493343 378593 493359 378627
rect 493393 378593 493431 378627
rect 493465 378593 493503 378627
rect 493537 378593 493575 378627
rect 493609 378593 493647 378627
rect 493681 378593 493719 378627
rect 493753 378593 493791 378627
rect 493825 378593 493863 378627
rect 493897 378593 493935 378627
rect 493969 378593 494007 378627
rect 494041 378593 494079 378627
rect 494113 378593 494151 378627
rect 494185 378593 494223 378627
rect 494257 378593 494295 378627
rect 494329 378593 494367 378627
rect 494401 378593 494439 378627
rect 494473 378593 494511 378627
rect 494545 378593 494583 378627
rect 494617 378593 494633 378627
rect 493343 378587 494633 378593
rect 493048 378307 493091 378341
rect 493125 378307 493168 378341
rect 493048 377941 493168 378307
rect 494928 378341 495048 378707
rect 494928 378307 494971 378341
rect 495005 378307 495048 378341
rect 493343 378169 494633 378175
rect 493343 378135 493359 378169
rect 493393 378135 493431 378169
rect 493465 378135 493503 378169
rect 493537 378135 493575 378169
rect 493609 378135 493647 378169
rect 493681 378135 493719 378169
rect 493753 378135 493791 378169
rect 493825 378135 493863 378169
rect 493897 378135 493935 378169
rect 493969 378135 494007 378169
rect 494041 378135 494079 378169
rect 494113 378135 494151 378169
rect 494185 378135 494223 378169
rect 494257 378135 494295 378169
rect 494329 378135 494367 378169
rect 494401 378135 494439 378169
rect 494473 378135 494511 378169
rect 494545 378135 494583 378169
rect 494617 378135 494633 378169
rect 493343 378129 494633 378135
rect 493048 377907 493091 377941
rect 493125 377907 493168 377941
rect 493048 377541 493168 377907
rect 494928 377941 495048 378307
rect 494928 377907 494971 377941
rect 495005 377907 495048 377941
rect 493343 377711 494633 377717
rect 493343 377677 493359 377711
rect 493393 377677 493431 377711
rect 493465 377677 493503 377711
rect 493537 377677 493575 377711
rect 493609 377677 493647 377711
rect 493681 377677 493719 377711
rect 493753 377677 493791 377711
rect 493825 377677 493863 377711
rect 493897 377677 493935 377711
rect 493969 377677 494007 377711
rect 494041 377677 494079 377711
rect 494113 377677 494151 377711
rect 494185 377677 494223 377711
rect 494257 377677 494295 377711
rect 494329 377677 494367 377711
rect 494401 377677 494439 377711
rect 494473 377677 494511 377711
rect 494545 377677 494583 377711
rect 494617 377677 494633 377711
rect 493343 377671 494633 377677
rect 493048 377507 493091 377541
rect 493125 377507 493168 377541
rect 493048 377141 493168 377507
rect 494928 377541 495048 377907
rect 494928 377507 494971 377541
rect 495005 377507 495048 377541
rect 493343 377253 494633 377259
rect 493343 377219 493359 377253
rect 493393 377219 493431 377253
rect 493465 377219 493503 377253
rect 493537 377219 493575 377253
rect 493609 377219 493647 377253
rect 493681 377219 493719 377253
rect 493753 377219 493791 377253
rect 493825 377219 493863 377253
rect 493897 377219 493935 377253
rect 493969 377219 494007 377253
rect 494041 377219 494079 377253
rect 494113 377219 494151 377253
rect 494185 377219 494223 377253
rect 494257 377219 494295 377253
rect 494329 377219 494367 377253
rect 494401 377219 494439 377253
rect 494473 377219 494511 377253
rect 494545 377219 494583 377253
rect 494617 377219 494633 377253
rect 493343 377213 494633 377219
rect 493048 377107 493091 377141
rect 493125 377107 493168 377141
rect 493048 376741 493168 377107
rect 494928 377141 495048 377507
rect 494928 377107 494971 377141
rect 495005 377107 495048 377141
rect 493343 376795 494633 376801
rect 493343 376761 493359 376795
rect 493393 376761 493431 376795
rect 493465 376761 493503 376795
rect 493537 376761 493575 376795
rect 493609 376761 493647 376795
rect 493681 376761 493719 376795
rect 493753 376761 493791 376795
rect 493825 376761 493863 376795
rect 493897 376761 493935 376795
rect 493969 376761 494007 376795
rect 494041 376761 494079 376795
rect 494113 376761 494151 376795
rect 494185 376761 494223 376795
rect 494257 376761 494295 376795
rect 494329 376761 494367 376795
rect 494401 376761 494439 376795
rect 494473 376761 494511 376795
rect 494545 376761 494583 376795
rect 494617 376761 494633 376795
rect 493343 376755 494633 376761
rect 493048 376707 493091 376741
rect 493125 376707 493168 376741
rect 493048 376341 493168 376707
rect 494928 376741 495048 377107
rect 494928 376707 494971 376741
rect 495005 376707 495048 376741
rect 493048 376307 493091 376341
rect 493125 376307 493168 376341
rect 493048 375941 493168 376307
rect 493343 376337 494633 376343
rect 493343 376303 493359 376337
rect 493393 376303 493431 376337
rect 493465 376303 493503 376337
rect 493537 376303 493575 376337
rect 493609 376303 493647 376337
rect 493681 376303 493719 376337
rect 493753 376303 493791 376337
rect 493825 376303 493863 376337
rect 493897 376303 493935 376337
rect 493969 376303 494007 376337
rect 494041 376303 494079 376337
rect 494113 376303 494151 376337
rect 494185 376303 494223 376337
rect 494257 376303 494295 376337
rect 494329 376303 494367 376337
rect 494401 376303 494439 376337
rect 494473 376303 494511 376337
rect 494545 376303 494583 376337
rect 494617 376303 494633 376337
rect 493343 376297 494633 376303
rect 494928 376341 495048 376707
rect 494928 376307 494971 376341
rect 495005 376307 495048 376341
rect 493048 375907 493091 375941
rect 493125 375907 493168 375941
rect 493048 375541 493168 375907
rect 494928 375941 495048 376307
rect 494928 375907 494971 375941
rect 495005 375907 495048 375941
rect 493343 375879 494633 375885
rect 493343 375845 493359 375879
rect 493393 375845 493431 375879
rect 493465 375845 493503 375879
rect 493537 375845 493575 375879
rect 493609 375845 493647 375879
rect 493681 375845 493719 375879
rect 493753 375845 493791 375879
rect 493825 375845 493863 375879
rect 493897 375845 493935 375879
rect 493969 375845 494007 375879
rect 494041 375845 494079 375879
rect 494113 375845 494151 375879
rect 494185 375845 494223 375879
rect 494257 375845 494295 375879
rect 494329 375845 494367 375879
rect 494401 375845 494439 375879
rect 494473 375845 494511 375879
rect 494545 375845 494583 375879
rect 494617 375845 494633 375879
rect 493343 375839 494633 375845
rect 493048 375507 493091 375541
rect 493125 375507 493168 375541
rect 493048 375141 493168 375507
rect 494928 375541 495048 375907
rect 494928 375507 494971 375541
rect 495005 375507 495048 375541
rect 493343 375421 494633 375427
rect 493343 375387 493359 375421
rect 493393 375387 493431 375421
rect 493465 375387 493503 375421
rect 493537 375387 493575 375421
rect 493609 375387 493647 375421
rect 493681 375387 493719 375421
rect 493753 375387 493791 375421
rect 493825 375387 493863 375421
rect 493897 375387 493935 375421
rect 493969 375387 494007 375421
rect 494041 375387 494079 375421
rect 494113 375387 494151 375421
rect 494185 375387 494223 375421
rect 494257 375387 494295 375421
rect 494329 375387 494367 375421
rect 494401 375387 494439 375421
rect 494473 375387 494511 375421
rect 494545 375387 494583 375421
rect 494617 375387 494633 375421
rect 493343 375381 494633 375387
rect 493048 375107 493091 375141
rect 493125 375107 493168 375141
rect 493048 374741 493168 375107
rect 494928 375141 495048 375507
rect 494928 375107 494971 375141
rect 495005 375107 495048 375141
rect 493343 374963 494633 374969
rect 493343 374929 493359 374963
rect 493393 374929 493431 374963
rect 493465 374929 493503 374963
rect 493537 374929 493575 374963
rect 493609 374929 493647 374963
rect 493681 374929 493719 374963
rect 493753 374929 493791 374963
rect 493825 374929 493863 374963
rect 493897 374929 493935 374963
rect 493969 374929 494007 374963
rect 494041 374929 494079 374963
rect 494113 374929 494151 374963
rect 494185 374929 494223 374963
rect 494257 374929 494295 374963
rect 494329 374929 494367 374963
rect 494401 374929 494439 374963
rect 494473 374929 494511 374963
rect 494545 374929 494583 374963
rect 494617 374929 494633 374963
rect 493343 374923 494633 374929
rect 493048 374707 493091 374741
rect 493125 374707 493168 374741
rect 493048 374341 493168 374707
rect 494928 374741 495048 375107
rect 494928 374707 494971 374741
rect 495005 374707 495048 374741
rect 493343 374505 494633 374511
rect 493343 374471 493359 374505
rect 493393 374471 493431 374505
rect 493465 374471 493503 374505
rect 493537 374471 493575 374505
rect 493609 374471 493647 374505
rect 493681 374471 493719 374505
rect 493753 374471 493791 374505
rect 493825 374471 493863 374505
rect 493897 374471 493935 374505
rect 493969 374471 494007 374505
rect 494041 374471 494079 374505
rect 494113 374471 494151 374505
rect 494185 374471 494223 374505
rect 494257 374471 494295 374505
rect 494329 374471 494367 374505
rect 494401 374471 494439 374505
rect 494473 374471 494511 374505
rect 494545 374471 494583 374505
rect 494617 374471 494633 374505
rect 493343 374465 494633 374471
rect 493048 374307 493091 374341
rect 493125 374307 493168 374341
rect 493048 373941 493168 374307
rect 494928 374341 495048 374707
rect 494928 374307 494971 374341
rect 495005 374307 495048 374341
rect 493343 374047 494633 374053
rect 493343 374013 493359 374047
rect 493393 374013 493431 374047
rect 493465 374013 493503 374047
rect 493537 374013 493575 374047
rect 493609 374013 493647 374047
rect 493681 374013 493719 374047
rect 493753 374013 493791 374047
rect 493825 374013 493863 374047
rect 493897 374013 493935 374047
rect 493969 374013 494007 374047
rect 494041 374013 494079 374047
rect 494113 374013 494151 374047
rect 494185 374013 494223 374047
rect 494257 374013 494295 374047
rect 494329 374013 494367 374047
rect 494401 374013 494439 374047
rect 494473 374013 494511 374047
rect 494545 374013 494583 374047
rect 494617 374013 494633 374047
rect 493343 374007 494633 374013
rect 493048 373907 493091 373941
rect 493125 373907 493168 373941
rect 493048 373541 493168 373907
rect 494928 373941 495048 374307
rect 494928 373907 494971 373941
rect 495005 373907 495048 373941
rect 493343 373589 494633 373595
rect 493343 373555 493359 373589
rect 493393 373555 493431 373589
rect 493465 373555 493503 373589
rect 493537 373555 493575 373589
rect 493609 373555 493647 373589
rect 493681 373555 493719 373589
rect 493753 373555 493791 373589
rect 493825 373555 493863 373589
rect 493897 373555 493935 373589
rect 493969 373555 494007 373589
rect 494041 373555 494079 373589
rect 494113 373555 494151 373589
rect 494185 373555 494223 373589
rect 494257 373555 494295 373589
rect 494329 373555 494367 373589
rect 494401 373555 494439 373589
rect 494473 373555 494511 373589
rect 494545 373555 494583 373589
rect 494617 373555 494633 373589
rect 493343 373549 494633 373555
rect 493048 373507 493091 373541
rect 493125 373507 493168 373541
rect 493048 373141 493168 373507
rect 493048 373107 493091 373141
rect 493125 373107 493168 373141
rect 494928 373541 495048 373907
rect 494928 373507 494971 373541
rect 495005 373507 495048 373541
rect 494928 373141 495048 373507
rect 493048 372741 493168 373107
rect 493343 373131 494633 373137
rect 493343 373097 493359 373131
rect 493393 373097 493431 373131
rect 493465 373097 493503 373131
rect 493537 373097 493575 373131
rect 493609 373097 493647 373131
rect 493681 373097 493719 373131
rect 493753 373097 493791 373131
rect 493825 373097 493863 373131
rect 493897 373097 493935 373131
rect 493969 373097 494007 373131
rect 494041 373097 494079 373131
rect 494113 373097 494151 373131
rect 494185 373097 494223 373131
rect 494257 373097 494295 373131
rect 494329 373097 494367 373131
rect 494401 373097 494439 373131
rect 494473 373097 494511 373131
rect 494545 373097 494583 373131
rect 494617 373097 494633 373131
rect 493343 373091 494633 373097
rect 494928 373107 494971 373141
rect 495005 373107 495048 373141
rect 493048 372707 493091 372741
rect 493125 372707 493168 372741
rect 493048 372341 493168 372707
rect 494928 372741 495048 373107
rect 494928 372707 494971 372741
rect 495005 372707 495048 372741
rect 493343 372673 494633 372679
rect 493343 372639 493359 372673
rect 493393 372639 493431 372673
rect 493465 372639 493503 372673
rect 493537 372639 493575 372673
rect 493609 372639 493647 372673
rect 493681 372639 493719 372673
rect 493753 372639 493791 372673
rect 493825 372639 493863 372673
rect 493897 372639 493935 372673
rect 493969 372639 494007 372673
rect 494041 372639 494079 372673
rect 494113 372639 494151 372673
rect 494185 372639 494223 372673
rect 494257 372639 494295 372673
rect 494329 372639 494367 372673
rect 494401 372639 494439 372673
rect 494473 372639 494511 372673
rect 494545 372639 494583 372673
rect 494617 372639 494633 372673
rect 493343 372633 494633 372639
rect 493048 372307 493091 372341
rect 493125 372307 493168 372341
rect 493048 371941 493168 372307
rect 494928 372341 495048 372707
rect 494928 372307 494971 372341
rect 495005 372307 495048 372341
rect 493343 372215 494633 372221
rect 493343 372181 493359 372215
rect 493393 372181 493431 372215
rect 493465 372181 493503 372215
rect 493537 372181 493575 372215
rect 493609 372181 493647 372215
rect 493681 372181 493719 372215
rect 493753 372181 493791 372215
rect 493825 372181 493863 372215
rect 493897 372181 493935 372215
rect 493969 372181 494007 372215
rect 494041 372181 494079 372215
rect 494113 372181 494151 372215
rect 494185 372181 494223 372215
rect 494257 372181 494295 372215
rect 494329 372181 494367 372215
rect 494401 372181 494439 372215
rect 494473 372181 494511 372215
rect 494545 372181 494583 372215
rect 494617 372181 494633 372215
rect 493343 372175 494633 372181
rect 493048 371907 493091 371941
rect 493125 371907 493168 371941
rect 493048 371541 493168 371907
rect 494928 371941 495048 372307
rect 494928 371907 494971 371941
rect 495005 371907 495048 371941
rect 493343 371757 494633 371763
rect 493343 371723 493359 371757
rect 493393 371723 493431 371757
rect 493465 371723 493503 371757
rect 493537 371723 493575 371757
rect 493609 371723 493647 371757
rect 493681 371723 493719 371757
rect 493753 371723 493791 371757
rect 493825 371723 493863 371757
rect 493897 371723 493935 371757
rect 493969 371723 494007 371757
rect 494041 371723 494079 371757
rect 494113 371723 494151 371757
rect 494185 371723 494223 371757
rect 494257 371723 494295 371757
rect 494329 371723 494367 371757
rect 494401 371723 494439 371757
rect 494473 371723 494511 371757
rect 494545 371723 494583 371757
rect 494617 371723 494633 371757
rect 493343 371717 494633 371723
rect 493048 371507 493091 371541
rect 493125 371507 493168 371541
rect 493048 371141 493168 371507
rect 494928 371541 495048 371907
rect 494928 371507 494971 371541
rect 495005 371507 495048 371541
rect 493343 371299 494633 371305
rect 493343 371265 493359 371299
rect 493393 371265 493431 371299
rect 493465 371265 493503 371299
rect 493537 371265 493575 371299
rect 493609 371265 493647 371299
rect 493681 371265 493719 371299
rect 493753 371265 493791 371299
rect 493825 371265 493863 371299
rect 493897 371265 493935 371299
rect 493969 371265 494007 371299
rect 494041 371265 494079 371299
rect 494113 371265 494151 371299
rect 494185 371265 494223 371299
rect 494257 371265 494295 371299
rect 494329 371265 494367 371299
rect 494401 371265 494439 371299
rect 494473 371265 494511 371299
rect 494545 371265 494583 371299
rect 494617 371265 494633 371299
rect 493343 371259 494633 371265
rect 493048 371107 493091 371141
rect 493125 371107 493168 371141
rect 493048 370741 493168 371107
rect 494928 371141 495048 371507
rect 494928 371107 494971 371141
rect 495005 371107 495048 371141
rect 493343 370841 494633 370847
rect 493343 370807 493359 370841
rect 493393 370807 493431 370841
rect 493465 370807 493503 370841
rect 493537 370807 493575 370841
rect 493609 370807 493647 370841
rect 493681 370807 493719 370841
rect 493753 370807 493791 370841
rect 493825 370807 493863 370841
rect 493897 370807 493935 370841
rect 493969 370807 494007 370841
rect 494041 370807 494079 370841
rect 494113 370807 494151 370841
rect 494185 370807 494223 370841
rect 494257 370807 494295 370841
rect 494329 370807 494367 370841
rect 494401 370807 494439 370841
rect 494473 370807 494511 370841
rect 494545 370807 494583 370841
rect 494617 370807 494633 370841
rect 493343 370801 494633 370807
rect 493048 370707 493091 370741
rect 493125 370707 493168 370741
rect 493048 370341 493168 370707
rect 494928 370741 495048 371107
rect 494928 370707 494971 370741
rect 495005 370707 495048 370741
rect 493343 370383 494633 370389
rect 493343 370349 493359 370383
rect 493393 370349 493431 370383
rect 493465 370349 493503 370383
rect 493537 370349 493575 370383
rect 493609 370349 493647 370383
rect 493681 370349 493719 370383
rect 493753 370349 493791 370383
rect 493825 370349 493863 370383
rect 493897 370349 493935 370383
rect 493969 370349 494007 370383
rect 494041 370349 494079 370383
rect 494113 370349 494151 370383
rect 494185 370349 494223 370383
rect 494257 370349 494295 370383
rect 494329 370349 494367 370383
rect 494401 370349 494439 370383
rect 494473 370349 494511 370383
rect 494545 370349 494583 370383
rect 494617 370349 494633 370383
rect 493343 370343 494633 370349
rect 493048 370307 493091 370341
rect 493125 370307 493168 370341
rect 493048 369941 493168 370307
rect 493048 369907 493091 369941
rect 493125 369907 493168 369941
rect 494928 370341 495048 370707
rect 494928 370307 494971 370341
rect 495005 370307 495048 370341
rect 494928 369941 495048 370307
rect 493048 369541 493168 369907
rect 493343 369925 494633 369931
rect 493343 369891 493359 369925
rect 493393 369891 493431 369925
rect 493465 369891 493503 369925
rect 493537 369891 493575 369925
rect 493609 369891 493647 369925
rect 493681 369891 493719 369925
rect 493753 369891 493791 369925
rect 493825 369891 493863 369925
rect 493897 369891 493935 369925
rect 493969 369891 494007 369925
rect 494041 369891 494079 369925
rect 494113 369891 494151 369925
rect 494185 369891 494223 369925
rect 494257 369891 494295 369925
rect 494329 369891 494367 369925
rect 494401 369891 494439 369925
rect 494473 369891 494511 369925
rect 494545 369891 494583 369925
rect 494617 369891 494633 369925
rect 493343 369885 494633 369891
rect 494928 369907 494971 369941
rect 495005 369907 495048 369941
rect 493048 369507 493091 369541
rect 493125 369507 493168 369541
rect 493048 369141 493168 369507
rect 494928 369541 495048 369907
rect 494928 369507 494971 369541
rect 495005 369507 495048 369541
rect 493343 369467 494633 369473
rect 493343 369433 493359 369467
rect 493393 369433 493431 369467
rect 493465 369433 493503 369467
rect 493537 369433 493575 369467
rect 493609 369433 493647 369467
rect 493681 369433 493719 369467
rect 493753 369433 493791 369467
rect 493825 369433 493863 369467
rect 493897 369433 493935 369467
rect 493969 369433 494007 369467
rect 494041 369433 494079 369467
rect 494113 369433 494151 369467
rect 494185 369433 494223 369467
rect 494257 369433 494295 369467
rect 494329 369433 494367 369467
rect 494401 369433 494439 369467
rect 494473 369433 494511 369467
rect 494545 369433 494583 369467
rect 494617 369433 494633 369467
rect 493343 369427 494633 369433
rect 493048 369107 493091 369141
rect 493125 369107 493168 369141
rect 493048 368741 493168 369107
rect 494928 369141 495048 369507
rect 494928 369107 494971 369141
rect 495005 369107 495048 369141
rect 493343 369009 494633 369015
rect 493343 368975 493359 369009
rect 493393 368975 493431 369009
rect 493465 368975 493503 369009
rect 493537 368975 493575 369009
rect 493609 368975 493647 369009
rect 493681 368975 493719 369009
rect 493753 368975 493791 369009
rect 493825 368975 493863 369009
rect 493897 368975 493935 369009
rect 493969 368975 494007 369009
rect 494041 368975 494079 369009
rect 494113 368975 494151 369009
rect 494185 368975 494223 369009
rect 494257 368975 494295 369009
rect 494329 368975 494367 369009
rect 494401 368975 494439 369009
rect 494473 368975 494511 369009
rect 494545 368975 494583 369009
rect 494617 368975 494633 369009
rect 493343 368969 494633 368975
rect 493048 368707 493091 368741
rect 493125 368707 493168 368741
rect 493048 368341 493168 368707
rect 494928 368741 495048 369107
rect 494928 368707 494971 368741
rect 495005 368707 495048 368741
rect 493343 368551 494633 368557
rect 493343 368517 493359 368551
rect 493393 368517 493431 368551
rect 493465 368517 493503 368551
rect 493537 368517 493575 368551
rect 493609 368517 493647 368551
rect 493681 368517 493719 368551
rect 493753 368517 493791 368551
rect 493825 368517 493863 368551
rect 493897 368517 493935 368551
rect 493969 368517 494007 368551
rect 494041 368517 494079 368551
rect 494113 368517 494151 368551
rect 494185 368517 494223 368551
rect 494257 368517 494295 368551
rect 494329 368517 494367 368551
rect 494401 368517 494439 368551
rect 494473 368517 494511 368551
rect 494545 368517 494583 368551
rect 494617 368517 494633 368551
rect 493343 368511 494633 368517
rect 493048 368307 493091 368341
rect 493125 368307 493168 368341
rect 493048 367941 493168 368307
rect 494928 368341 495048 368707
rect 494928 368307 494971 368341
rect 495005 368307 495048 368341
rect 493343 368093 494633 368099
rect 493343 368059 493359 368093
rect 493393 368059 493431 368093
rect 493465 368059 493503 368093
rect 493537 368059 493575 368093
rect 493609 368059 493647 368093
rect 493681 368059 493719 368093
rect 493753 368059 493791 368093
rect 493825 368059 493863 368093
rect 493897 368059 493935 368093
rect 493969 368059 494007 368093
rect 494041 368059 494079 368093
rect 494113 368059 494151 368093
rect 494185 368059 494223 368093
rect 494257 368059 494295 368093
rect 494329 368059 494367 368093
rect 494401 368059 494439 368093
rect 494473 368059 494511 368093
rect 494545 368059 494583 368093
rect 494617 368059 494633 368093
rect 493343 368053 494633 368059
rect 493048 367907 493091 367941
rect 493125 367907 493168 367941
rect 493048 367541 493168 367907
rect 494928 367941 495048 368307
rect 494928 367907 494971 367941
rect 495005 367907 495048 367941
rect 493343 367635 494633 367641
rect 493343 367601 493359 367635
rect 493393 367601 493431 367635
rect 493465 367601 493503 367635
rect 493537 367601 493575 367635
rect 493609 367601 493647 367635
rect 493681 367601 493719 367635
rect 493753 367601 493791 367635
rect 493825 367601 493863 367635
rect 493897 367601 493935 367635
rect 493969 367601 494007 367635
rect 494041 367601 494079 367635
rect 494113 367601 494151 367635
rect 494185 367601 494223 367635
rect 494257 367601 494295 367635
rect 494329 367601 494367 367635
rect 494401 367601 494439 367635
rect 494473 367601 494511 367635
rect 494545 367601 494583 367635
rect 494617 367601 494633 367635
rect 493343 367595 494633 367601
rect 493048 367507 493091 367541
rect 493125 367507 493168 367541
rect 493048 367141 493168 367507
rect 494928 367541 495048 367907
rect 494928 367507 494971 367541
rect 495005 367507 495048 367541
rect 493048 367107 493091 367141
rect 493125 367107 493168 367141
rect 493343 367177 494633 367183
rect 493343 367143 493359 367177
rect 493393 367143 493431 367177
rect 493465 367143 493503 367177
rect 493537 367143 493575 367177
rect 493609 367143 493647 367177
rect 493681 367143 493719 367177
rect 493753 367143 493791 367177
rect 493825 367143 493863 367177
rect 493897 367143 493935 367177
rect 493969 367143 494007 367177
rect 494041 367143 494079 367177
rect 494113 367143 494151 367177
rect 494185 367143 494223 367177
rect 494257 367143 494295 367177
rect 494329 367143 494367 367177
rect 494401 367143 494439 367177
rect 494473 367143 494511 367177
rect 494545 367143 494583 367177
rect 494617 367143 494633 367177
rect 493343 367137 494633 367143
rect 494928 367141 495048 367507
rect 493048 366741 493168 367107
rect 493048 366707 493091 366741
rect 493125 366707 493168 366741
rect 494928 367107 494971 367141
rect 495005 367107 495048 367141
rect 494928 366741 495048 367107
rect 493048 366341 493168 366707
rect 493343 366719 494633 366725
rect 493343 366685 493359 366719
rect 493393 366685 493431 366719
rect 493465 366685 493503 366719
rect 493537 366685 493575 366719
rect 493609 366685 493647 366719
rect 493681 366685 493719 366719
rect 493753 366685 493791 366719
rect 493825 366685 493863 366719
rect 493897 366685 493935 366719
rect 493969 366685 494007 366719
rect 494041 366685 494079 366719
rect 494113 366685 494151 366719
rect 494185 366685 494223 366719
rect 494257 366685 494295 366719
rect 494329 366685 494367 366719
rect 494401 366685 494439 366719
rect 494473 366685 494511 366719
rect 494545 366685 494583 366719
rect 494617 366685 494633 366719
rect 493343 366679 494633 366685
rect 494928 366707 494971 366741
rect 495005 366707 495048 366741
rect 494536 366634 494588 366640
rect 494536 366576 494588 366582
rect 493048 366307 493091 366341
rect 493125 366307 493168 366341
rect 493048 365941 493168 366307
rect 494548 366267 494576 366576
rect 494928 366341 495048 366707
rect 494928 366307 494971 366341
rect 495005 366307 495048 366341
rect 493343 366261 494633 366267
rect 493343 366227 493359 366261
rect 493393 366227 493431 366261
rect 493465 366227 493503 366261
rect 493537 366227 493575 366261
rect 493609 366227 493647 366261
rect 493681 366227 493719 366261
rect 493753 366227 493791 366261
rect 493825 366227 493863 366261
rect 493897 366227 493935 366261
rect 493969 366227 494007 366261
rect 494041 366227 494079 366261
rect 494113 366227 494151 366261
rect 494185 366227 494223 366261
rect 494257 366227 494295 366261
rect 494329 366227 494367 366261
rect 494401 366227 494439 366261
rect 494473 366227 494511 366261
rect 494545 366227 494583 366261
rect 494617 366227 494633 366261
rect 493343 366221 494633 366227
rect 493048 365907 493091 365941
rect 493125 365907 493168 365941
rect 493048 365541 493168 365907
rect 494928 365941 495048 366307
rect 494928 365907 494971 365941
rect 495005 365907 495048 365941
rect 493343 365803 494633 365809
rect 493343 365769 493359 365803
rect 493393 365769 493431 365803
rect 493465 365769 493503 365803
rect 493537 365769 493575 365803
rect 493609 365769 493647 365803
rect 493681 365769 493719 365803
rect 493753 365769 493791 365803
rect 493825 365769 493863 365803
rect 493897 365769 493935 365803
rect 493969 365769 494007 365803
rect 494041 365769 494079 365803
rect 494113 365769 494151 365803
rect 494185 365769 494223 365803
rect 494257 365769 494295 365803
rect 494329 365769 494367 365803
rect 494401 365769 494439 365803
rect 494473 365769 494511 365803
rect 494545 365769 494583 365803
rect 494617 365769 494633 365803
rect 493343 365763 494633 365769
rect 493048 365507 493091 365541
rect 493125 365507 493168 365541
rect 493048 365141 493168 365507
rect 494928 365541 495048 365907
rect 494928 365507 494971 365541
rect 495005 365507 495048 365541
rect 493343 365345 494633 365351
rect 493343 365311 493359 365345
rect 493393 365311 493431 365345
rect 493465 365311 493503 365345
rect 493537 365311 493575 365345
rect 493609 365311 493647 365345
rect 493681 365311 493719 365345
rect 493753 365311 493791 365345
rect 493825 365311 493863 365345
rect 493897 365311 493935 365345
rect 493969 365311 494007 365345
rect 494041 365311 494079 365345
rect 494113 365311 494151 365345
rect 494185 365311 494223 365345
rect 494257 365311 494295 365345
rect 494329 365311 494367 365345
rect 494401 365311 494439 365345
rect 494473 365311 494511 365345
rect 494545 365311 494583 365345
rect 494617 365311 494633 365345
rect 493343 365305 494633 365311
rect 493048 365107 493091 365141
rect 493125 365107 493168 365141
rect 493048 364741 493168 365107
rect 494928 365141 495048 365507
rect 494928 365107 494971 365141
rect 495005 365107 495048 365141
rect 493343 364887 494633 364893
rect 493343 364853 493359 364887
rect 493393 364853 493431 364887
rect 493465 364853 493503 364887
rect 493537 364853 493575 364887
rect 493609 364853 493647 364887
rect 493681 364853 493719 364887
rect 493753 364853 493791 364887
rect 493825 364853 493863 364887
rect 493897 364853 493935 364887
rect 493969 364853 494007 364887
rect 494041 364853 494079 364887
rect 494113 364853 494151 364887
rect 494185 364853 494223 364887
rect 494257 364853 494295 364887
rect 494329 364853 494367 364887
rect 494401 364853 494439 364887
rect 494473 364853 494511 364887
rect 494545 364853 494583 364887
rect 494617 364853 494633 364887
rect 493343 364847 494633 364853
rect 493048 364707 493091 364741
rect 493125 364707 493168 364741
rect 493048 364341 493168 364707
rect 494928 364741 495048 365107
rect 494928 364707 494971 364741
rect 495005 364707 495048 364741
rect 493343 364429 494633 364435
rect 493343 364395 493359 364429
rect 493393 364395 493431 364429
rect 493465 364395 493503 364429
rect 493537 364395 493575 364429
rect 493609 364395 493647 364429
rect 493681 364395 493719 364429
rect 493753 364395 493791 364429
rect 493825 364395 493863 364429
rect 493897 364395 493935 364429
rect 493969 364395 494007 364429
rect 494041 364395 494079 364429
rect 494113 364395 494151 364429
rect 494185 364395 494223 364429
rect 494257 364395 494295 364429
rect 494329 364395 494367 364429
rect 494401 364395 494439 364429
rect 494473 364395 494511 364429
rect 494545 364395 494583 364429
rect 494617 364395 494633 364429
rect 493343 364389 494633 364395
rect 493048 364307 493091 364341
rect 493125 364307 493168 364341
rect 493048 363941 493168 364307
rect 494928 364341 495048 364707
rect 494928 364307 494971 364341
rect 495005 364307 495048 364341
rect 493048 363907 493091 363941
rect 493125 363907 493168 363941
rect 493343 363971 494633 363977
rect 493343 363937 493359 363971
rect 493393 363937 493431 363971
rect 493465 363937 493503 363971
rect 493537 363937 493575 363971
rect 493609 363937 493647 363971
rect 493681 363937 493719 363971
rect 493753 363937 493791 363971
rect 493825 363937 493863 363971
rect 493897 363937 493935 363971
rect 493969 363937 494007 363971
rect 494041 363937 494079 363971
rect 494113 363937 494151 363971
rect 494185 363937 494223 363971
rect 494257 363937 494295 363971
rect 494329 363937 494367 363971
rect 494401 363937 494439 363971
rect 494473 363937 494511 363971
rect 494545 363937 494583 363971
rect 494617 363937 494633 363971
rect 493343 363931 494633 363937
rect 494928 363941 495048 364307
rect 493048 363541 493168 363907
rect 493048 363507 493091 363541
rect 493125 363507 493168 363541
rect 494928 363907 494971 363941
rect 495005 363907 495048 363941
rect 494928 363541 495048 363907
rect 493048 363141 493168 363507
rect 493343 363513 494633 363519
rect 493343 363479 493359 363513
rect 493393 363479 493431 363513
rect 493465 363479 493503 363513
rect 493537 363479 493575 363513
rect 493609 363479 493647 363513
rect 493681 363479 493719 363513
rect 493753 363479 493791 363513
rect 493825 363479 493863 363513
rect 493897 363479 493935 363513
rect 493969 363479 494007 363513
rect 494041 363479 494079 363513
rect 494113 363479 494151 363513
rect 494185 363479 494223 363513
rect 494257 363479 494295 363513
rect 494329 363479 494367 363513
rect 494401 363479 494439 363513
rect 494473 363479 494511 363513
rect 494545 363479 494583 363513
rect 494617 363479 494633 363513
rect 493343 363473 494633 363479
rect 494928 363507 494971 363541
rect 495005 363507 495048 363541
rect 493048 363107 493091 363141
rect 493125 363107 493168 363141
rect 493048 362741 493168 363107
rect 494928 363141 495048 363507
rect 494928 363107 494971 363141
rect 495005 363107 495048 363141
rect 493343 363055 494633 363061
rect 493343 363021 493359 363055
rect 493393 363021 493431 363055
rect 493465 363021 493503 363055
rect 493537 363021 493575 363055
rect 493609 363021 493647 363055
rect 493681 363021 493719 363055
rect 493753 363021 493791 363055
rect 493825 363021 493863 363055
rect 493897 363021 493935 363055
rect 493969 363021 494007 363055
rect 494041 363021 494079 363055
rect 494113 363021 494151 363055
rect 494185 363021 494223 363055
rect 494257 363021 494295 363055
rect 494329 363021 494367 363055
rect 494401 363021 494439 363055
rect 494473 363021 494511 363055
rect 494545 363021 494583 363055
rect 494617 363021 494633 363055
rect 493343 363015 494633 363021
rect 493048 362707 493091 362741
rect 493125 362707 493168 362741
rect 493048 361476 493168 362707
rect 494928 362741 495048 363107
rect 494928 362707 494971 362741
rect 495005 362707 495048 362741
rect 493343 362597 494633 362603
rect 493343 362563 493359 362597
rect 493393 362563 493431 362597
rect 493465 362563 493503 362597
rect 493537 362563 493575 362597
rect 493609 362563 493647 362597
rect 493681 362563 493719 362597
rect 493753 362563 493791 362597
rect 493825 362563 493863 362597
rect 493897 362563 493935 362597
rect 493969 362563 494007 362597
rect 494041 362563 494079 362597
rect 494113 362563 494151 362597
rect 494185 362563 494223 362597
rect 494257 362563 494295 362597
rect 494329 362563 494367 362597
rect 494401 362563 494439 362597
rect 494473 362563 494511 362597
rect 494545 362563 494583 362597
rect 494617 362563 494633 362597
rect 493343 362557 494633 362563
rect 493048 359888 493050 361476
rect 493166 359888 493168 361476
rect 493048 359866 493168 359888
rect 491168 357440 491170 359028
rect 491286 357440 491288 359028
rect 491168 357418 491288 357440
rect 494928 359028 495048 362707
rect 496808 411584 496928 411606
rect 496808 409996 496810 411584
rect 496926 409996 496928 411584
rect 496808 408853 496928 409996
rect 496808 408819 496851 408853
rect 496885 408819 496928 408853
rect 496808 408453 496928 408819
rect 496808 408419 496851 408453
rect 496885 408419 496928 408453
rect 496808 408053 496928 408419
rect 496808 408019 496851 408053
rect 496885 408019 496928 408053
rect 496808 407653 496928 408019
rect 496808 407619 496851 407653
rect 496885 407619 496928 407653
rect 496808 407253 496928 407619
rect 496808 407219 496851 407253
rect 496885 407219 496928 407253
rect 496808 406853 496928 407219
rect 496808 406819 496851 406853
rect 496885 406819 496928 406853
rect 496808 406453 496928 406819
rect 496808 406419 496851 406453
rect 496885 406419 496928 406453
rect 496808 406053 496928 406419
rect 496808 406019 496851 406053
rect 496885 406019 496928 406053
rect 496808 405653 496928 406019
rect 496808 405619 496851 405653
rect 496885 405619 496928 405653
rect 496808 405253 496928 405619
rect 496808 405219 496851 405253
rect 496885 405219 496928 405253
rect 496808 404853 496928 405219
rect 496808 404819 496851 404853
rect 496885 404819 496928 404853
rect 496808 404453 496928 404819
rect 496808 404419 496851 404453
rect 496885 404419 496928 404453
rect 496808 404053 496928 404419
rect 496808 404019 496851 404053
rect 496885 404019 496928 404053
rect 496808 403653 496928 404019
rect 496808 403619 496851 403653
rect 496885 403619 496928 403653
rect 496808 403253 496928 403619
rect 496808 403219 496851 403253
rect 496885 403219 496928 403253
rect 496808 402853 496928 403219
rect 496808 402819 496851 402853
rect 496885 402819 496928 402853
rect 496808 402453 496928 402819
rect 496808 402419 496851 402453
rect 496885 402419 496928 402453
rect 496808 402053 496928 402419
rect 496808 402019 496851 402053
rect 496885 402019 496928 402053
rect 496808 400653 496928 402019
rect 498688 408853 498808 412444
rect 502448 414032 502568 414054
rect 502448 412444 502450 414032
rect 502566 412444 502568 414032
rect 498688 408819 498731 408853
rect 498765 408819 498808 408853
rect 498688 408453 498808 408819
rect 498688 408419 498731 408453
rect 498765 408419 498808 408453
rect 498688 408053 498808 408419
rect 498688 408019 498731 408053
rect 498765 408019 498808 408053
rect 498688 407653 498808 408019
rect 498688 407619 498731 407653
rect 498765 407619 498808 407653
rect 498688 407253 498808 407619
rect 498688 407219 498731 407253
rect 498765 407219 498808 407253
rect 498688 406853 498808 407219
rect 498688 406819 498731 406853
rect 498765 406819 498808 406853
rect 498688 406654 498808 406819
rect 498688 406602 498752 406654
rect 498804 406602 498808 406654
rect 498688 406453 498808 406602
rect 498688 406419 498731 406453
rect 498765 406419 498808 406453
rect 498688 406053 498808 406419
rect 498688 406019 498731 406053
rect 498765 406019 498808 406053
rect 498688 405653 498808 406019
rect 498688 405619 498731 405653
rect 498765 405619 498808 405653
rect 498688 405253 498808 405619
rect 498688 405219 498731 405253
rect 498765 405219 498808 405253
rect 498688 404853 498808 405219
rect 498688 404819 498731 404853
rect 498765 404819 498808 404853
rect 498688 404453 498808 404819
rect 498688 404419 498731 404453
rect 498765 404419 498808 404453
rect 498688 404053 498808 404419
rect 498688 404019 498731 404053
rect 498765 404019 498808 404053
rect 498688 403653 498808 404019
rect 498688 403619 498731 403653
rect 498765 403619 498808 403653
rect 498688 403253 498808 403619
rect 498688 403219 498731 403253
rect 498765 403219 498808 403253
rect 498688 402853 498808 403219
rect 498688 402819 498731 402853
rect 498765 402819 498808 402853
rect 498688 402453 498808 402819
rect 498688 402419 498731 402453
rect 498765 402419 498808 402453
rect 498688 402053 498808 402419
rect 498688 402019 498731 402053
rect 498765 402019 498808 402053
rect 497348 400824 498148 400830
rect 497348 400790 497371 400824
rect 497405 400790 497443 400824
rect 497477 400790 497515 400824
rect 497549 400790 497587 400824
rect 497621 400790 497659 400824
rect 497693 400790 497731 400824
rect 497765 400790 497803 400824
rect 497837 400790 497875 400824
rect 497909 400790 497947 400824
rect 497981 400790 498019 400824
rect 498053 400790 498091 400824
rect 498125 400790 498148 400824
rect 497348 400784 498148 400790
rect 496808 400619 496851 400653
rect 496885 400619 496928 400653
rect 498688 400653 498808 402019
rect 496808 399741 496928 400619
rect 498356 400588 498384 400643
rect 498688 400619 498731 400653
rect 498765 400619 498808 400653
rect 498344 400582 498396 400588
rect 498344 400524 498396 400530
rect 498560 400404 498588 400459
rect 498548 400398 498600 400404
rect 497348 400366 498148 400372
rect 497348 400332 497371 400366
rect 497405 400332 497443 400366
rect 497477 400332 497515 400366
rect 497549 400332 497587 400366
rect 497621 400332 497659 400366
rect 497693 400332 497731 400366
rect 497765 400332 497803 400366
rect 497837 400332 497875 400366
rect 497909 400332 497947 400366
rect 497981 400332 498019 400366
rect 498053 400332 498091 400366
rect 498125 400332 498148 400366
rect 498548 400340 498600 400346
rect 497348 400326 498148 400332
rect 498084 400294 498112 400326
rect 498688 400294 498808 400619
rect 498084 400266 498808 400294
rect 498492 399944 498520 399999
rect 498480 399938 498532 399944
rect 497103 399877 498393 399883
rect 498480 399880 498532 399886
rect 497103 399843 497119 399877
rect 497153 399843 497191 399877
rect 497225 399843 497263 399877
rect 497297 399843 497335 399877
rect 497369 399843 497407 399877
rect 497441 399843 497479 399877
rect 497513 399843 497551 399877
rect 497585 399843 497623 399877
rect 497657 399843 497695 399877
rect 497729 399843 497767 399877
rect 497801 399843 497839 399877
rect 497873 399843 497911 399877
rect 497945 399843 497983 399877
rect 498017 399843 498055 399877
rect 498089 399843 498127 399877
rect 498161 399843 498199 399877
rect 498233 399843 498271 399877
rect 498305 399843 498343 399877
rect 498377 399843 498393 399877
rect 497103 399837 498393 399843
rect 496808 399707 496851 399741
rect 496885 399707 496928 399741
rect 496808 399341 496928 399707
rect 498688 399741 498808 400266
rect 498688 399707 498731 399741
rect 498765 399707 498808 399741
rect 497103 399419 498393 399425
rect 497103 399385 497119 399419
rect 497153 399385 497191 399419
rect 497225 399385 497263 399419
rect 497297 399385 497335 399419
rect 497369 399385 497407 399419
rect 497441 399385 497479 399419
rect 497513 399385 497551 399419
rect 497585 399385 497623 399419
rect 497657 399385 497695 399419
rect 497729 399385 497767 399419
rect 497801 399385 497839 399419
rect 497873 399385 497911 399419
rect 497945 399385 497983 399419
rect 498017 399385 498055 399419
rect 498089 399385 498127 399419
rect 498161 399385 498199 399419
rect 498233 399385 498271 399419
rect 498305 399385 498343 399419
rect 498377 399385 498393 399419
rect 497103 399379 498393 399385
rect 496808 399307 496851 399341
rect 496885 399307 496928 399341
rect 496808 398941 496928 399307
rect 498688 399341 498808 399707
rect 498688 399307 498731 399341
rect 498765 399307 498808 399341
rect 496808 398907 496851 398941
rect 496885 398907 496928 398941
rect 497103 398961 498393 398967
rect 497103 398927 497119 398961
rect 497153 398927 497191 398961
rect 497225 398927 497263 398961
rect 497297 398927 497335 398961
rect 497369 398927 497407 398961
rect 497441 398927 497479 398961
rect 497513 398927 497551 398961
rect 497585 398927 497623 398961
rect 497657 398927 497695 398961
rect 497729 398927 497767 398961
rect 497801 398927 497839 398961
rect 497873 398927 497911 398961
rect 497945 398927 497983 398961
rect 498017 398927 498055 398961
rect 498089 398927 498127 398961
rect 498161 398927 498199 398961
rect 498233 398927 498271 398961
rect 498305 398927 498343 398961
rect 498377 398927 498393 398961
rect 497103 398921 498393 398927
rect 498688 398941 498808 399307
rect 496808 398541 496928 398907
rect 496808 398507 496851 398541
rect 496885 398507 496928 398541
rect 498688 398907 498731 398941
rect 498765 398907 498808 398941
rect 498688 398541 498808 398907
rect 496808 398141 496928 398507
rect 497103 398503 498393 398509
rect 497103 398469 497119 398503
rect 497153 398469 497191 398503
rect 497225 398469 497263 398503
rect 497297 398469 497335 398503
rect 497369 398469 497407 398503
rect 497441 398469 497479 398503
rect 497513 398469 497551 398503
rect 497585 398469 497623 398503
rect 497657 398469 497695 398503
rect 497729 398469 497767 398503
rect 497801 398469 497839 398503
rect 497873 398469 497911 398503
rect 497945 398469 497983 398503
rect 498017 398469 498055 398503
rect 498089 398469 498127 398503
rect 498161 398469 498199 398503
rect 498233 398469 498271 398503
rect 498305 398469 498343 398503
rect 498377 398469 498393 398503
rect 497103 398463 498393 398469
rect 498688 398507 498731 398541
rect 498765 398507 498808 398541
rect 496808 398107 496851 398141
rect 496885 398107 496928 398141
rect 496808 397741 496928 398107
rect 498688 398141 498808 398507
rect 498688 398107 498731 398141
rect 498765 398107 498808 398141
rect 497103 398045 498393 398051
rect 497103 398011 497119 398045
rect 497153 398011 497191 398045
rect 497225 398011 497263 398045
rect 497297 398011 497335 398045
rect 497369 398011 497407 398045
rect 497441 398011 497479 398045
rect 497513 398011 497551 398045
rect 497585 398011 497623 398045
rect 497657 398011 497695 398045
rect 497729 398011 497767 398045
rect 497801 398011 497839 398045
rect 497873 398011 497911 398045
rect 497945 398011 497983 398045
rect 498017 398011 498055 398045
rect 498089 398011 498127 398045
rect 498161 398011 498199 398045
rect 498233 398011 498271 398045
rect 498305 398011 498343 398045
rect 498377 398011 498393 398045
rect 497103 398005 498393 398011
rect 496808 397707 496851 397741
rect 496885 397707 496928 397741
rect 496808 397341 496928 397707
rect 498688 397741 498808 398107
rect 498688 397707 498731 397741
rect 498765 397707 498808 397741
rect 497103 397587 498393 397593
rect 497103 397553 497119 397587
rect 497153 397553 497191 397587
rect 497225 397553 497263 397587
rect 497297 397553 497335 397587
rect 497369 397553 497407 397587
rect 497441 397553 497479 397587
rect 497513 397553 497551 397587
rect 497585 397553 497623 397587
rect 497657 397553 497695 397587
rect 497729 397553 497767 397587
rect 497801 397553 497839 397587
rect 497873 397553 497911 397587
rect 497945 397553 497983 397587
rect 498017 397553 498055 397587
rect 498089 397553 498127 397587
rect 498161 397553 498199 397587
rect 498233 397553 498271 397587
rect 498305 397553 498343 397587
rect 498377 397553 498393 397587
rect 497103 397547 498393 397553
rect 496808 397307 496851 397341
rect 496885 397307 496928 397341
rect 496808 396941 496928 397307
rect 498688 397341 498808 397707
rect 498688 397307 498731 397341
rect 498765 397307 498808 397341
rect 497103 397129 498393 397135
rect 497103 397095 497119 397129
rect 497153 397095 497191 397129
rect 497225 397095 497263 397129
rect 497297 397095 497335 397129
rect 497369 397095 497407 397129
rect 497441 397095 497479 397129
rect 497513 397095 497551 397129
rect 497585 397095 497623 397129
rect 497657 397095 497695 397129
rect 497729 397095 497767 397129
rect 497801 397095 497839 397129
rect 497873 397095 497911 397129
rect 497945 397095 497983 397129
rect 498017 397095 498055 397129
rect 498089 397095 498127 397129
rect 498161 397095 498199 397129
rect 498233 397095 498271 397129
rect 498305 397095 498343 397129
rect 498377 397095 498393 397129
rect 497103 397089 498393 397095
rect 496808 396907 496851 396941
rect 496885 396907 496928 396941
rect 496808 396541 496928 396907
rect 498688 396941 498808 397307
rect 498688 396907 498731 396941
rect 498765 396907 498808 396941
rect 497103 396671 498393 396677
rect 497103 396637 497119 396671
rect 497153 396637 497191 396671
rect 497225 396637 497263 396671
rect 497297 396637 497335 396671
rect 497369 396637 497407 396671
rect 497441 396637 497479 396671
rect 497513 396637 497551 396671
rect 497585 396637 497623 396671
rect 497657 396637 497695 396671
rect 497729 396637 497767 396671
rect 497801 396637 497839 396671
rect 497873 396637 497911 396671
rect 497945 396637 497983 396671
rect 498017 396637 498055 396671
rect 498089 396637 498127 396671
rect 498161 396637 498199 396671
rect 498233 396637 498271 396671
rect 498305 396637 498343 396671
rect 498377 396637 498393 396671
rect 497103 396631 498393 396637
rect 496808 396507 496851 396541
rect 496885 396507 496928 396541
rect 496808 396141 496928 396507
rect 498688 396541 498808 396907
rect 498688 396507 498731 396541
rect 498765 396507 498808 396541
rect 497103 396213 498393 396219
rect 497103 396179 497119 396213
rect 497153 396179 497191 396213
rect 497225 396179 497263 396213
rect 497297 396179 497335 396213
rect 497369 396179 497407 396213
rect 497441 396179 497479 396213
rect 497513 396179 497551 396213
rect 497585 396179 497623 396213
rect 497657 396179 497695 396213
rect 497729 396179 497767 396213
rect 497801 396179 497839 396213
rect 497873 396179 497911 396213
rect 497945 396179 497983 396213
rect 498017 396179 498055 396213
rect 498089 396179 498127 396213
rect 498161 396179 498199 396213
rect 498233 396179 498271 396213
rect 498305 396179 498343 396213
rect 498377 396179 498393 396213
rect 497103 396173 498393 396179
rect 496808 396107 496851 396141
rect 496885 396107 496928 396141
rect 496808 395741 496928 396107
rect 498688 396141 498808 396507
rect 498688 396107 498731 396141
rect 498765 396107 498808 396141
rect 496808 395707 496851 395741
rect 496885 395707 496928 395741
rect 497103 395755 498393 395761
rect 497103 395721 497119 395755
rect 497153 395721 497191 395755
rect 497225 395721 497263 395755
rect 497297 395721 497335 395755
rect 497369 395721 497407 395755
rect 497441 395721 497479 395755
rect 497513 395721 497551 395755
rect 497585 395721 497623 395755
rect 497657 395721 497695 395755
rect 497729 395721 497767 395755
rect 497801 395721 497839 395755
rect 497873 395721 497911 395755
rect 497945 395721 497983 395755
rect 498017 395721 498055 395755
rect 498089 395721 498127 395755
rect 498161 395721 498199 395755
rect 498233 395721 498271 395755
rect 498305 395721 498343 395755
rect 498377 395721 498393 395755
rect 497103 395715 498393 395721
rect 498688 395741 498808 396107
rect 496808 395341 496928 395707
rect 496808 395307 496851 395341
rect 496885 395307 496928 395341
rect 496808 394941 496928 395307
rect 498688 395707 498731 395741
rect 498765 395707 498808 395741
rect 498688 395341 498808 395707
rect 498688 395307 498731 395341
rect 498765 395307 498808 395341
rect 497103 395297 498393 395303
rect 497103 395263 497119 395297
rect 497153 395263 497191 395297
rect 497225 395263 497263 395297
rect 497297 395263 497335 395297
rect 497369 395263 497407 395297
rect 497441 395263 497479 395297
rect 497513 395263 497551 395297
rect 497585 395263 497623 395297
rect 497657 395263 497695 395297
rect 497729 395263 497767 395297
rect 497801 395263 497839 395297
rect 497873 395263 497911 395297
rect 497945 395263 497983 395297
rect 498017 395263 498055 395297
rect 498089 395263 498127 395297
rect 498161 395263 498199 395297
rect 498233 395263 498271 395297
rect 498305 395263 498343 395297
rect 498377 395263 498393 395297
rect 497103 395257 498393 395263
rect 496808 394907 496851 394941
rect 496885 394907 496928 394941
rect 496808 394541 496928 394907
rect 498688 394941 498808 395307
rect 498688 394907 498731 394941
rect 498765 394907 498808 394941
rect 497103 394839 498393 394845
rect 497103 394805 497119 394839
rect 497153 394805 497191 394839
rect 497225 394805 497263 394839
rect 497297 394805 497335 394839
rect 497369 394805 497407 394839
rect 497441 394805 497479 394839
rect 497513 394805 497551 394839
rect 497585 394805 497623 394839
rect 497657 394805 497695 394839
rect 497729 394805 497767 394839
rect 497801 394805 497839 394839
rect 497873 394805 497911 394839
rect 497945 394805 497983 394839
rect 498017 394805 498055 394839
rect 498089 394805 498127 394839
rect 498161 394805 498199 394839
rect 498233 394805 498271 394839
rect 498305 394805 498343 394839
rect 498377 394805 498393 394839
rect 497103 394799 498393 394805
rect 496808 394507 496851 394541
rect 496885 394507 496928 394541
rect 496808 394141 496928 394507
rect 498688 394541 498808 394907
rect 498688 394507 498731 394541
rect 498765 394507 498808 394541
rect 497103 394381 498393 394387
rect 497103 394347 497119 394381
rect 497153 394347 497191 394381
rect 497225 394347 497263 394381
rect 497297 394347 497335 394381
rect 497369 394347 497407 394381
rect 497441 394347 497479 394381
rect 497513 394347 497551 394381
rect 497585 394347 497623 394381
rect 497657 394347 497695 394381
rect 497729 394347 497767 394381
rect 497801 394347 497839 394381
rect 497873 394347 497911 394381
rect 497945 394347 497983 394381
rect 498017 394347 498055 394381
rect 498089 394347 498127 394381
rect 498161 394347 498199 394381
rect 498233 394347 498271 394381
rect 498305 394347 498343 394381
rect 498377 394347 498393 394381
rect 497103 394341 498393 394347
rect 496808 394107 496851 394141
rect 496885 394107 496928 394141
rect 496808 393741 496928 394107
rect 498688 394141 498808 394507
rect 498688 394107 498731 394141
rect 498765 394107 498808 394141
rect 497103 393923 498393 393929
rect 497103 393889 497119 393923
rect 497153 393889 497191 393923
rect 497225 393889 497263 393923
rect 497297 393889 497335 393923
rect 497369 393889 497407 393923
rect 497441 393889 497479 393923
rect 497513 393889 497551 393923
rect 497585 393889 497623 393923
rect 497657 393889 497695 393923
rect 497729 393889 497767 393923
rect 497801 393889 497839 393923
rect 497873 393889 497911 393923
rect 497945 393889 497983 393923
rect 498017 393889 498055 393923
rect 498089 393889 498127 393923
rect 498161 393889 498199 393923
rect 498233 393889 498271 393923
rect 498305 393889 498343 393923
rect 498377 393889 498393 393923
rect 497103 393883 498393 393889
rect 496808 393707 496851 393741
rect 496885 393707 496928 393741
rect 496808 393341 496928 393707
rect 498688 393741 498808 394107
rect 498688 393707 498731 393741
rect 498765 393707 498808 393741
rect 497103 393465 498393 393471
rect 497103 393431 497119 393465
rect 497153 393431 497191 393465
rect 497225 393431 497263 393465
rect 497297 393431 497335 393465
rect 497369 393431 497407 393465
rect 497441 393431 497479 393465
rect 497513 393431 497551 393465
rect 497585 393431 497623 393465
rect 497657 393431 497695 393465
rect 497729 393431 497767 393465
rect 497801 393431 497839 393465
rect 497873 393431 497911 393465
rect 497945 393431 497983 393465
rect 498017 393431 498055 393465
rect 498089 393431 498127 393465
rect 498161 393431 498199 393465
rect 498233 393431 498271 393465
rect 498305 393431 498343 393465
rect 498377 393431 498393 393465
rect 497103 393425 498393 393431
rect 496808 393307 496851 393341
rect 496885 393307 496928 393341
rect 496808 392941 496928 393307
rect 498688 393341 498808 393707
rect 498688 393307 498731 393341
rect 498765 393307 498808 393341
rect 497103 393007 498393 393013
rect 497103 392973 497119 393007
rect 497153 392973 497191 393007
rect 497225 392973 497263 393007
rect 497297 392973 497335 393007
rect 497369 392973 497407 393007
rect 497441 392973 497479 393007
rect 497513 392973 497551 393007
rect 497585 392973 497623 393007
rect 497657 392973 497695 393007
rect 497729 392973 497767 393007
rect 497801 392973 497839 393007
rect 497873 392973 497911 393007
rect 497945 392973 497983 393007
rect 498017 392973 498055 393007
rect 498089 392973 498127 393007
rect 498161 392973 498199 393007
rect 498233 392973 498271 393007
rect 498305 392973 498343 393007
rect 498377 392973 498393 393007
rect 497103 392967 498393 392973
rect 496808 392907 496851 392941
rect 496885 392907 496928 392941
rect 496808 392541 496928 392907
rect 498688 392941 498808 393307
rect 498688 392907 498731 392941
rect 498765 392907 498808 392941
rect 498344 392762 498396 392768
rect 498344 392704 498396 392710
rect 498356 392555 498384 392704
rect 496808 392507 496851 392541
rect 496885 392507 496928 392541
rect 497103 392549 498393 392555
rect 497103 392515 497119 392549
rect 497153 392515 497191 392549
rect 497225 392515 497263 392549
rect 497297 392515 497335 392549
rect 497369 392515 497407 392549
rect 497441 392515 497479 392549
rect 497513 392515 497551 392549
rect 497585 392515 497623 392549
rect 497657 392515 497695 392549
rect 497729 392515 497767 392549
rect 497801 392515 497839 392549
rect 497873 392515 497911 392549
rect 497945 392515 497983 392549
rect 498017 392515 498055 392549
rect 498089 392515 498127 392549
rect 498161 392515 498199 392549
rect 498233 392515 498271 392549
rect 498305 392515 498343 392549
rect 498377 392515 498393 392549
rect 497103 392509 498393 392515
rect 498688 392541 498808 392907
rect 496808 392141 496928 392507
rect 496808 392107 496851 392141
rect 496885 392107 496928 392141
rect 496808 391741 496928 392107
rect 498688 392507 498731 392541
rect 498765 392507 498808 392541
rect 498688 392141 498808 392507
rect 498688 392107 498731 392141
rect 498765 392107 498808 392141
rect 497103 392091 498393 392097
rect 497103 392057 497119 392091
rect 497153 392057 497191 392091
rect 497225 392057 497263 392091
rect 497297 392057 497335 392091
rect 497369 392057 497407 392091
rect 497441 392057 497479 392091
rect 497513 392057 497551 392091
rect 497585 392057 497623 392091
rect 497657 392057 497695 392091
rect 497729 392057 497767 392091
rect 497801 392057 497839 392091
rect 497873 392057 497911 392091
rect 497945 392057 497983 392091
rect 498017 392057 498055 392091
rect 498089 392057 498127 392091
rect 498161 392057 498199 392091
rect 498233 392057 498271 392091
rect 498305 392057 498343 392091
rect 498377 392057 498393 392091
rect 497103 392051 498393 392057
rect 496808 391707 496851 391741
rect 496885 391707 496928 391741
rect 496808 391341 496928 391707
rect 498688 391741 498808 392107
rect 498688 391707 498731 391741
rect 498765 391707 498808 391741
rect 497103 391633 498393 391639
rect 497103 391599 497119 391633
rect 497153 391599 497191 391633
rect 497225 391599 497263 391633
rect 497297 391599 497335 391633
rect 497369 391599 497407 391633
rect 497441 391599 497479 391633
rect 497513 391599 497551 391633
rect 497585 391599 497623 391633
rect 497657 391599 497695 391633
rect 497729 391599 497767 391633
rect 497801 391599 497839 391633
rect 497873 391599 497911 391633
rect 497945 391599 497983 391633
rect 498017 391599 498055 391633
rect 498089 391599 498127 391633
rect 498161 391599 498199 391633
rect 498233 391599 498271 391633
rect 498305 391599 498343 391633
rect 498377 391599 498393 391633
rect 497103 391593 498393 391599
rect 496808 391307 496851 391341
rect 496885 391307 496928 391341
rect 496808 390941 496928 391307
rect 498688 391341 498808 391707
rect 498688 391307 498731 391341
rect 498765 391307 498808 391341
rect 497103 391175 498393 391181
rect 497103 391141 497119 391175
rect 497153 391141 497191 391175
rect 497225 391141 497263 391175
rect 497297 391141 497335 391175
rect 497369 391141 497407 391175
rect 497441 391141 497479 391175
rect 497513 391141 497551 391175
rect 497585 391141 497623 391175
rect 497657 391141 497695 391175
rect 497729 391141 497767 391175
rect 497801 391141 497839 391175
rect 497873 391141 497911 391175
rect 497945 391141 497983 391175
rect 498017 391141 498055 391175
rect 498089 391141 498127 391175
rect 498161 391141 498199 391175
rect 498233 391141 498271 391175
rect 498305 391141 498343 391175
rect 498377 391141 498393 391175
rect 497103 391135 498393 391141
rect 496808 390907 496851 390941
rect 496885 390907 496928 390941
rect 496808 390541 496928 390907
rect 498688 390941 498808 391307
rect 498688 390907 498731 390941
rect 498765 390907 498808 390941
rect 497103 390717 498393 390723
rect 497103 390683 497119 390717
rect 497153 390683 497191 390717
rect 497225 390683 497263 390717
rect 497297 390683 497335 390717
rect 497369 390683 497407 390717
rect 497441 390683 497479 390717
rect 497513 390683 497551 390717
rect 497585 390683 497623 390717
rect 497657 390683 497695 390717
rect 497729 390683 497767 390717
rect 497801 390683 497839 390717
rect 497873 390683 497911 390717
rect 497945 390683 497983 390717
rect 498017 390683 498055 390717
rect 498089 390683 498127 390717
rect 498161 390683 498199 390717
rect 498233 390683 498271 390717
rect 498305 390683 498343 390717
rect 498377 390683 498393 390717
rect 497103 390677 498393 390683
rect 496808 390507 496851 390541
rect 496885 390507 496928 390541
rect 496808 390141 496928 390507
rect 498688 390541 498808 390907
rect 498688 390507 498731 390541
rect 498765 390507 498808 390541
rect 497103 390259 498393 390265
rect 497103 390225 497119 390259
rect 497153 390225 497191 390259
rect 497225 390225 497263 390259
rect 497297 390225 497335 390259
rect 497369 390225 497407 390259
rect 497441 390225 497479 390259
rect 497513 390225 497551 390259
rect 497585 390225 497623 390259
rect 497657 390225 497695 390259
rect 497729 390225 497767 390259
rect 497801 390225 497839 390259
rect 497873 390225 497911 390259
rect 497945 390225 497983 390259
rect 498017 390225 498055 390259
rect 498089 390225 498127 390259
rect 498161 390225 498199 390259
rect 498233 390225 498271 390259
rect 498305 390225 498343 390259
rect 498377 390225 498393 390259
rect 497103 390219 498393 390225
rect 496808 390107 496851 390141
rect 496885 390107 496928 390141
rect 496808 389741 496928 390107
rect 498688 390141 498808 390507
rect 498688 390107 498731 390141
rect 498765 390107 498808 390141
rect 497103 389801 498393 389807
rect 497103 389767 497119 389801
rect 497153 389767 497191 389801
rect 497225 389767 497263 389801
rect 497297 389767 497335 389801
rect 497369 389767 497407 389801
rect 497441 389767 497479 389801
rect 497513 389767 497551 389801
rect 497585 389767 497623 389801
rect 497657 389767 497695 389801
rect 497729 389767 497767 389801
rect 497801 389767 497839 389801
rect 497873 389767 497911 389801
rect 497945 389767 497983 389801
rect 498017 389767 498055 389801
rect 498089 389767 498127 389801
rect 498161 389767 498199 389801
rect 498233 389767 498271 389801
rect 498305 389767 498343 389801
rect 498377 389767 498393 389801
rect 497103 389761 498393 389767
rect 496808 389707 496851 389741
rect 496885 389707 496928 389741
rect 496808 389346 496928 389707
rect 498688 389741 498808 390107
rect 498688 389707 498731 389741
rect 498765 389707 498808 389741
rect 497103 389346 498393 389349
rect 496808 389343 498393 389346
rect 496808 389341 497119 389343
rect 496808 389307 496851 389341
rect 496885 389318 497119 389341
rect 496885 389307 496928 389318
rect 496808 388941 496928 389307
rect 497103 389309 497119 389318
rect 497153 389309 497191 389343
rect 497225 389309 497263 389343
rect 497297 389309 497335 389343
rect 497369 389309 497407 389343
rect 497441 389309 497479 389343
rect 497513 389309 497551 389343
rect 497585 389309 497623 389343
rect 497657 389309 497695 389343
rect 497729 389309 497767 389343
rect 497801 389309 497839 389343
rect 497873 389309 497911 389343
rect 497945 389309 497983 389343
rect 498017 389309 498055 389343
rect 498089 389309 498127 389343
rect 498161 389309 498199 389343
rect 498233 389309 498271 389343
rect 498305 389309 498343 389343
rect 498377 389309 498393 389343
rect 497103 389303 498393 389309
rect 498688 389341 498808 389707
rect 498688 389307 498731 389341
rect 498765 389307 498808 389341
rect 496808 388907 496851 388941
rect 496885 388907 496928 388941
rect 496808 388541 496928 388907
rect 498688 388941 498808 389307
rect 498688 388907 498731 388941
rect 498765 388907 498808 388941
rect 497103 388885 498393 388891
rect 497103 388851 497119 388885
rect 497153 388851 497191 388885
rect 497225 388851 497263 388885
rect 497297 388851 497335 388885
rect 497369 388851 497407 388885
rect 497441 388851 497479 388885
rect 497513 388851 497551 388885
rect 497585 388851 497623 388885
rect 497657 388851 497695 388885
rect 497729 388851 497767 388885
rect 497801 388851 497839 388885
rect 497873 388851 497911 388885
rect 497945 388851 497983 388885
rect 498017 388851 498055 388885
rect 498089 388851 498127 388885
rect 498161 388851 498199 388885
rect 498233 388851 498271 388885
rect 498305 388851 498343 388885
rect 498377 388851 498393 388885
rect 497103 388845 498393 388851
rect 496808 388507 496851 388541
rect 496885 388507 496928 388541
rect 496808 388141 496928 388507
rect 498688 388541 498808 388907
rect 498688 388507 498731 388541
rect 498765 388507 498808 388541
rect 497103 388427 498393 388433
rect 497103 388393 497119 388427
rect 497153 388393 497191 388427
rect 497225 388393 497263 388427
rect 497297 388393 497335 388427
rect 497369 388393 497407 388427
rect 497441 388393 497479 388427
rect 497513 388393 497551 388427
rect 497585 388393 497623 388427
rect 497657 388393 497695 388427
rect 497729 388393 497767 388427
rect 497801 388393 497839 388427
rect 497873 388393 497911 388427
rect 497945 388393 497983 388427
rect 498017 388393 498055 388427
rect 498089 388393 498127 388427
rect 498161 388393 498199 388427
rect 498233 388393 498271 388427
rect 498305 388393 498343 388427
rect 498377 388393 498393 388427
rect 497103 388387 498393 388393
rect 496808 388107 496851 388141
rect 496885 388107 496928 388141
rect 496808 387741 496928 388107
rect 498688 388141 498808 388507
rect 498688 388107 498731 388141
rect 498765 388107 498808 388141
rect 497103 387969 498393 387975
rect 497103 387935 497119 387969
rect 497153 387935 497191 387969
rect 497225 387935 497263 387969
rect 497297 387935 497335 387969
rect 497369 387935 497407 387969
rect 497441 387935 497479 387969
rect 497513 387935 497551 387969
rect 497585 387935 497623 387969
rect 497657 387935 497695 387969
rect 497729 387935 497767 387969
rect 497801 387935 497839 387969
rect 497873 387935 497911 387969
rect 497945 387935 497983 387969
rect 498017 387935 498055 387969
rect 498089 387935 498127 387969
rect 498161 387935 498199 387969
rect 498233 387935 498271 387969
rect 498305 387935 498343 387969
rect 498377 387935 498393 387969
rect 497103 387929 498393 387935
rect 496808 387707 496851 387741
rect 496885 387707 496928 387741
rect 496808 387341 496928 387707
rect 498688 387741 498808 388107
rect 498688 387707 498731 387741
rect 498765 387707 498808 387741
rect 497103 387511 498393 387517
rect 497103 387477 497119 387511
rect 497153 387477 497191 387511
rect 497225 387477 497263 387511
rect 497297 387477 497335 387511
rect 497369 387477 497407 387511
rect 497441 387477 497479 387511
rect 497513 387477 497551 387511
rect 497585 387477 497623 387511
rect 497657 387477 497695 387511
rect 497729 387477 497767 387511
rect 497801 387477 497839 387511
rect 497873 387477 497911 387511
rect 497945 387477 497983 387511
rect 498017 387477 498055 387511
rect 498089 387477 498127 387511
rect 498161 387477 498199 387511
rect 498233 387477 498271 387511
rect 498305 387477 498343 387511
rect 498377 387477 498393 387511
rect 497103 387471 498393 387477
rect 496808 387307 496851 387341
rect 496885 387307 496928 387341
rect 496808 386941 496928 387307
rect 498688 387341 498808 387707
rect 498688 387307 498731 387341
rect 498765 387307 498808 387341
rect 497103 387053 498393 387059
rect 497103 387019 497119 387053
rect 497153 387019 497191 387053
rect 497225 387019 497263 387053
rect 497297 387019 497335 387053
rect 497369 387019 497407 387053
rect 497441 387019 497479 387053
rect 497513 387019 497551 387053
rect 497585 387019 497623 387053
rect 497657 387019 497695 387053
rect 497729 387019 497767 387053
rect 497801 387019 497839 387053
rect 497873 387019 497911 387053
rect 497945 387019 497983 387053
rect 498017 387019 498055 387053
rect 498089 387019 498127 387053
rect 498161 387019 498199 387053
rect 498233 387019 498271 387053
rect 498305 387019 498343 387053
rect 498377 387019 498393 387053
rect 497103 387013 498393 387019
rect 496808 386907 496851 386941
rect 496885 386907 496928 386941
rect 496808 386541 496928 386907
rect 498688 386941 498808 387307
rect 498688 386907 498731 386941
rect 498765 386907 498808 386941
rect 497103 386595 498393 386601
rect 497103 386561 497119 386595
rect 497153 386561 497191 386595
rect 497225 386561 497263 386595
rect 497297 386561 497335 386595
rect 497369 386561 497407 386595
rect 497441 386561 497479 386595
rect 497513 386561 497551 386595
rect 497585 386561 497623 386595
rect 497657 386561 497695 386595
rect 497729 386561 497767 386595
rect 497801 386561 497839 386595
rect 497873 386561 497911 386595
rect 497945 386561 497983 386595
rect 498017 386561 498055 386595
rect 498089 386561 498127 386595
rect 498161 386561 498199 386595
rect 498233 386561 498271 386595
rect 498305 386561 498343 386595
rect 498377 386561 498393 386595
rect 497103 386555 498393 386561
rect 496808 386507 496851 386541
rect 496885 386507 496928 386541
rect 496808 386141 496928 386507
rect 498688 386541 498808 386907
rect 498688 386507 498731 386541
rect 498765 386507 498808 386541
rect 496808 386107 496851 386141
rect 496885 386107 496928 386141
rect 496808 385741 496928 386107
rect 497103 386137 498393 386143
rect 497103 386103 497119 386137
rect 497153 386103 497191 386137
rect 497225 386103 497263 386137
rect 497297 386103 497335 386137
rect 497369 386103 497407 386137
rect 497441 386103 497479 386137
rect 497513 386103 497551 386137
rect 497585 386103 497623 386137
rect 497657 386103 497695 386137
rect 497729 386103 497767 386137
rect 497801 386103 497839 386137
rect 497873 386103 497911 386137
rect 497945 386103 497983 386137
rect 498017 386103 498055 386137
rect 498089 386103 498127 386137
rect 498161 386103 498199 386137
rect 498233 386103 498271 386137
rect 498305 386103 498343 386137
rect 498377 386103 498393 386137
rect 497103 386097 498393 386103
rect 498688 386141 498808 386507
rect 498688 386107 498731 386141
rect 498765 386107 498808 386141
rect 496808 385707 496851 385741
rect 496885 385707 496928 385741
rect 496808 385341 496928 385707
rect 498688 385741 498808 386107
rect 498688 385707 498731 385741
rect 498765 385707 498808 385741
rect 497103 385679 498393 385685
rect 497103 385645 497119 385679
rect 497153 385645 497191 385679
rect 497225 385645 497263 385679
rect 497297 385645 497335 385679
rect 497369 385645 497407 385679
rect 497441 385645 497479 385679
rect 497513 385645 497551 385679
rect 497585 385645 497623 385679
rect 497657 385645 497695 385679
rect 497729 385645 497767 385679
rect 497801 385645 497839 385679
rect 497873 385645 497911 385679
rect 497945 385645 497983 385679
rect 498017 385645 498055 385679
rect 498089 385645 498127 385679
rect 498161 385645 498199 385679
rect 498233 385645 498271 385679
rect 498305 385645 498343 385679
rect 498377 385645 498393 385679
rect 497103 385639 498393 385645
rect 498594 385500 498622 385555
rect 498582 385494 498634 385500
rect 498582 385436 498634 385442
rect 496808 385307 496851 385341
rect 496885 385307 496928 385341
rect 496808 384941 496928 385307
rect 498688 385341 498808 385707
rect 498688 385307 498731 385341
rect 498765 385307 498808 385341
rect 497103 385221 498393 385227
rect 497103 385187 497119 385221
rect 497153 385187 497191 385221
rect 497225 385187 497263 385221
rect 497297 385187 497335 385221
rect 497369 385187 497407 385221
rect 497441 385187 497479 385221
rect 497513 385187 497551 385221
rect 497585 385187 497623 385221
rect 497657 385187 497695 385221
rect 497729 385187 497767 385221
rect 497801 385187 497839 385221
rect 497873 385187 497911 385221
rect 497945 385187 497983 385221
rect 498017 385187 498055 385221
rect 498089 385187 498127 385221
rect 498161 385187 498199 385221
rect 498233 385187 498271 385221
rect 498305 385187 498343 385221
rect 498377 385187 498393 385221
rect 497103 385181 498393 385187
rect 496808 384907 496851 384941
rect 496885 384907 496928 384941
rect 496808 384541 496928 384907
rect 498688 384941 498808 385307
rect 498688 384907 498731 384941
rect 498765 384907 498808 384941
rect 497103 384763 498393 384769
rect 497103 384729 497119 384763
rect 497153 384729 497191 384763
rect 497225 384729 497263 384763
rect 497297 384729 497335 384763
rect 497369 384729 497407 384763
rect 497441 384729 497479 384763
rect 497513 384729 497551 384763
rect 497585 384729 497623 384763
rect 497657 384729 497695 384763
rect 497729 384729 497767 384763
rect 497801 384729 497839 384763
rect 497873 384729 497911 384763
rect 497945 384729 497983 384763
rect 498017 384729 498055 384763
rect 498089 384729 498127 384763
rect 498161 384729 498199 384763
rect 498233 384729 498271 384763
rect 498305 384729 498343 384763
rect 498377 384729 498393 384763
rect 497103 384723 498393 384729
rect 496808 384507 496851 384541
rect 496885 384507 496928 384541
rect 496808 384141 496928 384507
rect 498688 384541 498808 384907
rect 498688 384507 498731 384541
rect 498765 384507 498808 384541
rect 497103 384305 498393 384311
rect 497103 384271 497119 384305
rect 497153 384271 497191 384305
rect 497225 384271 497263 384305
rect 497297 384271 497335 384305
rect 497369 384271 497407 384305
rect 497441 384271 497479 384305
rect 497513 384271 497551 384305
rect 497585 384271 497623 384305
rect 497657 384271 497695 384305
rect 497729 384271 497767 384305
rect 497801 384271 497839 384305
rect 497873 384271 497911 384305
rect 497945 384271 497983 384305
rect 498017 384271 498055 384305
rect 498089 384271 498127 384305
rect 498161 384271 498199 384305
rect 498233 384271 498271 384305
rect 498305 384271 498343 384305
rect 498377 384271 498393 384305
rect 497103 384265 498393 384271
rect 496808 384107 496851 384141
rect 496885 384107 496928 384141
rect 496808 383741 496928 384107
rect 498688 384141 498808 384507
rect 498688 384107 498731 384141
rect 498765 384107 498808 384141
rect 497103 383847 498393 383853
rect 497103 383813 497119 383847
rect 497153 383813 497191 383847
rect 497225 383813 497263 383847
rect 497297 383813 497335 383847
rect 497369 383813 497407 383847
rect 497441 383813 497479 383847
rect 497513 383813 497551 383847
rect 497585 383813 497623 383847
rect 497657 383813 497695 383847
rect 497729 383813 497767 383847
rect 497801 383813 497839 383847
rect 497873 383813 497911 383847
rect 497945 383813 497983 383847
rect 498017 383813 498055 383847
rect 498089 383813 498127 383847
rect 498161 383813 498199 383847
rect 498233 383813 498271 383847
rect 498305 383813 498343 383847
rect 498377 383813 498393 383847
rect 497103 383807 498393 383813
rect 496808 383707 496851 383741
rect 496885 383707 496928 383741
rect 496808 383341 496928 383707
rect 498688 383741 498808 384107
rect 498688 383707 498731 383741
rect 498765 383707 498808 383741
rect 497103 383389 498393 383395
rect 497103 383355 497119 383389
rect 497153 383355 497191 383389
rect 497225 383355 497263 383389
rect 497297 383355 497335 383389
rect 497369 383355 497407 383389
rect 497441 383355 497479 383389
rect 497513 383355 497551 383389
rect 497585 383355 497623 383389
rect 497657 383355 497695 383389
rect 497729 383355 497767 383389
rect 497801 383355 497839 383389
rect 497873 383355 497911 383389
rect 497945 383355 497983 383389
rect 498017 383355 498055 383389
rect 498089 383355 498127 383389
rect 498161 383355 498199 383389
rect 498233 383355 498271 383389
rect 498305 383355 498343 383389
rect 498377 383355 498393 383389
rect 497103 383349 498393 383355
rect 496808 383307 496851 383341
rect 496885 383307 496928 383341
rect 496808 382941 496928 383307
rect 496808 382907 496851 382941
rect 496885 382907 496928 382941
rect 498688 383341 498808 383707
rect 498688 383307 498731 383341
rect 498765 383307 498808 383341
rect 498688 382941 498808 383307
rect 496808 382541 496928 382907
rect 497103 382931 498393 382937
rect 497103 382897 497119 382931
rect 497153 382897 497191 382931
rect 497225 382897 497263 382931
rect 497297 382897 497335 382931
rect 497369 382897 497407 382931
rect 497441 382897 497479 382931
rect 497513 382897 497551 382931
rect 497585 382897 497623 382931
rect 497657 382897 497695 382931
rect 497729 382897 497767 382931
rect 497801 382897 497839 382931
rect 497873 382897 497911 382931
rect 497945 382897 497983 382931
rect 498017 382897 498055 382931
rect 498089 382897 498127 382931
rect 498161 382897 498199 382931
rect 498233 382897 498271 382931
rect 498305 382897 498343 382931
rect 498377 382897 498393 382931
rect 497103 382891 498393 382897
rect 498688 382907 498731 382941
rect 498765 382907 498808 382941
rect 496808 382507 496851 382541
rect 496885 382507 496928 382541
rect 496808 382141 496928 382507
rect 498688 382541 498808 382907
rect 498688 382507 498731 382541
rect 498765 382507 498808 382541
rect 497103 382473 498393 382479
rect 497103 382439 497119 382473
rect 497153 382439 497191 382473
rect 497225 382439 497263 382473
rect 497297 382439 497335 382473
rect 497369 382439 497407 382473
rect 497441 382439 497479 382473
rect 497513 382439 497551 382473
rect 497585 382439 497623 382473
rect 497657 382439 497695 382473
rect 497729 382439 497767 382473
rect 497801 382439 497839 382473
rect 497873 382439 497911 382473
rect 497945 382439 497983 382473
rect 498017 382439 498055 382473
rect 498089 382439 498127 382473
rect 498161 382439 498199 382473
rect 498233 382439 498271 382473
rect 498305 382439 498343 382473
rect 498377 382439 498393 382473
rect 497103 382433 498393 382439
rect 496808 382107 496851 382141
rect 496885 382107 496928 382141
rect 496808 381741 496928 382107
rect 498688 382141 498808 382507
rect 498688 382107 498731 382141
rect 498765 382107 498808 382141
rect 497103 382015 498393 382021
rect 497103 381981 497119 382015
rect 497153 381981 497191 382015
rect 497225 381981 497263 382015
rect 497297 381981 497335 382015
rect 497369 381981 497407 382015
rect 497441 381981 497479 382015
rect 497513 381981 497551 382015
rect 497585 381981 497623 382015
rect 497657 381981 497695 382015
rect 497729 381981 497767 382015
rect 497801 381981 497839 382015
rect 497873 381981 497911 382015
rect 497945 381981 497983 382015
rect 498017 381981 498055 382015
rect 498089 381981 498127 382015
rect 498161 381981 498199 382015
rect 498233 381981 498271 382015
rect 498305 381981 498343 382015
rect 498377 381981 498393 382015
rect 497103 381975 498393 381981
rect 496808 381707 496851 381741
rect 496885 381707 496928 381741
rect 496808 381341 496928 381707
rect 498688 381741 498808 382107
rect 498688 381707 498731 381741
rect 498765 381707 498808 381741
rect 497103 381557 498393 381563
rect 497103 381523 497119 381557
rect 497153 381523 497191 381557
rect 497225 381523 497263 381557
rect 497297 381523 497335 381557
rect 497369 381523 497407 381557
rect 497441 381523 497479 381557
rect 497513 381523 497551 381557
rect 497585 381523 497623 381557
rect 497657 381523 497695 381557
rect 497729 381523 497767 381557
rect 497801 381523 497839 381557
rect 497873 381523 497911 381557
rect 497945 381523 497983 381557
rect 498017 381523 498055 381557
rect 498089 381523 498127 381557
rect 498161 381523 498199 381557
rect 498233 381523 498271 381557
rect 498305 381523 498343 381557
rect 498377 381523 498393 381557
rect 497103 381517 498393 381523
rect 496808 381307 496851 381341
rect 496885 381307 496928 381341
rect 496808 380941 496928 381307
rect 498688 381341 498808 381707
rect 498688 381307 498731 381341
rect 498765 381307 498808 381341
rect 497103 381099 498393 381105
rect 497103 381065 497119 381099
rect 497153 381065 497191 381099
rect 497225 381065 497263 381099
rect 497297 381065 497335 381099
rect 497369 381065 497407 381099
rect 497441 381065 497479 381099
rect 497513 381065 497551 381099
rect 497585 381065 497623 381099
rect 497657 381065 497695 381099
rect 497729 381065 497767 381099
rect 497801 381065 497839 381099
rect 497873 381065 497911 381099
rect 497945 381065 497983 381099
rect 498017 381065 498055 381099
rect 498089 381065 498127 381099
rect 498161 381065 498199 381099
rect 498233 381065 498271 381099
rect 498305 381065 498343 381099
rect 498377 381065 498393 381099
rect 497103 381059 498393 381065
rect 496808 380907 496851 380941
rect 496885 380907 496928 380941
rect 496808 380541 496928 380907
rect 498688 380941 498808 381307
rect 498688 380907 498731 380941
rect 498765 380907 498808 380941
rect 497103 380641 498393 380647
rect 497103 380607 497119 380641
rect 497153 380607 497191 380641
rect 497225 380607 497263 380641
rect 497297 380607 497335 380641
rect 497369 380607 497407 380641
rect 497441 380607 497479 380641
rect 497513 380607 497551 380641
rect 497585 380607 497623 380641
rect 497657 380607 497695 380641
rect 497729 380607 497767 380641
rect 497801 380607 497839 380641
rect 497873 380607 497911 380641
rect 497945 380607 497983 380641
rect 498017 380607 498055 380641
rect 498089 380607 498127 380641
rect 498161 380607 498199 380641
rect 498233 380607 498271 380641
rect 498305 380607 498343 380641
rect 498377 380607 498393 380641
rect 497103 380601 498393 380607
rect 496808 380507 496851 380541
rect 496885 380507 496928 380541
rect 496808 380141 496928 380507
rect 498688 380541 498808 380907
rect 498688 380507 498731 380541
rect 498765 380507 498808 380541
rect 497103 380183 498393 380189
rect 497103 380149 497119 380183
rect 497153 380149 497191 380183
rect 497225 380149 497263 380183
rect 497297 380149 497335 380183
rect 497369 380149 497407 380183
rect 497441 380149 497479 380183
rect 497513 380149 497551 380183
rect 497585 380149 497623 380183
rect 497657 380149 497695 380183
rect 497729 380149 497767 380183
rect 497801 380149 497839 380183
rect 497873 380149 497911 380183
rect 497945 380149 497983 380183
rect 498017 380149 498055 380183
rect 498089 380149 498127 380183
rect 498161 380149 498199 380183
rect 498233 380149 498271 380183
rect 498305 380149 498343 380183
rect 498377 380149 498393 380183
rect 497103 380143 498393 380149
rect 496808 380107 496851 380141
rect 496885 380107 496928 380141
rect 496808 379741 496928 380107
rect 496808 379707 496851 379741
rect 496885 379707 496928 379741
rect 498688 380141 498808 380507
rect 498688 380107 498731 380141
rect 498765 380107 498808 380141
rect 498688 379741 498808 380107
rect 496808 379341 496928 379707
rect 497103 379725 498393 379731
rect 497103 379691 497119 379725
rect 497153 379691 497191 379725
rect 497225 379691 497263 379725
rect 497297 379691 497335 379725
rect 497369 379691 497407 379725
rect 497441 379691 497479 379725
rect 497513 379691 497551 379725
rect 497585 379691 497623 379725
rect 497657 379691 497695 379725
rect 497729 379691 497767 379725
rect 497801 379691 497839 379725
rect 497873 379691 497911 379725
rect 497945 379691 497983 379725
rect 498017 379691 498055 379725
rect 498089 379691 498127 379725
rect 498161 379691 498199 379725
rect 498233 379691 498271 379725
rect 498305 379691 498343 379725
rect 498377 379691 498393 379725
rect 497103 379685 498393 379691
rect 498688 379707 498731 379741
rect 498765 379707 498808 379741
rect 496808 379307 496851 379341
rect 496885 379307 496928 379341
rect 496808 378941 496928 379307
rect 498688 379341 498808 379707
rect 498688 379307 498731 379341
rect 498765 379307 498808 379341
rect 497103 379267 498393 379273
rect 497103 379233 497119 379267
rect 497153 379233 497191 379267
rect 497225 379233 497263 379267
rect 497297 379233 497335 379267
rect 497369 379233 497407 379267
rect 497441 379233 497479 379267
rect 497513 379233 497551 379267
rect 497585 379233 497623 379267
rect 497657 379233 497695 379267
rect 497729 379233 497767 379267
rect 497801 379233 497839 379267
rect 497873 379233 497911 379267
rect 497945 379233 497983 379267
rect 498017 379233 498055 379267
rect 498089 379233 498127 379267
rect 498161 379233 498199 379267
rect 498233 379233 498271 379267
rect 498305 379233 498343 379267
rect 498377 379233 498393 379267
rect 497103 379227 498393 379233
rect 496808 378907 496851 378941
rect 496885 378907 496928 378941
rect 496808 378541 496928 378907
rect 498688 378941 498808 379307
rect 498688 378907 498731 378941
rect 498765 378907 498808 378941
rect 497103 378809 498393 378815
rect 497103 378775 497119 378809
rect 497153 378775 497191 378809
rect 497225 378775 497263 378809
rect 497297 378775 497335 378809
rect 497369 378775 497407 378809
rect 497441 378775 497479 378809
rect 497513 378775 497551 378809
rect 497585 378775 497623 378809
rect 497657 378775 497695 378809
rect 497729 378775 497767 378809
rect 497801 378775 497839 378809
rect 497873 378775 497911 378809
rect 497945 378775 497983 378809
rect 498017 378775 498055 378809
rect 498089 378775 498127 378809
rect 498161 378775 498199 378809
rect 498233 378775 498271 378809
rect 498305 378775 498343 378809
rect 498377 378775 498393 378809
rect 497103 378769 498393 378775
rect 496808 378507 496851 378541
rect 496885 378507 496928 378541
rect 496808 378141 496928 378507
rect 498688 378541 498808 378907
rect 498688 378507 498731 378541
rect 498765 378507 498808 378541
rect 497103 378351 498393 378357
rect 497103 378317 497119 378351
rect 497153 378317 497191 378351
rect 497225 378317 497263 378351
rect 497297 378317 497335 378351
rect 497369 378317 497407 378351
rect 497441 378317 497479 378351
rect 497513 378317 497551 378351
rect 497585 378317 497623 378351
rect 497657 378317 497695 378351
rect 497729 378317 497767 378351
rect 497801 378317 497839 378351
rect 497873 378317 497911 378351
rect 497945 378317 497983 378351
rect 498017 378317 498055 378351
rect 498089 378317 498127 378351
rect 498161 378317 498199 378351
rect 498233 378317 498271 378351
rect 498305 378317 498343 378351
rect 498377 378317 498393 378351
rect 497103 378311 498393 378317
rect 496808 378107 496851 378141
rect 496885 378107 496928 378141
rect 496808 377741 496928 378107
rect 498688 378141 498808 378507
rect 498688 378107 498731 378141
rect 498765 378107 498808 378141
rect 497103 377893 498393 377899
rect 497103 377859 497119 377893
rect 497153 377859 497191 377893
rect 497225 377859 497263 377893
rect 497297 377859 497335 377893
rect 497369 377859 497407 377893
rect 497441 377859 497479 377893
rect 497513 377859 497551 377893
rect 497585 377859 497623 377893
rect 497657 377859 497695 377893
rect 497729 377859 497767 377893
rect 497801 377859 497839 377893
rect 497873 377859 497911 377893
rect 497945 377859 497983 377893
rect 498017 377859 498055 377893
rect 498089 377859 498127 377893
rect 498161 377859 498199 377893
rect 498233 377859 498271 377893
rect 498305 377859 498343 377893
rect 498377 377859 498393 377893
rect 497103 377853 498393 377859
rect 496808 377707 496851 377741
rect 496885 377707 496928 377741
rect 496808 377341 496928 377707
rect 498688 377741 498808 378107
rect 498688 377707 498731 377741
rect 498765 377707 498808 377741
rect 497103 377435 498393 377441
rect 497103 377401 497119 377435
rect 497153 377401 497191 377435
rect 497225 377401 497263 377435
rect 497297 377401 497335 377435
rect 497369 377401 497407 377435
rect 497441 377401 497479 377435
rect 497513 377401 497551 377435
rect 497585 377401 497623 377435
rect 497657 377401 497695 377435
rect 497729 377401 497767 377435
rect 497801 377401 497839 377435
rect 497873 377401 497911 377435
rect 497945 377401 497983 377435
rect 498017 377401 498055 377435
rect 498089 377401 498127 377435
rect 498161 377401 498199 377435
rect 498233 377401 498271 377435
rect 498305 377401 498343 377435
rect 498377 377401 498393 377435
rect 497103 377395 498393 377401
rect 496808 377307 496851 377341
rect 496885 377307 496928 377341
rect 496808 376941 496928 377307
rect 498688 377341 498808 377707
rect 498688 377307 498731 377341
rect 498765 377307 498808 377341
rect 496808 376907 496851 376941
rect 496885 376907 496928 376941
rect 497103 376977 498393 376983
rect 497103 376943 497119 376977
rect 497153 376943 497191 376977
rect 497225 376943 497263 376977
rect 497297 376943 497335 376977
rect 497369 376943 497407 376977
rect 497441 376943 497479 376977
rect 497513 376943 497551 376977
rect 497585 376943 497623 376977
rect 497657 376943 497695 376977
rect 497729 376943 497767 376977
rect 497801 376943 497839 376977
rect 497873 376943 497911 376977
rect 497945 376943 497983 376977
rect 498017 376943 498055 376977
rect 498089 376943 498127 376977
rect 498161 376943 498199 376977
rect 498233 376943 498271 376977
rect 498305 376943 498343 376977
rect 498377 376943 498393 376977
rect 497103 376937 498393 376943
rect 498688 376941 498808 377307
rect 496808 376541 496928 376907
rect 496808 376507 496851 376541
rect 496885 376507 496928 376541
rect 498688 376907 498731 376941
rect 498765 376907 498808 376941
rect 498688 376541 498808 376907
rect 496808 376141 496928 376507
rect 497103 376519 498393 376525
rect 497103 376485 497119 376519
rect 497153 376485 497191 376519
rect 497225 376485 497263 376519
rect 497297 376485 497335 376519
rect 497369 376485 497407 376519
rect 497441 376485 497479 376519
rect 497513 376485 497551 376519
rect 497585 376485 497623 376519
rect 497657 376485 497695 376519
rect 497729 376485 497767 376519
rect 497801 376485 497839 376519
rect 497873 376485 497911 376519
rect 497945 376485 497983 376519
rect 498017 376485 498055 376519
rect 498089 376485 498127 376519
rect 498161 376485 498199 376519
rect 498233 376485 498271 376519
rect 498305 376485 498343 376519
rect 498377 376485 498393 376519
rect 497103 376479 498393 376485
rect 498688 376507 498731 376541
rect 498765 376507 498808 376541
rect 496808 376107 496851 376141
rect 496885 376107 496928 376141
rect 496808 375741 496928 376107
rect 498688 376141 498808 376507
rect 498688 376107 498731 376141
rect 498765 376107 498808 376141
rect 497103 376061 498393 376067
rect 497103 376027 497119 376061
rect 497153 376027 497191 376061
rect 497225 376027 497263 376061
rect 497297 376027 497335 376061
rect 497369 376027 497407 376061
rect 497441 376027 497479 376061
rect 497513 376027 497551 376061
rect 497585 376027 497623 376061
rect 497657 376027 497695 376061
rect 497729 376027 497767 376061
rect 497801 376027 497839 376061
rect 497873 376027 497911 376061
rect 497945 376027 497983 376061
rect 498017 376027 498055 376061
rect 498089 376027 498127 376061
rect 498161 376027 498199 376061
rect 498233 376027 498271 376061
rect 498305 376027 498343 376061
rect 498377 376027 498393 376061
rect 497103 376021 498393 376027
rect 496808 375707 496851 375741
rect 496885 375707 496928 375741
rect 496808 375341 496928 375707
rect 498688 375741 498808 376107
rect 498688 375707 498731 375741
rect 498765 375707 498808 375741
rect 497103 375603 498393 375609
rect 497103 375569 497119 375603
rect 497153 375569 497191 375603
rect 497225 375569 497263 375603
rect 497297 375569 497335 375603
rect 497369 375569 497407 375603
rect 497441 375569 497479 375603
rect 497513 375569 497551 375603
rect 497585 375569 497623 375603
rect 497657 375569 497695 375603
rect 497729 375569 497767 375603
rect 497801 375569 497839 375603
rect 497873 375569 497911 375603
rect 497945 375569 497983 375603
rect 498017 375569 498055 375603
rect 498089 375569 498127 375603
rect 498161 375569 498199 375603
rect 498233 375569 498271 375603
rect 498305 375569 498343 375603
rect 498377 375569 498393 375603
rect 497103 375563 498393 375569
rect 496808 375307 496851 375341
rect 496885 375307 496928 375341
rect 496808 374941 496928 375307
rect 498688 375341 498808 375707
rect 498688 375307 498731 375341
rect 498765 375307 498808 375341
rect 497103 375145 498393 375151
rect 497103 375111 497119 375145
rect 497153 375111 497191 375145
rect 497225 375111 497263 375145
rect 497297 375111 497335 375145
rect 497369 375111 497407 375145
rect 497441 375111 497479 375145
rect 497513 375111 497551 375145
rect 497585 375111 497623 375145
rect 497657 375111 497695 375145
rect 497729 375111 497767 375145
rect 497801 375111 497839 375145
rect 497873 375111 497911 375145
rect 497945 375111 497983 375145
rect 498017 375111 498055 375145
rect 498089 375111 498127 375145
rect 498161 375111 498199 375145
rect 498233 375111 498271 375145
rect 498305 375111 498343 375145
rect 498377 375111 498393 375145
rect 497103 375105 498393 375111
rect 496808 374907 496851 374941
rect 496885 374907 496928 374941
rect 496808 374541 496928 374907
rect 498688 374941 498808 375307
rect 498688 374907 498731 374941
rect 498765 374907 498808 374941
rect 497103 374687 498393 374693
rect 497103 374653 497119 374687
rect 497153 374653 497191 374687
rect 497225 374653 497263 374687
rect 497297 374653 497335 374687
rect 497369 374653 497407 374687
rect 497441 374653 497479 374687
rect 497513 374653 497551 374687
rect 497585 374653 497623 374687
rect 497657 374653 497695 374687
rect 497729 374653 497767 374687
rect 497801 374653 497839 374687
rect 497873 374653 497911 374687
rect 497945 374653 497983 374687
rect 498017 374653 498055 374687
rect 498089 374653 498127 374687
rect 498161 374653 498199 374687
rect 498233 374653 498271 374687
rect 498305 374653 498343 374687
rect 498377 374653 498393 374687
rect 497103 374647 498393 374653
rect 496808 374507 496851 374541
rect 496885 374507 496928 374541
rect 496808 374141 496928 374507
rect 498688 374541 498808 374907
rect 498688 374507 498731 374541
rect 498765 374507 498808 374541
rect 497103 374229 498393 374235
rect 497103 374195 497119 374229
rect 497153 374195 497191 374229
rect 497225 374195 497263 374229
rect 497297 374195 497335 374229
rect 497369 374195 497407 374229
rect 497441 374195 497479 374229
rect 497513 374195 497551 374229
rect 497585 374195 497623 374229
rect 497657 374195 497695 374229
rect 497729 374195 497767 374229
rect 497801 374195 497839 374229
rect 497873 374195 497911 374229
rect 497945 374195 497983 374229
rect 498017 374195 498055 374229
rect 498089 374195 498127 374229
rect 498161 374195 498199 374229
rect 498233 374195 498271 374229
rect 498305 374195 498343 374229
rect 498377 374195 498393 374229
rect 497103 374189 498393 374195
rect 496808 374107 496851 374141
rect 496885 374107 496928 374141
rect 496808 373741 496928 374107
rect 498688 374141 498808 374507
rect 498688 374107 498731 374141
rect 498765 374107 498808 374141
rect 496808 373707 496851 373741
rect 496885 373707 496928 373741
rect 497103 373771 498393 373777
rect 497103 373737 497119 373771
rect 497153 373737 497191 373771
rect 497225 373737 497263 373771
rect 497297 373737 497335 373771
rect 497369 373737 497407 373771
rect 497441 373737 497479 373771
rect 497513 373737 497551 373771
rect 497585 373737 497623 373771
rect 497657 373737 497695 373771
rect 497729 373737 497767 373771
rect 497801 373737 497839 373771
rect 497873 373737 497911 373771
rect 497945 373737 497983 373771
rect 498017 373737 498055 373771
rect 498089 373737 498127 373771
rect 498161 373737 498199 373771
rect 498233 373737 498271 373771
rect 498305 373737 498343 373771
rect 498377 373737 498393 373771
rect 497103 373731 498393 373737
rect 498688 373741 498808 374107
rect 496808 373341 496928 373707
rect 496808 373307 496851 373341
rect 496885 373307 496928 373341
rect 498688 373707 498731 373741
rect 498765 373707 498808 373741
rect 498688 373341 498808 373707
rect 496808 372941 496928 373307
rect 497103 373313 498393 373319
rect 497103 373279 497119 373313
rect 497153 373279 497191 373313
rect 497225 373279 497263 373313
rect 497297 373279 497335 373313
rect 497369 373279 497407 373313
rect 497441 373279 497479 373313
rect 497513 373279 497551 373313
rect 497585 373279 497623 373313
rect 497657 373279 497695 373313
rect 497729 373279 497767 373313
rect 497801 373279 497839 373313
rect 497873 373279 497911 373313
rect 497945 373279 497983 373313
rect 498017 373279 498055 373313
rect 498089 373279 498127 373313
rect 498161 373279 498199 373313
rect 498233 373279 498271 373313
rect 498305 373279 498343 373313
rect 498377 373279 498393 373313
rect 497103 373273 498393 373279
rect 498688 373307 498731 373341
rect 498765 373307 498808 373341
rect 496808 372907 496851 372941
rect 496885 372907 496928 372941
rect 496808 372541 496928 372907
rect 498688 372941 498808 373307
rect 498688 372907 498731 372941
rect 498765 372907 498808 372941
rect 497103 372855 498393 372861
rect 497103 372821 497119 372855
rect 497153 372821 497191 372855
rect 497225 372821 497263 372855
rect 497297 372821 497335 372855
rect 497369 372821 497407 372855
rect 497441 372821 497479 372855
rect 497513 372821 497551 372855
rect 497585 372821 497623 372855
rect 497657 372821 497695 372855
rect 497729 372821 497767 372855
rect 497801 372821 497839 372855
rect 497873 372821 497911 372855
rect 497945 372821 497983 372855
rect 498017 372821 498055 372855
rect 498089 372821 498127 372855
rect 498161 372821 498199 372855
rect 498233 372821 498271 372855
rect 498305 372821 498343 372855
rect 498377 372821 498393 372855
rect 497103 372815 498393 372821
rect 496808 372507 496851 372541
rect 496885 372507 496928 372541
rect 496808 371811 496928 372507
rect 498688 372541 498808 372907
rect 498688 372507 498731 372541
rect 498765 372507 498808 372541
rect 497103 372397 498393 372403
rect 497103 372363 497119 372397
rect 497153 372363 497191 372397
rect 497225 372363 497263 372397
rect 497297 372363 497335 372397
rect 497369 372363 497407 372397
rect 497441 372363 497479 372397
rect 497513 372363 497551 372397
rect 497585 372363 497623 372397
rect 497657 372363 497695 372397
rect 497729 372363 497767 372397
rect 497801 372363 497839 372397
rect 497873 372363 497911 372397
rect 497945 372363 497983 372397
rect 498017 372363 498055 372397
rect 498089 372363 498127 372397
rect 498161 372363 498199 372397
rect 498233 372363 498271 372397
rect 498305 372363 498343 372397
rect 498377 372363 498393 372397
rect 497103 372357 498393 372363
rect 496808 371777 496851 371811
rect 496885 371777 496928 371811
rect 496808 371611 496928 371777
rect 496808 371577 496851 371611
rect 496885 371577 496928 371611
rect 496808 371411 496928 371577
rect 496808 371377 496851 371411
rect 496885 371377 496928 371411
rect 496808 371211 496928 371377
rect 496808 371177 496851 371211
rect 496885 371177 496928 371211
rect 496808 371011 496928 371177
rect 496808 370977 496851 371011
rect 496885 370977 496928 371011
rect 496808 370811 496928 370977
rect 496808 370777 496851 370811
rect 496885 370777 496928 370811
rect 496808 370611 496928 370777
rect 496808 370577 496851 370611
rect 496885 370577 496928 370611
rect 496808 370411 496928 370577
rect 496808 370377 496851 370411
rect 496885 370377 496928 370411
rect 496808 370211 496928 370377
rect 496808 370177 496851 370211
rect 496885 370177 496928 370211
rect 496808 370011 496928 370177
rect 496808 369977 496851 370011
rect 496885 369977 496928 370011
rect 496808 369811 496928 369977
rect 496808 369777 496851 369811
rect 496885 369777 496928 369811
rect 496808 369611 496928 369777
rect 496808 369577 496851 369611
rect 496885 369577 496928 369611
rect 496808 369411 496928 369577
rect 496808 369377 496851 369411
rect 496885 369377 496928 369411
rect 496808 369211 496928 369377
rect 496808 369177 496851 369211
rect 496885 369177 496928 369211
rect 496808 369011 496928 369177
rect 496808 368977 496851 369011
rect 496885 368977 496928 369011
rect 496808 368811 496928 368977
rect 496808 368777 496851 368811
rect 496885 368777 496928 368811
rect 496808 368611 496928 368777
rect 496808 368577 496851 368611
rect 496885 368577 496928 368611
rect 496808 368411 496928 368577
rect 496808 368377 496851 368411
rect 496885 368377 496928 368411
rect 496808 368211 496928 368377
rect 496808 368177 496851 368211
rect 496885 368177 496928 368211
rect 496808 368011 496928 368177
rect 496808 367977 496851 368011
rect 496885 367977 496928 368011
rect 496808 367811 496928 367977
rect 496808 367777 496851 367811
rect 496885 367777 496928 367811
rect 496808 367611 496928 367777
rect 496808 367577 496851 367611
rect 496885 367577 496928 367611
rect 496808 367411 496928 367577
rect 496808 367377 496851 367411
rect 496885 367377 496928 367411
rect 496808 367211 496928 367377
rect 496808 367177 496851 367211
rect 496885 367177 496928 367211
rect 496808 367011 496928 367177
rect 496808 366977 496851 367011
rect 496885 366977 496928 367011
rect 496808 366811 496928 366977
rect 496808 366777 496851 366811
rect 496885 366777 496928 366811
rect 496808 366611 496928 366777
rect 496808 366577 496851 366611
rect 496885 366577 496928 366611
rect 496808 366411 496928 366577
rect 496808 366377 496851 366411
rect 496885 366377 496928 366411
rect 496808 366211 496928 366377
rect 496808 366177 496851 366211
rect 496885 366177 496928 366211
rect 496808 366011 496928 366177
rect 496808 365977 496851 366011
rect 496885 365977 496928 366011
rect 496808 365811 496928 365977
rect 496808 365777 496851 365811
rect 496885 365777 496928 365811
rect 496808 365611 496928 365777
rect 496808 365577 496851 365611
rect 496885 365577 496928 365611
rect 496808 365411 496928 365577
rect 496808 365377 496851 365411
rect 496885 365377 496928 365411
rect 496808 365211 496928 365377
rect 496808 365177 496851 365211
rect 496885 365177 496928 365211
rect 496808 365011 496928 365177
rect 496808 364977 496851 365011
rect 496885 364977 496928 365011
rect 496808 364811 496928 364977
rect 496808 364777 496851 364811
rect 496885 364777 496928 364811
rect 496808 364611 496928 364777
rect 496808 364577 496851 364611
rect 496885 364577 496928 364611
rect 496808 364411 496928 364577
rect 496808 364377 496851 364411
rect 496885 364377 496928 364411
rect 496808 364211 496928 364377
rect 496808 364177 496851 364211
rect 496885 364177 496928 364211
rect 496808 364011 496928 364177
rect 496808 363977 496851 364011
rect 496885 363977 496928 364011
rect 496808 363811 496928 363977
rect 496808 363777 496851 363811
rect 496885 363777 496928 363811
rect 496808 363611 496928 363777
rect 496808 363577 496851 363611
rect 496885 363577 496928 363611
rect 496808 363411 496928 363577
rect 496808 363377 496851 363411
rect 496885 363377 496928 363411
rect 496808 363211 496928 363377
rect 496808 363177 496851 363211
rect 496885 363177 496928 363211
rect 496808 363011 496928 363177
rect 496808 362977 496851 363011
rect 496885 362977 496928 363011
rect 496808 362811 496928 362977
rect 496808 362777 496851 362811
rect 496885 362777 496928 362811
rect 496808 361476 496928 362777
rect 497178 371948 497248 371968
rect 497178 371914 497184 371948
rect 497218 371914 497248 371948
rect 497178 371858 497248 371914
rect 497178 371824 497184 371858
rect 497218 371824 497248 371858
rect 497178 371768 497248 371824
rect 498688 371811 498808 372507
rect 497178 371734 497184 371768
rect 497218 371734 497248 371768
rect 497178 371682 497248 371734
rect 497328 371784 497398 371804
rect 497328 371750 497344 371784
rect 497378 371750 497398 371784
rect 497328 371700 497398 371750
rect 497324 371694 497398 371700
rect 497178 371678 497324 371682
rect 497178 371644 497184 371678
rect 497218 371654 497324 371678
rect 497378 371660 497398 371694
rect 497218 371644 497248 371654
rect 497178 371588 497248 371644
rect 497376 371642 497398 371660
rect 497324 371636 497398 371642
rect 497178 371554 497184 371588
rect 497218 371554 497248 371588
rect 497178 371498 497248 371554
rect 497178 371464 497184 371498
rect 497218 371464 497248 371498
rect 497178 371408 497248 371464
rect 497178 371374 497184 371408
rect 497218 371374 497248 371408
rect 497178 371318 497248 371374
rect 497178 371284 497184 371318
rect 497218 371284 497248 371318
rect 497178 371228 497248 371284
rect 497178 371194 497184 371228
rect 497218 371194 497248 371228
rect 497178 371138 497248 371194
rect 497178 371104 497184 371138
rect 497218 371104 497248 371138
rect 497178 371048 497248 371104
rect 497178 371014 497184 371048
rect 497218 371014 497248 371048
rect 497178 370958 497248 371014
rect 497178 370924 497184 370958
rect 497218 370924 497248 370958
rect 497178 370868 497248 370924
rect 497178 370834 497184 370868
rect 497218 370834 497248 370868
rect 497178 370778 497248 370834
rect 497178 370744 497184 370778
rect 497218 370744 497248 370778
rect 497178 370608 497248 370744
rect 497178 370574 497184 370608
rect 497218 370574 497248 370608
rect 497178 370518 497248 370574
rect 497178 370484 497184 370518
rect 497218 370484 497248 370518
rect 497178 370428 497248 370484
rect 497178 370394 497184 370428
rect 497218 370394 497248 370428
rect 497178 370338 497248 370394
rect 497178 370304 497184 370338
rect 497218 370304 497248 370338
rect 497178 370248 497248 370304
rect 497178 370214 497184 370248
rect 497218 370214 497248 370248
rect 497178 370158 497248 370214
rect 497178 370124 497184 370158
rect 497218 370124 497248 370158
rect 497178 370068 497248 370124
rect 497178 370034 497184 370068
rect 497218 370034 497248 370068
rect 497178 369978 497248 370034
rect 497178 369944 497184 369978
rect 497218 369944 497248 369978
rect 497178 369888 497248 369944
rect 497178 369854 497184 369888
rect 497218 369854 497248 369888
rect 497178 369798 497248 369854
rect 497178 369764 497184 369798
rect 497218 369764 497248 369798
rect 497178 369708 497248 369764
rect 497178 369674 497184 369708
rect 497218 369674 497248 369708
rect 497178 369618 497248 369674
rect 497178 369584 497184 369618
rect 497218 369584 497248 369618
rect 497178 369528 497248 369584
rect 497178 369494 497184 369528
rect 497218 369494 497248 369528
rect 497178 369438 497248 369494
rect 497178 369404 497184 369438
rect 497218 369404 497248 369438
rect 497178 369268 497248 369404
rect 497178 369234 497184 369268
rect 497218 369234 497248 369268
rect 497178 369178 497248 369234
rect 497178 369144 497184 369178
rect 497218 369144 497248 369178
rect 497178 369088 497248 369144
rect 497178 369054 497184 369088
rect 497218 369054 497248 369088
rect 497178 368998 497248 369054
rect 497178 368964 497184 368998
rect 497218 368964 497248 368998
rect 497178 368908 497248 368964
rect 497178 368874 497184 368908
rect 497218 368874 497248 368908
rect 497178 368818 497248 368874
rect 497178 368784 497184 368818
rect 497218 368784 497248 368818
rect 497178 368728 497248 368784
rect 497178 368694 497184 368728
rect 497218 368694 497248 368728
rect 497178 368638 497248 368694
rect 497178 368604 497184 368638
rect 497218 368604 497248 368638
rect 497178 368548 497248 368604
rect 497178 368514 497184 368548
rect 497218 368514 497248 368548
rect 497178 368458 497248 368514
rect 497178 368424 497184 368458
rect 497218 368424 497248 368458
rect 497178 368368 497248 368424
rect 497178 368334 497184 368368
rect 497218 368334 497248 368368
rect 497178 368278 497248 368334
rect 497178 368244 497184 368278
rect 497218 368244 497248 368278
rect 497178 368188 497248 368244
rect 497178 368154 497184 368188
rect 497218 368154 497248 368188
rect 497178 368098 497248 368154
rect 497178 368064 497184 368098
rect 497218 368064 497248 368098
rect 497178 367928 497248 368064
rect 497178 367894 497184 367928
rect 497218 367894 497248 367928
rect 497178 367838 497248 367894
rect 497178 367804 497184 367838
rect 497218 367804 497248 367838
rect 497178 367748 497248 367804
rect 497178 367714 497184 367748
rect 497218 367714 497248 367748
rect 497178 367658 497248 367714
rect 497178 367624 497184 367658
rect 497218 367624 497248 367658
rect 497178 367568 497248 367624
rect 497178 367534 497184 367568
rect 497218 367534 497248 367568
rect 497178 367478 497248 367534
rect 497178 367444 497184 367478
rect 497218 367444 497248 367478
rect 497178 367388 497248 367444
rect 497178 367354 497184 367388
rect 497218 367354 497248 367388
rect 497178 367298 497248 367354
rect 497178 367264 497184 367298
rect 497218 367264 497248 367298
rect 497178 367208 497248 367264
rect 497178 367174 497184 367208
rect 497218 367174 497248 367208
rect 497178 367118 497248 367174
rect 497178 367084 497184 367118
rect 497218 367084 497248 367118
rect 497178 367028 497248 367084
rect 497178 366994 497184 367028
rect 497218 366994 497248 367028
rect 497178 366938 497248 366994
rect 497178 366904 497184 366938
rect 497218 366904 497248 366938
rect 497178 366848 497248 366904
rect 497178 366814 497184 366848
rect 497218 366814 497248 366848
rect 497178 366758 497248 366814
rect 497178 366724 497184 366758
rect 497218 366724 497248 366758
rect 497178 366588 497248 366724
rect 497178 366554 497184 366588
rect 497218 366554 497248 366588
rect 497178 366498 497248 366554
rect 497178 366464 497184 366498
rect 497218 366464 497248 366498
rect 497178 366408 497248 366464
rect 497178 366374 497184 366408
rect 497218 366374 497248 366408
rect 497178 366318 497248 366374
rect 497178 366284 497184 366318
rect 497218 366284 497248 366318
rect 497178 366228 497248 366284
rect 497178 366194 497184 366228
rect 497218 366194 497248 366228
rect 497178 366138 497248 366194
rect 497178 366104 497184 366138
rect 497218 366104 497248 366138
rect 497178 366048 497248 366104
rect 497178 366014 497184 366048
rect 497218 366014 497248 366048
rect 497178 365958 497248 366014
rect 497178 365924 497184 365958
rect 497218 365924 497248 365958
rect 497178 365868 497248 365924
rect 497178 365834 497184 365868
rect 497218 365834 497248 365868
rect 497178 365778 497248 365834
rect 497178 365744 497184 365778
rect 497218 365744 497248 365778
rect 497178 365688 497248 365744
rect 497178 365654 497184 365688
rect 497218 365654 497248 365688
rect 497178 365598 497248 365654
rect 497178 365564 497184 365598
rect 497218 365564 497248 365598
rect 497178 365508 497248 365564
rect 497178 365474 497184 365508
rect 497218 365474 497248 365508
rect 497178 365418 497248 365474
rect 497178 365384 497184 365418
rect 497218 365384 497248 365418
rect 497178 365248 497248 365384
rect 497178 365214 497184 365248
rect 497218 365214 497248 365248
rect 497178 365158 497248 365214
rect 497178 365124 497184 365158
rect 497218 365124 497248 365158
rect 497178 365068 497248 365124
rect 497178 365034 497184 365068
rect 497218 365034 497248 365068
rect 497178 364978 497248 365034
rect 497178 364944 497184 364978
rect 497218 364944 497248 364978
rect 497178 364888 497248 364944
rect 497178 364854 497184 364888
rect 497218 364854 497248 364888
rect 497178 364798 497248 364854
rect 497178 364764 497184 364798
rect 497218 364764 497248 364798
rect 497178 364708 497248 364764
rect 497178 364674 497184 364708
rect 497218 364674 497248 364708
rect 497178 364618 497248 364674
rect 497178 364584 497184 364618
rect 497218 364584 497248 364618
rect 497178 364528 497248 364584
rect 497178 364494 497184 364528
rect 497218 364494 497248 364528
rect 497178 364438 497248 364494
rect 497178 364404 497184 364438
rect 497218 364404 497248 364438
rect 497178 364348 497248 364404
rect 497178 364314 497184 364348
rect 497218 364314 497248 364348
rect 497178 364258 497248 364314
rect 497178 364224 497184 364258
rect 497218 364224 497248 364258
rect 497178 364168 497248 364224
rect 497178 364134 497184 364168
rect 497218 364134 497248 364168
rect 497178 364078 497248 364134
rect 497178 364044 497184 364078
rect 497218 364044 497248 364078
rect 497178 363908 497248 364044
rect 497178 363874 497184 363908
rect 497218 363874 497248 363908
rect 497178 363818 497248 363874
rect 497178 363784 497184 363818
rect 497218 363784 497248 363818
rect 497178 363728 497248 363784
rect 497178 363694 497184 363728
rect 497218 363694 497248 363728
rect 497178 363638 497248 363694
rect 497178 363604 497184 363638
rect 497218 363604 497248 363638
rect 497178 363548 497248 363604
rect 497178 363514 497184 363548
rect 497218 363514 497248 363548
rect 497178 363458 497248 363514
rect 497178 363424 497184 363458
rect 497218 363424 497248 363458
rect 497178 363368 497248 363424
rect 497178 363334 497184 363368
rect 497218 363334 497248 363368
rect 497178 363278 497248 363334
rect 497178 363244 497184 363278
rect 497218 363244 497248 363278
rect 497178 363188 497248 363244
rect 497178 363154 497184 363188
rect 497218 363154 497248 363188
rect 497178 363098 497248 363154
rect 497178 363064 497184 363098
rect 497218 363064 497248 363098
rect 497178 363008 497248 363064
rect 497178 362974 497184 363008
rect 497218 362974 497248 363008
rect 497178 362918 497248 362974
rect 497178 362884 497184 362918
rect 497218 362884 497248 362918
rect 497178 362828 497248 362884
rect 497178 362794 497184 362828
rect 497218 362794 497248 362828
rect 497328 371604 497398 371636
rect 498688 371777 498731 371811
rect 498765 371777 498808 371811
rect 498688 371694 498808 371777
rect 498688 371642 498752 371694
rect 498804 371642 498808 371694
rect 497328 371570 497344 371604
rect 497378 371570 497398 371604
rect 497328 371514 497398 371570
rect 497328 371480 497344 371514
rect 497378 371480 497398 371514
rect 497328 371424 497398 371480
rect 497328 371390 497344 371424
rect 497378 371390 497398 371424
rect 497328 371334 497398 371390
rect 497328 371300 497344 371334
rect 497378 371300 497398 371334
rect 497328 371244 497398 371300
rect 497328 371210 497344 371244
rect 497378 371210 497398 371244
rect 497328 371154 497398 371210
rect 497328 371120 497344 371154
rect 497378 371120 497398 371154
rect 497328 371064 497398 371120
rect 497328 371030 497344 371064
rect 497378 371030 497398 371064
rect 497328 370974 497398 371030
rect 497328 370940 497344 370974
rect 497378 370940 497398 370974
rect 497328 370884 497398 370940
rect 497328 370850 497344 370884
rect 497378 370850 497398 370884
rect 497328 370444 497398 370850
rect 497328 370410 497344 370444
rect 497378 370410 497398 370444
rect 497328 370354 497398 370410
rect 497328 370320 497344 370354
rect 497378 370320 497398 370354
rect 497328 370264 497398 370320
rect 497328 370230 497344 370264
rect 497378 370230 497398 370264
rect 497328 370174 497398 370230
rect 497328 370140 497344 370174
rect 497378 370140 497398 370174
rect 497328 370084 497398 370140
rect 497328 370050 497344 370084
rect 497378 370050 497398 370084
rect 497328 369994 497398 370050
rect 497328 369960 497344 369994
rect 497378 369960 497398 369994
rect 497328 369904 497398 369960
rect 497328 369870 497344 369904
rect 497378 369870 497398 369904
rect 497328 369814 497398 369870
rect 497328 369780 497344 369814
rect 497378 369780 497398 369814
rect 497328 369724 497398 369780
rect 497328 369690 497344 369724
rect 497378 369690 497398 369724
rect 497328 369634 497398 369690
rect 497328 369600 497344 369634
rect 497378 369600 497398 369634
rect 497328 369544 497398 369600
rect 497328 369510 497344 369544
rect 497378 369510 497398 369544
rect 497328 369104 497398 369510
rect 497328 369070 497344 369104
rect 497378 369070 497398 369104
rect 497328 369014 497398 369070
rect 497328 368980 497344 369014
rect 497378 368980 497398 369014
rect 497328 368924 497398 368980
rect 497328 368890 497344 368924
rect 497378 368890 497398 368924
rect 497328 368834 497398 368890
rect 497328 368800 497344 368834
rect 497378 368800 497398 368834
rect 497328 368744 497398 368800
rect 497328 368710 497344 368744
rect 497378 368710 497398 368744
rect 497328 368654 497398 368710
rect 497328 368620 497344 368654
rect 497378 368620 497398 368654
rect 497328 368564 497398 368620
rect 497328 368530 497344 368564
rect 497378 368530 497398 368564
rect 497328 368474 497398 368530
rect 497328 368440 497344 368474
rect 497378 368440 497398 368474
rect 497328 368384 497398 368440
rect 497328 368350 497344 368384
rect 497378 368350 497398 368384
rect 497328 368294 497398 368350
rect 497328 368260 497344 368294
rect 497378 368260 497398 368294
rect 497328 368204 497398 368260
rect 497328 368170 497344 368204
rect 497378 368170 497398 368204
rect 497328 367764 497398 368170
rect 497328 367730 497344 367764
rect 497378 367730 497398 367764
rect 497328 367674 497398 367730
rect 497328 367640 497344 367674
rect 497378 367640 497398 367674
rect 497328 367584 497398 367640
rect 497328 367550 497344 367584
rect 497378 367550 497398 367584
rect 497328 367494 497398 367550
rect 497328 367460 497344 367494
rect 497378 367460 497398 367494
rect 497328 367404 497398 367460
rect 497328 367370 497344 367404
rect 497378 367370 497398 367404
rect 497328 367314 497398 367370
rect 497328 367280 497344 367314
rect 497378 367280 497398 367314
rect 497328 367224 497398 367280
rect 497328 367190 497344 367224
rect 497378 367190 497398 367224
rect 497328 367134 497398 367190
rect 497328 367100 497344 367134
rect 497378 367100 497398 367134
rect 497328 367044 497398 367100
rect 497328 367010 497344 367044
rect 497378 367010 497398 367044
rect 497328 366954 497398 367010
rect 497328 366920 497344 366954
rect 497378 366920 497398 366954
rect 497328 366864 497398 366920
rect 497328 366830 497344 366864
rect 497378 366830 497398 366864
rect 497328 366424 497398 366830
rect 497328 366390 497344 366424
rect 497378 366390 497398 366424
rect 497328 366334 497398 366390
rect 497328 366300 497344 366334
rect 497378 366300 497398 366334
rect 497328 366244 497398 366300
rect 497328 366210 497344 366244
rect 497378 366210 497398 366244
rect 497328 366154 497398 366210
rect 497328 366120 497344 366154
rect 497378 366120 497398 366154
rect 497328 366064 497398 366120
rect 497328 366030 497344 366064
rect 497378 366030 497398 366064
rect 497328 365974 497398 366030
rect 497328 365940 497344 365974
rect 497378 365940 497398 365974
rect 497328 365884 497398 365940
rect 497328 365850 497344 365884
rect 497378 365850 497398 365884
rect 497328 365794 497398 365850
rect 497328 365760 497344 365794
rect 497378 365760 497398 365794
rect 497328 365704 497398 365760
rect 497328 365670 497344 365704
rect 497378 365670 497398 365704
rect 497328 365614 497398 365670
rect 497328 365580 497344 365614
rect 497378 365580 497398 365614
rect 497328 365524 497398 365580
rect 497328 365490 497344 365524
rect 497378 365490 497398 365524
rect 497328 365084 497398 365490
rect 497328 365050 497344 365084
rect 497378 365050 497398 365084
rect 497328 364994 497398 365050
rect 497328 364960 497344 364994
rect 497378 364960 497398 364994
rect 497328 364904 497398 364960
rect 497328 364870 497344 364904
rect 497378 364870 497398 364904
rect 497328 364814 497398 364870
rect 497328 364780 497344 364814
rect 497378 364780 497398 364814
rect 497328 364724 497398 364780
rect 497328 364690 497344 364724
rect 497378 364690 497398 364724
rect 497328 364634 497398 364690
rect 497328 364600 497344 364634
rect 497378 364600 497398 364634
rect 497328 364544 497398 364600
rect 497328 364510 497344 364544
rect 497378 364510 497398 364544
rect 497328 364454 497398 364510
rect 497328 364420 497344 364454
rect 497378 364420 497398 364454
rect 497328 364364 497398 364420
rect 497328 364330 497344 364364
rect 497378 364330 497398 364364
rect 497328 364274 497398 364330
rect 497328 364240 497344 364274
rect 497378 364240 497398 364274
rect 497328 364184 497398 364240
rect 497328 364150 497344 364184
rect 497378 364150 497398 364184
rect 497328 363744 497398 364150
rect 497328 363710 497344 363744
rect 497378 363710 497398 363744
rect 497328 363654 497398 363710
rect 497328 363620 497344 363654
rect 497378 363620 497398 363654
rect 497328 363564 497398 363620
rect 497328 363530 497344 363564
rect 497378 363530 497398 363564
rect 497328 363474 497398 363530
rect 497328 363440 497344 363474
rect 497378 363440 497398 363474
rect 497328 363384 497398 363440
rect 497328 363350 497344 363384
rect 497378 363350 497398 363384
rect 497328 363294 497398 363350
rect 497328 363260 497344 363294
rect 497378 363260 497398 363294
rect 497328 363204 497398 363260
rect 497328 363170 497344 363204
rect 497378 363170 497398 363204
rect 497328 363114 497398 363170
rect 497328 363080 497344 363114
rect 497378 363080 497398 363114
rect 497328 363024 497398 363080
rect 497328 362990 497344 363024
rect 497378 362990 497398 363024
rect 497328 362934 497398 362990
rect 497502 371598 498114 371630
rect 497502 371564 497548 371598
rect 497582 371564 497648 371598
rect 497682 371564 497748 371598
rect 497782 371564 497848 371598
rect 497882 371564 497948 371598
rect 497982 371564 498048 371598
rect 498082 371564 498114 371598
rect 497502 371498 498114 371564
rect 497502 371464 497548 371498
rect 497582 371464 497648 371498
rect 497682 371464 497748 371498
rect 497782 371464 497848 371498
rect 497882 371464 497948 371498
rect 497982 371464 498048 371498
rect 498082 371464 498114 371498
rect 497502 371398 498114 371464
rect 497502 371364 497548 371398
rect 497582 371364 497648 371398
rect 497682 371364 497748 371398
rect 497782 371364 497848 371398
rect 497882 371364 497948 371398
rect 497982 371364 498048 371398
rect 498082 371364 498114 371398
rect 497502 371298 498114 371364
rect 497502 371264 497548 371298
rect 497582 371264 497648 371298
rect 497682 371264 497748 371298
rect 497782 371264 497848 371298
rect 497882 371264 497948 371298
rect 497982 371264 498048 371298
rect 498082 371264 498114 371298
rect 497502 371198 498114 371264
rect 497502 371164 497548 371198
rect 497582 371164 497648 371198
rect 497682 371164 497748 371198
rect 497782 371164 497848 371198
rect 497882 371164 497948 371198
rect 497982 371164 498048 371198
rect 498082 371164 498114 371198
rect 497502 371098 498114 371164
rect 497502 371064 497548 371098
rect 497582 371064 497648 371098
rect 497682 371064 497748 371098
rect 497782 371064 497848 371098
rect 497882 371064 497948 371098
rect 497982 371064 498048 371098
rect 498082 371064 498114 371098
rect 497502 370854 498114 371064
rect 498688 371611 498808 371642
rect 498688 371577 498731 371611
rect 498765 371577 498808 371611
rect 498688 371411 498808 371577
rect 498688 371377 498731 371411
rect 498765 371377 498808 371411
rect 498688 371211 498808 371377
rect 498688 371177 498731 371211
rect 498765 371177 498808 371211
rect 498688 371011 498808 371177
rect 498688 370977 498731 371011
rect 498765 370977 498808 371011
rect 498208 370866 498260 370872
rect 497502 370826 498208 370854
rect 497502 370258 498114 370826
rect 498208 370808 498260 370814
rect 498688 370811 498808 370977
rect 497502 370224 497548 370258
rect 497582 370224 497648 370258
rect 497682 370224 497748 370258
rect 497782 370224 497848 370258
rect 497882 370224 497948 370258
rect 497982 370224 498048 370258
rect 498082 370224 498114 370258
rect 497502 370158 498114 370224
rect 497502 370124 497548 370158
rect 497582 370124 497648 370158
rect 497682 370124 497748 370158
rect 497782 370124 497848 370158
rect 497882 370124 497948 370158
rect 497982 370124 498048 370158
rect 498082 370124 498114 370158
rect 497502 370058 498114 370124
rect 497502 370024 497548 370058
rect 497582 370024 497648 370058
rect 497682 370024 497748 370058
rect 497782 370024 497848 370058
rect 497882 370024 497948 370058
rect 497982 370024 498048 370058
rect 498082 370024 498114 370058
rect 497502 369958 498114 370024
rect 497502 369924 497548 369958
rect 497582 369924 497648 369958
rect 497682 369924 497748 369958
rect 497782 369924 497848 369958
rect 497882 369924 497948 369958
rect 497982 369924 498048 369958
rect 498082 369924 498114 369958
rect 497502 369858 498114 369924
rect 497502 369824 497548 369858
rect 497582 369824 497648 369858
rect 497682 369824 497748 369858
rect 497782 369824 497848 369858
rect 497882 369824 497948 369858
rect 497982 369824 498048 369858
rect 498082 369824 498114 369858
rect 497502 369758 498114 369824
rect 497502 369724 497548 369758
rect 497582 369724 497648 369758
rect 497682 369724 497748 369758
rect 497782 369724 497848 369758
rect 497882 369724 497948 369758
rect 497982 369724 498048 369758
rect 498082 369724 498114 369758
rect 497502 368918 498114 369724
rect 497502 368884 497548 368918
rect 497582 368884 497648 368918
rect 497682 368884 497748 368918
rect 497782 368884 497848 368918
rect 497882 368884 497948 368918
rect 497982 368884 498048 368918
rect 498082 368884 498114 368918
rect 497502 368818 498114 368884
rect 497502 368784 497548 368818
rect 497582 368784 497648 368818
rect 497682 368784 497748 368818
rect 497782 368784 497848 368818
rect 497882 368784 497948 368818
rect 497982 368784 498048 368818
rect 498082 368784 498114 368818
rect 497502 368718 498114 368784
rect 497502 368684 497548 368718
rect 497582 368684 497648 368718
rect 497682 368684 497748 368718
rect 497782 368684 497848 368718
rect 497882 368684 497948 368718
rect 497982 368684 498048 368718
rect 498082 368684 498114 368718
rect 497502 368618 498114 368684
rect 497502 368584 497548 368618
rect 497582 368584 497648 368618
rect 497682 368584 497748 368618
rect 497782 368584 497848 368618
rect 497882 368584 497948 368618
rect 497982 368584 498048 368618
rect 498082 368584 498114 368618
rect 497502 368518 498114 368584
rect 497502 368484 497548 368518
rect 497582 368484 497648 368518
rect 497682 368484 497748 368518
rect 497782 368484 497848 368518
rect 497882 368484 497948 368518
rect 497982 368484 498048 368518
rect 498082 368484 498114 368518
rect 497502 368418 498114 368484
rect 497502 368384 497548 368418
rect 497582 368384 497648 368418
rect 497682 368384 497748 368418
rect 497782 368384 497848 368418
rect 497882 368384 497948 368418
rect 497982 368384 498048 368418
rect 498082 368384 498114 368418
rect 497502 367578 498114 368384
rect 497502 367544 497548 367578
rect 497582 367544 497648 367578
rect 497682 367544 497748 367578
rect 497782 367544 497848 367578
rect 497882 367544 497948 367578
rect 497982 367544 498048 367578
rect 498082 367544 498114 367578
rect 497502 367478 498114 367544
rect 497502 367444 497548 367478
rect 497582 367444 497648 367478
rect 497682 367444 497748 367478
rect 497782 367444 497848 367478
rect 497882 367444 497948 367478
rect 497982 367444 498048 367478
rect 498082 367444 498114 367478
rect 497502 367378 498114 367444
rect 497502 367344 497548 367378
rect 497582 367344 497648 367378
rect 497682 367344 497748 367378
rect 497782 367344 497848 367378
rect 497882 367344 497948 367378
rect 497982 367344 498048 367378
rect 498082 367344 498114 367378
rect 497502 367278 498114 367344
rect 497502 367244 497548 367278
rect 497582 367244 497648 367278
rect 497682 367244 497748 367278
rect 497782 367244 497848 367278
rect 497882 367244 497948 367278
rect 497982 367244 498048 367278
rect 498082 367244 498114 367278
rect 497502 367178 498114 367244
rect 497502 367144 497548 367178
rect 497582 367144 497648 367178
rect 497682 367144 497748 367178
rect 497782 367144 497848 367178
rect 497882 367144 497948 367178
rect 497982 367144 498048 367178
rect 498082 367144 498114 367178
rect 497502 367078 498114 367144
rect 497502 367044 497548 367078
rect 497582 367044 497648 367078
rect 497682 367044 497748 367078
rect 497782 367044 497848 367078
rect 497882 367044 497948 367078
rect 497982 367044 498048 367078
rect 498082 367044 498114 367078
rect 497502 366238 498114 367044
rect 497502 366204 497548 366238
rect 497582 366204 497648 366238
rect 497682 366204 497748 366238
rect 497782 366204 497848 366238
rect 497882 366204 497948 366238
rect 497982 366204 498048 366238
rect 498082 366204 498114 366238
rect 497502 366138 498114 366204
rect 497502 366104 497548 366138
rect 497582 366104 497648 366138
rect 497682 366104 497748 366138
rect 497782 366104 497848 366138
rect 497882 366104 497948 366138
rect 497982 366104 498048 366138
rect 498082 366104 498114 366138
rect 497502 366038 498114 366104
rect 497502 366004 497548 366038
rect 497582 366004 497648 366038
rect 497682 366004 497748 366038
rect 497782 366004 497848 366038
rect 497882 366004 497948 366038
rect 497982 366004 498048 366038
rect 498082 366004 498114 366038
rect 497502 365938 498114 366004
rect 497502 365904 497548 365938
rect 497582 365904 497648 365938
rect 497682 365904 497748 365938
rect 497782 365904 497848 365938
rect 497882 365904 497948 365938
rect 497982 365904 498048 365938
rect 498082 365904 498114 365938
rect 497502 365838 498114 365904
rect 497502 365804 497548 365838
rect 497582 365804 497648 365838
rect 497682 365804 497748 365838
rect 497782 365804 497848 365838
rect 497882 365804 497948 365838
rect 497982 365804 498048 365838
rect 498082 365804 498114 365838
rect 497502 365738 498114 365804
rect 497502 365704 497548 365738
rect 497582 365704 497648 365738
rect 497682 365704 497748 365738
rect 497782 365704 497848 365738
rect 497882 365704 497948 365738
rect 497982 365704 498048 365738
rect 498082 365704 498114 365738
rect 497502 364898 498114 365704
rect 497502 364864 497548 364898
rect 497582 364864 497648 364898
rect 497682 364864 497748 364898
rect 497782 364864 497848 364898
rect 497882 364864 497948 364898
rect 497982 364864 498048 364898
rect 498082 364864 498114 364898
rect 497502 364798 498114 364864
rect 497502 364764 497548 364798
rect 497582 364764 497648 364798
rect 497682 364764 497748 364798
rect 497782 364764 497848 364798
rect 497882 364764 497948 364798
rect 497982 364764 498048 364798
rect 498082 364764 498114 364798
rect 497502 364698 498114 364764
rect 497502 364664 497548 364698
rect 497582 364664 497648 364698
rect 497682 364664 497748 364698
rect 497782 364664 497848 364698
rect 497882 364664 497948 364698
rect 497982 364664 498048 364698
rect 498082 364664 498114 364698
rect 497502 364598 498114 364664
rect 497502 364564 497548 364598
rect 497582 364564 497648 364598
rect 497682 364564 497748 364598
rect 497782 364564 497848 364598
rect 497882 364564 497948 364598
rect 497982 364564 498048 364598
rect 498082 364564 498114 364598
rect 497502 364498 498114 364564
rect 497502 364464 497548 364498
rect 497582 364464 497648 364498
rect 497682 364464 497748 364498
rect 497782 364464 497848 364498
rect 497882 364464 497948 364498
rect 497982 364464 498048 364498
rect 498082 364464 498114 364498
rect 497502 364398 498114 364464
rect 497502 364364 497548 364398
rect 497582 364364 497648 364398
rect 497682 364364 497748 364398
rect 497782 364364 497848 364398
rect 497882 364364 497948 364398
rect 497982 364364 498048 364398
rect 498082 364364 498114 364398
rect 497502 363558 498114 364364
rect 497502 363524 497548 363558
rect 497582 363524 497648 363558
rect 497682 363524 497748 363558
rect 497782 363524 497848 363558
rect 497882 363524 497948 363558
rect 497982 363524 498048 363558
rect 498082 363524 498114 363558
rect 497502 363458 498114 363524
rect 497502 363424 497548 363458
rect 497582 363424 497648 363458
rect 497682 363424 497748 363458
rect 497782 363424 497848 363458
rect 497882 363424 497948 363458
rect 497982 363424 498048 363458
rect 498082 363424 498114 363458
rect 497502 363358 498114 363424
rect 497502 363324 497548 363358
rect 497582 363324 497648 363358
rect 497682 363324 497748 363358
rect 497782 363324 497848 363358
rect 497882 363324 497948 363358
rect 497982 363324 498048 363358
rect 498082 363324 498114 363358
rect 497502 363258 498114 363324
rect 497502 363224 497548 363258
rect 497582 363224 497648 363258
rect 497682 363224 497748 363258
rect 497782 363224 497848 363258
rect 497882 363224 497948 363258
rect 497982 363224 498048 363258
rect 498082 363224 498114 363258
rect 497502 363158 498114 363224
rect 497502 363124 497548 363158
rect 497582 363124 497648 363158
rect 497682 363124 497748 363158
rect 497782 363124 497848 363158
rect 497882 363124 497948 363158
rect 497982 363124 498048 363158
rect 498082 363124 498114 363158
rect 497502 363058 498114 363124
rect 497502 363024 497548 363058
rect 497582 363024 497648 363058
rect 497682 363024 497748 363058
rect 497782 363024 497848 363058
rect 497882 363024 497948 363058
rect 497982 363024 498048 363058
rect 498082 363024 498114 363058
rect 497502 362978 498114 363024
rect 498688 370777 498731 370811
rect 498765 370777 498808 370811
rect 498688 370611 498808 370777
rect 498688 370577 498731 370611
rect 498765 370577 498808 370611
rect 498688 370411 498808 370577
rect 498688 370377 498731 370411
rect 498765 370377 498808 370411
rect 498688 370211 498808 370377
rect 498688 370177 498731 370211
rect 498765 370177 498808 370211
rect 498688 370011 498808 370177
rect 498688 369977 498731 370011
rect 498765 369977 498808 370011
rect 498688 369811 498808 369977
rect 498688 369777 498731 369811
rect 498765 369777 498808 369811
rect 498688 369611 498808 369777
rect 498688 369577 498731 369611
rect 498765 369577 498808 369611
rect 498688 369411 498808 369577
rect 498688 369377 498731 369411
rect 498765 369377 498808 369411
rect 498688 369211 498808 369377
rect 498688 369177 498731 369211
rect 498765 369177 498808 369211
rect 498688 369011 498808 369177
rect 498688 368977 498731 369011
rect 498765 368977 498808 369011
rect 498688 368811 498808 368977
rect 498688 368777 498731 368811
rect 498765 368777 498808 368811
rect 498688 368611 498808 368777
rect 498688 368577 498731 368611
rect 498765 368577 498808 368611
rect 498688 368411 498808 368577
rect 498688 368377 498731 368411
rect 498765 368377 498808 368411
rect 498688 368211 498808 368377
rect 498688 368177 498731 368211
rect 498765 368177 498808 368211
rect 498688 368011 498808 368177
rect 498688 367977 498731 368011
rect 498765 367977 498808 368011
rect 498688 367811 498808 367977
rect 498688 367777 498731 367811
rect 498765 367777 498808 367811
rect 498688 367611 498808 367777
rect 498688 367577 498731 367611
rect 498765 367577 498808 367611
rect 498688 367411 498808 367577
rect 498688 367377 498731 367411
rect 498765 367377 498808 367411
rect 498688 367211 498808 367377
rect 498688 367177 498731 367211
rect 498765 367177 498808 367211
rect 498688 367011 498808 367177
rect 498688 366977 498731 367011
rect 498765 366977 498808 367011
rect 498688 366811 498808 366977
rect 498688 366777 498731 366811
rect 498765 366777 498808 366811
rect 498688 366611 498808 366777
rect 498688 366577 498731 366611
rect 498765 366577 498808 366611
rect 498688 366411 498808 366577
rect 498688 366377 498731 366411
rect 498765 366377 498808 366411
rect 498688 366211 498808 366377
rect 498688 366177 498731 366211
rect 498765 366177 498808 366211
rect 498688 366011 498808 366177
rect 498688 365977 498731 366011
rect 498765 365977 498808 366011
rect 498688 365811 498808 365977
rect 498688 365777 498731 365811
rect 498765 365777 498808 365811
rect 498688 365611 498808 365777
rect 498688 365577 498731 365611
rect 498765 365577 498808 365611
rect 498688 365411 498808 365577
rect 498688 365377 498731 365411
rect 498765 365377 498808 365411
rect 498688 365211 498808 365377
rect 498688 365177 498731 365211
rect 498765 365177 498808 365211
rect 498688 365011 498808 365177
rect 498688 364977 498731 365011
rect 498765 364977 498808 365011
rect 498688 364811 498808 364977
rect 498688 364777 498731 364811
rect 498765 364777 498808 364811
rect 498688 364611 498808 364777
rect 498688 364577 498731 364611
rect 498765 364577 498808 364611
rect 498688 364411 498808 364577
rect 498688 364377 498731 364411
rect 498765 364377 498808 364411
rect 498688 364211 498808 364377
rect 498688 364177 498731 364211
rect 498765 364177 498808 364211
rect 498688 364011 498808 364177
rect 498688 363977 498731 364011
rect 498765 363977 498808 364011
rect 498688 363811 498808 363977
rect 498688 363777 498731 363811
rect 498765 363777 498808 363811
rect 498688 363611 498808 363777
rect 498688 363577 498731 363611
rect 498765 363577 498808 363611
rect 498688 363411 498808 363577
rect 498688 363377 498731 363411
rect 498765 363377 498808 363411
rect 498688 363211 498808 363377
rect 498688 363177 498731 363211
rect 498765 363177 498808 363211
rect 498688 363011 498808 363177
rect 497328 362900 497344 362934
rect 497378 362900 497398 362934
rect 497328 362844 497398 362900
rect 497328 362810 497344 362844
rect 497378 362810 497398 362844
rect 497328 362804 497398 362810
rect 498688 362977 498731 363011
rect 498765 362977 498808 363011
rect 498688 362811 498808 362977
rect 497178 362738 497248 362794
rect 497178 362704 497184 362738
rect 497218 362704 497248 362738
rect 497178 362640 497248 362704
rect 498688 362777 498731 362811
rect 498765 362777 498808 362811
rect 496808 359888 496810 361476
rect 496926 359888 496928 361476
rect 496808 359866 496928 359888
rect 494928 357440 494930 359028
rect 495046 357440 495048 359028
rect 494928 357418 495048 357440
rect 498688 359028 498808 362777
rect 500568 411584 500688 411606
rect 500568 409996 500570 411584
rect 500686 409996 500688 411584
rect 500568 408461 500688 409996
rect 500568 408427 500611 408461
rect 500645 408427 500688 408461
rect 500568 408061 500688 408427
rect 500568 408027 500611 408061
rect 500645 408027 500688 408061
rect 500568 407661 500688 408027
rect 500568 407627 500611 407661
rect 500645 407627 500688 407661
rect 500568 407261 500688 407627
rect 500568 407227 500611 407261
rect 500645 407227 500688 407261
rect 500568 406861 500688 407227
rect 500568 406827 500611 406861
rect 500645 406827 500688 406861
rect 500568 406461 500688 406827
rect 500568 406427 500611 406461
rect 500645 406427 500688 406461
rect 500568 406061 500688 406427
rect 500568 406027 500611 406061
rect 500645 406027 500688 406061
rect 500568 405661 500688 406027
rect 500568 405627 500611 405661
rect 500645 405627 500688 405661
rect 500568 405261 500688 405627
rect 500568 405227 500611 405261
rect 500645 405227 500688 405261
rect 500568 404861 500688 405227
rect 500568 404827 500611 404861
rect 500645 404827 500688 404861
rect 500568 404461 500688 404827
rect 500568 404427 500611 404461
rect 500645 404427 500688 404461
rect 500568 404061 500688 404427
rect 500568 404027 500611 404061
rect 500645 404027 500688 404061
rect 500568 403661 500688 404027
rect 500568 403627 500611 403661
rect 500645 403627 500688 403661
rect 500568 403261 500688 403627
rect 500568 403227 500611 403261
rect 500645 403227 500688 403261
rect 500568 402861 500688 403227
rect 500568 402827 500611 402861
rect 500645 402827 500688 402861
rect 500568 402461 500688 402827
rect 500568 402427 500611 402461
rect 500645 402427 500688 402461
rect 500568 402061 500688 402427
rect 500568 402027 500611 402061
rect 500645 402027 500688 402061
rect 500568 401661 500688 402027
rect 500568 401627 500611 401661
rect 500645 401627 500688 401661
rect 500568 399641 500688 401627
rect 500568 399607 500611 399641
rect 500645 399607 500688 399641
rect 500568 399241 500688 399607
rect 500568 399207 500611 399241
rect 500645 399207 500688 399241
rect 500568 398841 500688 399207
rect 500568 398807 500611 398841
rect 500645 398807 500688 398841
rect 500568 398441 500688 398807
rect 500568 398407 500611 398441
rect 500645 398407 500688 398441
rect 500568 398041 500688 398407
rect 500568 398007 500611 398041
rect 500645 398007 500688 398041
rect 500568 397641 500688 398007
rect 500568 397607 500611 397641
rect 500645 397607 500688 397641
rect 500568 397241 500688 397607
rect 500568 397207 500611 397241
rect 500645 397207 500688 397241
rect 500568 396841 500688 397207
rect 500568 396807 500611 396841
rect 500645 396807 500688 396841
rect 500568 396441 500688 396807
rect 500568 396407 500611 396441
rect 500645 396407 500688 396441
rect 500568 396041 500688 396407
rect 500568 396007 500611 396041
rect 500645 396007 500688 396041
rect 500568 395641 500688 396007
rect 500568 395607 500611 395641
rect 500645 395607 500688 395641
rect 500568 395241 500688 395607
rect 500568 395207 500611 395241
rect 500645 395207 500688 395241
rect 500568 394841 500688 395207
rect 500568 394807 500611 394841
rect 500645 394807 500688 394841
rect 500568 394441 500688 394807
rect 500568 394407 500611 394441
rect 500645 394407 500688 394441
rect 500568 394041 500688 394407
rect 500568 394007 500611 394041
rect 500645 394007 500688 394041
rect 500568 393641 500688 394007
rect 500568 393607 500611 393641
rect 500645 393607 500688 393641
rect 500568 393241 500688 393607
rect 500568 393207 500611 393241
rect 500645 393207 500688 393241
rect 500568 392841 500688 393207
rect 500568 392807 500611 392841
rect 500645 392807 500688 392841
rect 500568 392097 500688 392807
rect 502448 408461 502568 412444
rect 506208 414032 506328 414054
rect 506208 412444 506210 414032
rect 506326 412444 506328 414032
rect 502448 408427 502491 408461
rect 502525 408427 502568 408461
rect 502448 408061 502568 408427
rect 502448 408027 502491 408061
rect 502525 408027 502568 408061
rect 502448 407661 502568 408027
rect 502448 407627 502491 407661
rect 502525 407627 502568 407661
rect 502448 407261 502568 407627
rect 502448 407227 502491 407261
rect 502525 407227 502568 407261
rect 502448 406861 502568 407227
rect 502448 406827 502491 406861
rect 502525 406827 502568 406861
rect 502448 406461 502568 406827
rect 502448 406427 502491 406461
rect 502525 406427 502568 406461
rect 502448 406061 502568 406427
rect 502448 406027 502491 406061
rect 502525 406027 502568 406061
rect 502448 405661 502568 406027
rect 502448 405627 502491 405661
rect 502525 405627 502568 405661
rect 502448 405261 502568 405627
rect 502448 405227 502491 405261
rect 502525 405227 502568 405261
rect 502448 404861 502568 405227
rect 502448 404827 502491 404861
rect 502525 404827 502568 404861
rect 502448 404461 502568 404827
rect 502448 404427 502491 404461
rect 502525 404427 502568 404461
rect 502448 404061 502568 404427
rect 502448 404027 502491 404061
rect 502525 404027 502568 404061
rect 502448 403661 502568 404027
rect 502448 403627 502491 403661
rect 502525 403627 502568 403661
rect 502448 403261 502568 403627
rect 502448 403227 502491 403261
rect 502525 403227 502568 403261
rect 502448 402861 502568 403227
rect 502448 402827 502491 402861
rect 502525 402827 502568 402861
rect 502448 402461 502568 402827
rect 502448 402427 502491 402461
rect 502525 402427 502568 402461
rect 502448 402061 502568 402427
rect 502448 402027 502491 402061
rect 502525 402027 502568 402061
rect 502448 401661 502568 402027
rect 502448 401627 502491 401661
rect 502525 401627 502568 401661
rect 502448 399641 502568 401627
rect 504328 411584 504448 411606
rect 504328 409996 504330 411584
rect 504446 409996 504448 411584
rect 504328 402779 504448 409996
rect 504328 402745 504371 402779
rect 504405 402745 504448 402779
rect 504328 402579 504448 402745
rect 506208 402779 506328 412444
rect 509968 414032 510088 414054
rect 509968 412444 509970 414032
rect 510086 412444 510088 414032
rect 506208 402745 506251 402779
rect 506285 402745 506328 402779
rect 504328 402545 504371 402579
rect 504405 402545 504448 402579
rect 504328 402379 504448 402545
rect 504328 402345 504371 402379
rect 504405 402345 504448 402379
rect 504328 402179 504448 402345
rect 504328 402145 504371 402179
rect 504405 402145 504448 402179
rect 504328 401979 504448 402145
rect 505023 402566 505633 402597
rect 505023 402532 505068 402566
rect 505102 402532 505168 402566
rect 505202 402532 505268 402566
rect 505302 402532 505368 402566
rect 505402 402532 505468 402566
rect 505502 402532 505568 402566
rect 505602 402532 505633 402566
rect 505023 402466 505633 402532
rect 505023 402432 505068 402466
rect 505102 402432 505168 402466
rect 505202 402432 505268 402466
rect 505302 402432 505368 402466
rect 505402 402432 505468 402466
rect 505502 402432 505568 402466
rect 505602 402432 505633 402466
rect 505023 402366 505633 402432
rect 505023 402332 505068 402366
rect 505102 402332 505168 402366
rect 505202 402332 505268 402366
rect 505302 402332 505368 402366
rect 505402 402332 505468 402366
rect 505502 402332 505568 402366
rect 505602 402332 505633 402366
rect 505023 402266 505633 402332
rect 505023 402232 505068 402266
rect 505102 402232 505168 402266
rect 505202 402232 505268 402266
rect 505302 402232 505368 402266
rect 505402 402232 505468 402266
rect 505502 402232 505568 402266
rect 505602 402232 505633 402266
rect 505023 402166 505633 402232
rect 505023 402132 505068 402166
rect 505102 402132 505168 402166
rect 505202 402132 505268 402166
rect 505302 402132 505368 402166
rect 505402 402132 505468 402166
rect 505502 402132 505568 402166
rect 505602 402132 505633 402166
rect 505023 402066 505633 402132
rect 504872 402054 504924 402060
rect 505023 402042 505068 402066
rect 504924 402032 505068 402042
rect 505102 402032 505168 402066
rect 505202 402032 505268 402066
rect 505302 402032 505368 402066
rect 505402 402032 505468 402066
rect 505502 402032 505568 402066
rect 505602 402032 505633 402066
rect 504924 402014 505633 402032
rect 504872 401996 504924 402002
rect 505023 401987 505633 402014
rect 506208 402579 506328 402745
rect 506208 402545 506251 402579
rect 506285 402545 506328 402579
rect 506208 402379 506328 402545
rect 506208 402345 506251 402379
rect 506285 402345 506328 402379
rect 506208 402179 506328 402345
rect 506208 402145 506251 402179
rect 506285 402145 506328 402179
rect 504328 401945 504371 401979
rect 504405 401945 504448 401979
rect 504328 401779 504448 401945
rect 506208 401979 506328 402145
rect 506208 401945 506251 401979
rect 506285 401945 506328 401979
rect 505759 401861 505805 401873
rect 505759 401827 505765 401861
rect 505799 401858 505805 401861
rect 505799 401830 505932 401858
rect 505799 401827 505805 401830
rect 505759 401815 505805 401827
rect 504328 401745 504371 401779
rect 504405 401745 504448 401779
rect 504328 401093 504448 401745
rect 505904 401689 505932 401830
rect 506208 401779 506328 401945
rect 506208 401745 506251 401779
rect 506285 401745 506328 401779
rect 505895 401677 505941 401689
rect 505895 401643 505901 401677
rect 505935 401674 505941 401677
rect 506208 401674 506328 401745
rect 505935 401646 506328 401674
rect 505935 401643 505941 401646
rect 505895 401631 505941 401643
rect 504328 401059 504371 401093
rect 504405 401059 504448 401093
rect 504328 400893 504448 401059
rect 504328 400859 504371 400893
rect 504405 400859 504448 400893
rect 504328 400693 504448 400859
rect 504627 401257 505189 401265
rect 504627 400863 504639 401257
rect 505177 400863 505189 401257
rect 504627 400855 505189 400863
rect 505587 401257 506149 401265
rect 505587 400863 505599 401257
rect 506137 401042 506149 401257
rect 506148 400990 506149 401042
rect 506137 400863 506149 400990
rect 505587 400855 506149 400863
rect 506208 401093 506328 401646
rect 506208 401059 506251 401093
rect 506285 401059 506328 401093
rect 506208 400893 506328 401059
rect 506208 400859 506251 400893
rect 506285 400859 506328 400893
rect 504328 400659 504371 400693
rect 504405 400659 504448 400693
rect 503920 400582 503972 400588
rect 503972 400542 504028 400570
rect 503920 400524 503972 400530
rect 502448 399607 502491 399641
rect 502525 399607 502568 399641
rect 502448 399478 502568 399607
rect 502448 399426 502492 399478
rect 502544 399426 502568 399478
rect 502448 399241 502568 399426
rect 502448 399207 502491 399241
rect 502525 399207 502568 399241
rect 502448 398841 502568 399207
rect 502448 398807 502491 398841
rect 502525 398807 502568 398841
rect 502448 398441 502568 398807
rect 502448 398407 502491 398441
rect 502525 398407 502568 398441
rect 502448 398041 502568 398407
rect 502448 398007 502491 398041
rect 502525 398007 502568 398041
rect 502448 397641 502568 398007
rect 502448 397607 502491 397641
rect 502525 397607 502568 397641
rect 502448 397241 502568 397607
rect 502448 397207 502491 397241
rect 502525 397207 502568 397241
rect 502448 396841 502568 397207
rect 502448 396807 502491 396841
rect 502525 396807 502568 396841
rect 502448 396441 502568 396807
rect 502448 396407 502491 396441
rect 502525 396407 502568 396441
rect 502448 396041 502568 396407
rect 502448 396007 502491 396041
rect 502525 396007 502568 396041
rect 502448 395641 502568 396007
rect 502448 395607 502491 395641
rect 502525 395607 502568 395641
rect 502448 395241 502568 395607
rect 502448 395207 502491 395241
rect 502525 395207 502568 395241
rect 502448 394841 502568 395207
rect 502448 394807 502491 394841
rect 502525 394807 502568 394841
rect 502448 394441 502568 394807
rect 502448 394407 502491 394441
rect 502525 394407 502568 394441
rect 502448 394041 502568 394407
rect 502448 394007 502491 394041
rect 502525 394007 502568 394041
rect 502448 393641 502568 394007
rect 502448 393607 502491 393641
rect 502525 393607 502568 393641
rect 502448 393241 502568 393607
rect 502448 393207 502491 393241
rect 502525 393207 502568 393241
rect 502448 392841 502568 393207
rect 502448 392807 502491 392841
rect 502525 392807 502568 392841
rect 502220 392762 502272 392768
rect 502220 392704 502272 392710
rect 500863 392233 502153 392239
rect 500863 392199 500879 392233
rect 500913 392199 500951 392233
rect 500985 392199 501023 392233
rect 501057 392199 501095 392233
rect 501129 392199 501167 392233
rect 501201 392199 501239 392233
rect 501273 392199 501311 392233
rect 501345 392199 501383 392233
rect 501417 392199 501455 392233
rect 501489 392199 501527 392233
rect 501561 392199 501599 392233
rect 501633 392199 501671 392233
rect 501705 392199 501743 392233
rect 501777 392199 501815 392233
rect 501849 392199 501887 392233
rect 501921 392199 501959 392233
rect 501993 392199 502031 392233
rect 502065 392199 502103 392233
rect 502137 392199 502153 392233
rect 502232 392213 502260 392704
rect 500863 392193 502153 392199
rect 502223 392201 502269 392213
rect 502223 392167 502229 392201
rect 502263 392167 502269 392201
rect 502223 392155 502269 392167
rect 500568 392063 500611 392097
rect 500645 392063 500688 392097
rect 500568 391697 500688 392063
rect 502448 392097 502568 392807
rect 502448 392063 502491 392097
rect 502525 392063 502568 392097
rect 500863 391775 502153 391781
rect 500863 391741 500879 391775
rect 500913 391741 500951 391775
rect 500985 391741 501023 391775
rect 501057 391741 501095 391775
rect 501129 391741 501167 391775
rect 501201 391741 501239 391775
rect 501273 391741 501311 391775
rect 501345 391741 501383 391775
rect 501417 391741 501455 391775
rect 501489 391741 501527 391775
rect 501561 391741 501599 391775
rect 501633 391741 501671 391775
rect 501705 391741 501743 391775
rect 501777 391741 501815 391775
rect 501849 391741 501887 391775
rect 501921 391741 501959 391775
rect 501993 391741 502031 391775
rect 502065 391741 502103 391775
rect 502137 391741 502153 391775
rect 500863 391735 502153 391741
rect 500568 391663 500611 391697
rect 500645 391663 500688 391697
rect 500568 391297 500688 391663
rect 502448 391697 502568 392063
rect 502448 391663 502491 391697
rect 502525 391663 502568 391697
rect 500568 391263 500611 391297
rect 500645 391263 500688 391297
rect 500863 391317 502153 391323
rect 500863 391283 500879 391317
rect 500913 391283 500951 391317
rect 500985 391283 501023 391317
rect 501057 391283 501095 391317
rect 501129 391283 501167 391317
rect 501201 391283 501239 391317
rect 501273 391283 501311 391317
rect 501345 391283 501383 391317
rect 501417 391283 501455 391317
rect 501489 391283 501527 391317
rect 501561 391283 501599 391317
rect 501633 391283 501671 391317
rect 501705 391283 501743 391317
rect 501777 391283 501815 391317
rect 501849 391283 501887 391317
rect 501921 391283 501959 391317
rect 501993 391283 502031 391317
rect 502065 391283 502103 391317
rect 502137 391283 502153 391317
rect 500863 391277 502153 391283
rect 502448 391297 502568 391663
rect 500568 390897 500688 391263
rect 502448 391263 502491 391297
rect 502525 391263 502568 391297
rect 502220 391198 502272 391204
rect 502220 391140 502272 391146
rect 500568 390863 500611 390897
rect 500645 390863 500688 390897
rect 500568 390497 500688 390863
rect 500863 390859 502153 390865
rect 500863 390825 500879 390859
rect 500913 390825 500951 390859
rect 500985 390825 501023 390859
rect 501057 390825 501095 390859
rect 501129 390825 501167 390859
rect 501201 390825 501239 390859
rect 501273 390825 501311 390859
rect 501345 390825 501383 390859
rect 501417 390825 501455 390859
rect 501489 390825 501527 390859
rect 501561 390825 501599 390859
rect 501633 390825 501671 390859
rect 501705 390825 501743 390859
rect 501777 390825 501815 390859
rect 501849 390825 501887 390859
rect 501921 390825 501959 390859
rect 501993 390825 502031 390859
rect 502065 390825 502103 390859
rect 502137 390825 502153 390859
rect 500863 390819 502153 390825
rect 500568 390463 500611 390497
rect 500645 390463 500688 390497
rect 500568 390097 500688 390463
rect 500863 390401 502153 390407
rect 500863 390367 500879 390401
rect 500913 390367 500951 390401
rect 500985 390367 501023 390401
rect 501057 390367 501095 390401
rect 501129 390367 501167 390401
rect 501201 390367 501239 390401
rect 501273 390367 501311 390401
rect 501345 390367 501383 390401
rect 501417 390367 501455 390401
rect 501489 390367 501527 390401
rect 501561 390367 501599 390401
rect 501633 390367 501671 390401
rect 501705 390367 501743 390401
rect 501777 390367 501815 390401
rect 501849 390367 501887 390401
rect 501921 390367 501959 390401
rect 501993 390367 502031 390401
rect 502065 390367 502103 390401
rect 502137 390367 502153 390401
rect 500863 390361 502153 390367
rect 500568 390063 500611 390097
rect 500645 390082 500688 390097
rect 500795 390085 500841 390097
rect 500795 390082 500801 390085
rect 500645 390063 500801 390082
rect 500568 390054 500801 390063
rect 500568 389697 500688 390054
rect 500795 390051 500801 390054
rect 500835 390051 500841 390085
rect 500795 390039 500841 390051
rect 500863 389943 502153 389949
rect 500863 389909 500879 389943
rect 500913 389909 500951 389943
rect 500985 389909 501023 389943
rect 501057 389909 501095 389943
rect 501129 389909 501167 389943
rect 501201 389909 501239 389943
rect 501273 389909 501311 389943
rect 501345 389909 501383 389943
rect 501417 389909 501455 389943
rect 501489 389909 501527 389943
rect 501561 389909 501599 389943
rect 501633 389909 501671 389943
rect 501705 389909 501743 389943
rect 501777 389909 501815 389943
rect 501849 389909 501887 389943
rect 501921 389909 501959 389943
rect 501993 389909 502031 389943
rect 502065 389909 502103 389943
rect 502137 389909 502153 389943
rect 500863 389903 502153 389909
rect 500568 389663 500611 389697
rect 500645 389663 500688 389697
rect 500568 389297 500688 389663
rect 500863 389485 502153 389491
rect 500863 389451 500879 389485
rect 500913 389451 500951 389485
rect 500985 389451 501023 389485
rect 501057 389451 501095 389485
rect 501129 389451 501167 389485
rect 501201 389451 501239 389485
rect 501273 389451 501311 389485
rect 501345 389451 501383 389485
rect 501417 389451 501455 389485
rect 501489 389451 501527 389485
rect 501561 389451 501599 389485
rect 501633 389451 501671 389485
rect 501705 389451 501743 389485
rect 501777 389451 501815 389485
rect 501849 389451 501887 389485
rect 501921 389451 501959 389485
rect 501993 389451 502031 389485
rect 502065 389451 502103 389485
rect 502137 389451 502153 389485
rect 500863 389445 502153 389451
rect 500568 389263 500611 389297
rect 500645 389263 500688 389297
rect 500568 388897 500688 389263
rect 500863 389027 502153 389033
rect 500863 388993 500879 389027
rect 500913 388993 500951 389027
rect 500985 388993 501023 389027
rect 501057 388993 501095 389027
rect 501129 388993 501167 389027
rect 501201 388993 501239 389027
rect 501273 388993 501311 389027
rect 501345 388993 501383 389027
rect 501417 388993 501455 389027
rect 501489 388993 501527 389027
rect 501561 388993 501599 389027
rect 501633 388993 501671 389027
rect 501705 388993 501743 389027
rect 501777 388993 501815 389027
rect 501849 388993 501887 389027
rect 501921 388993 501959 389027
rect 501993 388993 502031 389027
rect 502065 388993 502103 389027
rect 502137 388993 502153 389027
rect 500863 388987 502153 388993
rect 500568 388863 500611 388897
rect 500645 388863 500688 388897
rect 500568 388497 500688 388863
rect 500863 388569 502153 388575
rect 500863 388535 500879 388569
rect 500913 388535 500951 388569
rect 500985 388535 501023 388569
rect 501057 388535 501095 388569
rect 501129 388535 501167 388569
rect 501201 388535 501239 388569
rect 501273 388535 501311 388569
rect 501345 388535 501383 388569
rect 501417 388535 501455 388569
rect 501489 388535 501527 388569
rect 501561 388535 501599 388569
rect 501633 388535 501671 388569
rect 501705 388535 501743 388569
rect 501777 388535 501815 388569
rect 501849 388535 501887 388569
rect 501921 388535 501959 388569
rect 501993 388535 502031 388569
rect 502065 388535 502103 388569
rect 502137 388535 502153 388569
rect 500863 388529 502153 388535
rect 500568 388463 500611 388497
rect 500645 388463 500688 388497
rect 500568 388097 500688 388463
rect 500568 388063 500611 388097
rect 500645 388063 500688 388097
rect 500863 388111 502153 388117
rect 500863 388077 500879 388111
rect 500913 388077 500951 388111
rect 500985 388077 501023 388111
rect 501057 388077 501095 388111
rect 501129 388077 501167 388111
rect 501201 388077 501239 388111
rect 501273 388077 501311 388111
rect 501345 388077 501383 388111
rect 501417 388077 501455 388111
rect 501489 388077 501527 388111
rect 501561 388077 501599 388111
rect 501633 388077 501671 388111
rect 501705 388077 501743 388111
rect 501777 388077 501815 388111
rect 501849 388077 501887 388111
rect 501921 388077 501959 388111
rect 501993 388077 502031 388111
rect 502065 388077 502103 388111
rect 502137 388077 502153 388111
rect 500863 388071 502153 388077
rect 500568 387697 500688 388063
rect 500568 387663 500611 387697
rect 500645 387663 500688 387697
rect 500568 387297 500688 387663
rect 500863 387653 502153 387659
rect 500863 387619 500879 387653
rect 500913 387619 500951 387653
rect 500985 387619 501023 387653
rect 501057 387619 501095 387653
rect 501129 387619 501167 387653
rect 501201 387619 501239 387653
rect 501273 387619 501311 387653
rect 501345 387619 501383 387653
rect 501417 387619 501455 387653
rect 501489 387619 501527 387653
rect 501561 387619 501599 387653
rect 501633 387619 501671 387653
rect 501705 387619 501743 387653
rect 501777 387619 501815 387653
rect 501849 387619 501887 387653
rect 501921 387619 501959 387653
rect 501993 387619 502031 387653
rect 502065 387619 502103 387653
rect 502137 387619 502153 387653
rect 500863 387613 502153 387619
rect 500568 387263 500611 387297
rect 500645 387263 500688 387297
rect 500568 386897 500688 387263
rect 500863 387195 502153 387201
rect 500863 387161 500879 387195
rect 500913 387161 500951 387195
rect 500985 387161 501023 387195
rect 501057 387161 501095 387195
rect 501129 387161 501167 387195
rect 501201 387161 501239 387195
rect 501273 387161 501311 387195
rect 501345 387161 501383 387195
rect 501417 387161 501455 387195
rect 501489 387161 501527 387195
rect 501561 387161 501599 387195
rect 501633 387161 501671 387195
rect 501705 387161 501743 387195
rect 501777 387161 501815 387195
rect 501849 387161 501887 387195
rect 501921 387161 501959 387195
rect 501993 387161 502031 387195
rect 502065 387161 502103 387195
rect 502137 387161 502153 387195
rect 500863 387155 502153 387161
rect 502232 387046 502260 391140
rect 502448 390897 502568 391263
rect 502448 390863 502491 390897
rect 502525 390863 502568 390897
rect 502448 390497 502568 390863
rect 502448 390463 502491 390497
rect 502525 390463 502568 390497
rect 502448 390097 502568 390463
rect 502448 390063 502491 390097
rect 502525 390063 502568 390097
rect 502448 389697 502568 390063
rect 502448 389663 502491 389697
rect 502525 389663 502568 389697
rect 502448 389297 502568 389663
rect 502448 389263 502491 389297
rect 502525 389263 502568 389297
rect 502448 388897 502568 389263
rect 504000 389180 504028 400542
rect 504328 400493 504448 400659
rect 504328 400459 504371 400493
rect 504405 400459 504448 400493
rect 504328 400293 504448 400459
rect 504328 400259 504371 400293
rect 504405 400259 504448 400293
rect 504328 400093 504448 400259
rect 504328 400059 504371 400093
rect 504405 400059 504448 400093
rect 504328 399893 504448 400059
rect 504328 399859 504371 399893
rect 504405 399859 504448 399893
rect 504328 399693 504448 399859
rect 504328 399659 504371 399693
rect 504405 399659 504448 399693
rect 504328 399493 504448 399659
rect 504328 399459 504371 399493
rect 504405 399459 504448 399493
rect 504328 399293 504448 399459
rect 505156 399392 505184 400855
rect 506208 400693 506328 400859
rect 506208 400659 506251 400693
rect 506285 400659 506328 400693
rect 506208 400493 506328 400659
rect 506208 400459 506251 400493
rect 506285 400459 506328 400493
rect 506208 400293 506328 400459
rect 506208 400259 506251 400293
rect 506285 400259 506328 400293
rect 506208 400093 506328 400259
rect 506208 400059 506251 400093
rect 506285 400059 506328 400093
rect 506208 399893 506328 400059
rect 506208 399859 506251 399893
rect 506285 399859 506328 399893
rect 506208 399693 506328 399859
rect 506208 399659 506251 399693
rect 506285 399659 506328 399693
rect 506208 399493 506328 399659
rect 506208 399459 506251 399493
rect 506285 399459 506328 399493
rect 505144 399386 505196 399392
rect 505144 399328 505196 399334
rect 504328 399259 504371 399293
rect 504405 399259 504448 399293
rect 506208 399293 506328 399459
rect 504328 399093 504448 399259
rect 505189 399257 506153 399268
rect 504328 399059 504371 399093
rect 504405 399059 504448 399093
rect 504328 398349 504448 399059
rect 504627 399250 506153 399257
rect 504627 398856 504639 399250
rect 505177 398856 505599 399250
rect 506137 398856 506153 399250
rect 504627 398847 506153 398856
rect 505189 398836 506153 398847
rect 506208 399259 506251 399293
rect 506285 399259 506328 399293
rect 506208 399093 506328 399259
rect 506208 399059 506251 399093
rect 506285 399059 506328 399093
rect 505620 398742 505672 398748
rect 505620 398684 505672 398690
rect 505632 398521 505660 398684
rect 504328 398315 504371 398349
rect 504405 398315 504448 398349
rect 504328 398149 504448 398315
rect 504328 398115 504371 398149
rect 504405 398115 504448 398149
rect 504328 397949 504448 398115
rect 504627 398513 505189 398521
rect 504627 398119 504639 398513
rect 505177 398380 505189 398513
rect 505587 398513 506149 398521
rect 505177 398374 505196 398380
rect 505177 398316 505196 398322
rect 505177 398119 505189 398316
rect 504627 398111 505189 398119
rect 505587 398119 505599 398513
rect 506137 398119 506149 398513
rect 505587 398111 506149 398119
rect 506208 398349 506328 399059
rect 506208 398315 506251 398349
rect 506285 398315 506328 398349
rect 506208 398149 506328 398315
rect 506208 398115 506251 398149
rect 506285 398115 506328 398149
rect 504328 397915 504371 397949
rect 504405 397915 504448 397949
rect 504328 397749 504448 397915
rect 504328 397715 504371 397749
rect 504405 397715 504448 397749
rect 504328 397549 504448 397715
rect 504328 397515 504371 397549
rect 504405 397515 504448 397549
rect 504328 397349 504448 397515
rect 504328 397315 504371 397349
rect 504405 397315 504448 397349
rect 504328 397149 504448 397315
rect 504328 397115 504371 397149
rect 504405 397115 504448 397149
rect 504328 396949 504448 397115
rect 504328 396915 504371 396949
rect 504405 396915 504448 396949
rect 504328 396749 504448 396915
rect 504328 396715 504371 396749
rect 504405 396715 504448 396749
rect 504328 396549 504448 396715
rect 504328 396515 504371 396549
rect 504405 396515 504448 396549
rect 506208 397949 506328 398115
rect 506208 397915 506251 397949
rect 506285 397915 506328 397949
rect 506208 397749 506328 397915
rect 506208 397715 506251 397749
rect 506285 397715 506328 397749
rect 506208 397549 506328 397715
rect 506208 397515 506251 397549
rect 506285 397515 506328 397549
rect 506208 397349 506328 397515
rect 506208 397315 506251 397349
rect 506285 397315 506328 397349
rect 506208 397149 506328 397315
rect 506208 397115 506251 397149
rect 506285 397115 506328 397149
rect 506208 396949 506328 397115
rect 506208 396915 506251 396949
rect 506285 396915 506328 396949
rect 506208 396749 506328 396915
rect 506208 396715 506251 396749
rect 506285 396715 506328 396749
rect 506208 396549 506328 396715
rect 504328 396349 504448 396515
rect 505189 396513 506153 396524
rect 504328 396315 504371 396349
rect 504405 396315 504448 396349
rect 504328 395603 504448 396315
rect 504627 396506 506153 396513
rect 504627 396112 504639 396506
rect 505177 396112 505599 396506
rect 506137 396112 506153 396506
rect 504627 396103 506153 396112
rect 505189 396092 506153 396103
rect 506208 396515 506251 396549
rect 506285 396515 506328 396549
rect 506208 396349 506328 396515
rect 506208 396315 506251 396349
rect 506285 396315 506328 396349
rect 504328 395569 504371 395603
rect 504405 395569 504448 395603
rect 504328 395403 504448 395569
rect 504328 395369 504371 395403
rect 504405 395369 504448 395403
rect 504328 395203 504448 395369
rect 504627 395768 505189 395776
rect 504627 395374 504639 395768
rect 505177 395374 505189 395768
rect 504627 395366 505189 395374
rect 505587 395768 506149 395776
rect 505587 395374 505599 395768
rect 506137 395694 506149 395768
rect 506208 395694 506328 396315
rect 506137 395666 506328 395694
rect 506137 395374 506149 395666
rect 505587 395366 506149 395374
rect 506208 395603 506328 395666
rect 506208 395569 506251 395603
rect 506285 395569 506328 395603
rect 506208 395403 506328 395569
rect 506208 395369 506251 395403
rect 506285 395369 506328 395403
rect 504328 395169 504371 395203
rect 504405 395169 504448 395203
rect 504328 395003 504448 395169
rect 504328 394969 504371 395003
rect 504405 394969 504448 395003
rect 504328 394803 504448 394969
rect 504328 394769 504371 394803
rect 504405 394769 504448 394803
rect 504328 394603 504448 394769
rect 504328 394569 504371 394603
rect 504405 394569 504448 394603
rect 504328 394403 504448 394569
rect 504328 394369 504371 394403
rect 504405 394369 504448 394403
rect 504328 394203 504448 394369
rect 504328 394169 504371 394203
rect 504405 394169 504448 394203
rect 504328 394003 504448 394169
rect 504328 393969 504371 394003
rect 504405 393969 504448 394003
rect 504328 393803 504448 393969
rect 504328 393769 504371 393803
rect 504405 393769 504448 393803
rect 504328 393603 504448 393769
rect 504328 393569 504371 393603
rect 504405 393569 504448 393603
rect 504328 393403 504448 393569
rect 504328 393369 504371 393403
rect 504405 393369 504448 393403
rect 504328 393203 504448 393369
rect 504680 393302 504708 395366
rect 504328 393169 504371 393203
rect 504405 393169 504448 393203
rect 504328 393003 504448 393169
rect 504328 392969 504371 393003
rect 504405 392969 504448 393003
rect 504328 392273 504448 392969
rect 504544 393274 504708 393302
rect 506208 395203 506328 395369
rect 506208 395169 506251 395203
rect 506285 395169 506328 395203
rect 506208 395003 506328 395169
rect 506208 394969 506251 395003
rect 506285 394969 506328 395003
rect 506208 394803 506328 394969
rect 506208 394769 506251 394803
rect 506285 394769 506328 394803
rect 506208 394603 506328 394769
rect 506208 394569 506251 394603
rect 506285 394569 506328 394603
rect 506208 394403 506328 394569
rect 506208 394369 506251 394403
rect 506285 394369 506328 394403
rect 506208 394203 506328 394369
rect 506208 394169 506251 394203
rect 506285 394169 506328 394203
rect 506208 394003 506328 394169
rect 506208 393969 506251 394003
rect 506285 393969 506328 394003
rect 506208 393803 506328 393969
rect 506208 393769 506251 393803
rect 506285 393769 506328 393803
rect 506208 393603 506328 393769
rect 506208 393569 506251 393603
rect 506285 393569 506328 393603
rect 506208 393403 506328 393569
rect 506208 393369 506251 393403
rect 506285 393369 506328 393403
rect 504544 392676 504572 393274
rect 505189 393194 506153 393205
rect 504627 393187 506153 393194
rect 504627 392793 504639 393187
rect 505177 392793 505599 393187
rect 506137 392793 506153 393187
rect 504627 392784 506153 392793
rect 505189 392773 506153 392784
rect 506208 393203 506328 393369
rect 506208 393169 506251 393203
rect 506285 393169 506328 393203
rect 506208 393003 506328 393169
rect 506208 392969 506251 393003
rect 506285 392969 506328 393003
rect 504532 392670 504584 392676
rect 504532 392612 504584 392618
rect 505620 392670 505672 392676
rect 505620 392612 505672 392618
rect 505144 392578 505196 392584
rect 505144 392520 505196 392526
rect 505156 392445 505184 392520
rect 505632 392445 505660 392612
rect 504328 392239 504371 392273
rect 504405 392239 504448 392273
rect 504328 392073 504448 392239
rect 504328 392039 504371 392073
rect 504405 392039 504448 392073
rect 504328 391873 504448 392039
rect 504627 392437 505189 392445
rect 504627 392043 504639 392437
rect 505177 392043 505189 392437
rect 504627 392035 505189 392043
rect 505587 392437 506149 392445
rect 505587 392043 505599 392437
rect 506137 392043 506149 392437
rect 505587 392035 506149 392043
rect 506208 392273 506328 392969
rect 506208 392239 506251 392273
rect 506285 392239 506328 392273
rect 506208 392073 506328 392239
rect 506208 392039 506251 392073
rect 506285 392039 506328 392073
rect 504328 391839 504371 391873
rect 504405 391839 504448 391873
rect 504328 391673 504448 391839
rect 504328 391639 504371 391673
rect 504405 391639 504448 391673
rect 504328 391473 504448 391639
rect 504328 391439 504371 391473
rect 504405 391439 504448 391473
rect 504328 391273 504448 391439
rect 504328 391239 504371 391273
rect 504405 391239 504448 391273
rect 504328 391073 504448 391239
rect 504328 391039 504371 391073
rect 504405 391039 504448 391073
rect 504328 390873 504448 391039
rect 504328 390839 504371 390873
rect 504405 390839 504448 390873
rect 504328 390673 504448 390839
rect 504328 390639 504371 390673
rect 504405 390639 504448 390673
rect 504328 390473 504448 390639
rect 504328 390439 504371 390473
rect 504405 390439 504448 390473
rect 506208 391873 506328 392039
rect 506208 391839 506251 391873
rect 506285 391839 506328 391873
rect 506208 391673 506328 391839
rect 506208 391639 506251 391673
rect 506285 391639 506328 391673
rect 506208 391473 506328 391639
rect 506208 391439 506251 391473
rect 506285 391439 506328 391473
rect 506208 391273 506328 391439
rect 506208 391239 506251 391273
rect 506285 391239 506328 391273
rect 506208 391073 506328 391239
rect 506208 391039 506251 391073
rect 506285 391039 506328 391073
rect 506208 390873 506328 391039
rect 506208 390839 506251 390873
rect 506285 390839 506328 390873
rect 506208 390673 506328 390839
rect 506208 390639 506251 390673
rect 506285 390639 506328 390673
rect 506208 390473 506328 390639
rect 504328 390273 504448 390439
rect 505189 390437 506153 390448
rect 504328 390239 504371 390273
rect 504405 390239 504448 390273
rect 504328 389353 504448 390239
rect 504627 390430 506153 390437
rect 504627 390036 504639 390430
rect 505177 390036 505599 390430
rect 506137 390036 506153 390430
rect 504627 390027 506153 390036
rect 505189 390016 506153 390027
rect 506208 390439 506251 390473
rect 506285 390439 506328 390473
rect 506208 390273 506328 390439
rect 506208 390239 506251 390273
rect 506285 390239 506328 390273
rect 504868 389524 505668 389530
rect 504868 389490 504891 389524
rect 504925 389490 504963 389524
rect 504997 389490 505035 389524
rect 505069 389490 505107 389524
rect 505141 389490 505179 389524
rect 505213 389490 505251 389524
rect 505285 389490 505323 389524
rect 505357 389490 505395 389524
rect 505429 389490 505467 389524
rect 505501 389490 505539 389524
rect 505573 389490 505611 389524
rect 505645 389490 505668 389524
rect 504868 389484 505668 389490
rect 504328 389319 504371 389353
rect 504405 389319 504448 389353
rect 503988 389174 504040 389180
rect 503988 389116 504040 389122
rect 502448 388863 502491 388897
rect 502525 388863 502568 388897
rect 502448 388497 502568 388863
rect 502448 388463 502491 388497
rect 502525 388463 502568 388497
rect 502448 388097 502568 388463
rect 502448 388063 502491 388097
rect 502525 388063 502568 388097
rect 502448 387697 502568 388063
rect 502448 387663 502491 387697
rect 502525 387663 502568 387697
rect 502448 387297 502568 387663
rect 502448 387263 502491 387297
rect 502525 387263 502568 387297
rect 502232 387018 502328 387046
rect 500568 386863 500611 386897
rect 500645 386863 500688 386897
rect 502232 386880 502260 386935
rect 500568 385433 500688 386863
rect 502220 386874 502272 386880
rect 502220 386816 502272 386822
rect 502300 386788 502328 387018
rect 502448 386897 502568 387263
rect 502448 386863 502491 386897
rect 502525 386863 502568 386897
rect 502288 386782 502340 386788
rect 500863 386737 502153 386743
rect 500863 386703 500879 386737
rect 500913 386703 500951 386737
rect 500985 386703 501023 386737
rect 501057 386703 501095 386737
rect 501129 386703 501167 386737
rect 501201 386703 501239 386737
rect 501273 386703 501311 386737
rect 501345 386703 501383 386737
rect 501417 386703 501455 386737
rect 501489 386703 501527 386737
rect 501561 386703 501599 386737
rect 501633 386703 501671 386737
rect 501705 386703 501743 386737
rect 501777 386703 501815 386737
rect 501849 386703 501887 386737
rect 501921 386703 501959 386737
rect 501993 386703 502031 386737
rect 502065 386703 502103 386737
rect 502137 386703 502153 386737
rect 502288 386724 502340 386730
rect 500863 386697 502153 386703
rect 502359 386681 502405 386693
rect 502359 386678 502365 386681
rect 502300 386650 502365 386678
rect 502084 386598 502136 386604
rect 502084 386540 502136 386546
rect 502096 385575 502124 386540
rect 500863 385569 502153 385575
rect 500863 385535 500879 385569
rect 500913 385535 500951 385569
rect 500985 385535 501023 385569
rect 501057 385535 501095 385569
rect 501129 385535 501167 385569
rect 501201 385535 501239 385569
rect 501273 385535 501311 385569
rect 501345 385535 501383 385569
rect 501417 385535 501455 385569
rect 501489 385535 501527 385569
rect 501561 385535 501599 385569
rect 501633 385535 501671 385569
rect 501705 385535 501743 385569
rect 501777 385535 501815 385569
rect 501849 385535 501887 385569
rect 501921 385535 501959 385569
rect 501993 385535 502031 385569
rect 502065 385535 502103 385569
rect 502137 385535 502153 385569
rect 500863 385529 502153 385535
rect 502300 385482 502328 386650
rect 502359 386647 502365 386650
rect 502399 386647 502405 386681
rect 502359 386635 502405 386647
rect 502368 385500 502396 385555
rect 500568 385399 500611 385433
rect 500645 385399 500688 385433
rect 500568 385033 500688 385399
rect 502096 385454 502328 385482
rect 502356 385494 502408 385500
rect 502096 385117 502124 385454
rect 502356 385436 502408 385442
rect 502448 385433 502568 386863
rect 502448 385399 502491 385433
rect 502525 385399 502568 385433
rect 500863 385111 502153 385117
rect 500863 385077 500879 385111
rect 500913 385077 500951 385111
rect 500985 385077 501023 385111
rect 501057 385077 501095 385111
rect 501129 385077 501167 385111
rect 501201 385077 501239 385111
rect 501273 385077 501311 385111
rect 501345 385077 501383 385111
rect 501417 385077 501455 385111
rect 501489 385077 501527 385111
rect 501561 385077 501599 385111
rect 501633 385077 501671 385111
rect 501705 385077 501743 385111
rect 501777 385077 501815 385111
rect 501849 385077 501887 385111
rect 501921 385077 501959 385111
rect 501993 385077 502031 385111
rect 502065 385077 502103 385111
rect 502137 385077 502153 385111
rect 500863 385071 502153 385077
rect 500568 384999 500611 385033
rect 500645 384999 500688 385033
rect 500568 384633 500688 384999
rect 502448 385033 502568 385399
rect 502448 384999 502491 385033
rect 502525 384999 502568 385033
rect 500568 384599 500611 384633
rect 500645 384599 500688 384633
rect 500863 384653 502153 384659
rect 500863 384619 500879 384653
rect 500913 384619 500951 384653
rect 500985 384619 501023 384653
rect 501057 384619 501095 384653
rect 501129 384619 501167 384653
rect 501201 384619 501239 384653
rect 501273 384619 501311 384653
rect 501345 384619 501383 384653
rect 501417 384619 501455 384653
rect 501489 384619 501527 384653
rect 501561 384619 501599 384653
rect 501633 384619 501671 384653
rect 501705 384619 501743 384653
rect 501777 384619 501815 384653
rect 501849 384619 501887 384653
rect 501921 384619 501959 384653
rect 501993 384619 502031 384653
rect 502065 384619 502103 384653
rect 502137 384619 502153 384653
rect 500863 384613 502153 384619
rect 502448 384633 502568 384999
rect 500568 384233 500688 384599
rect 500568 384199 500611 384233
rect 500645 384199 500688 384233
rect 502448 384599 502491 384633
rect 502525 384599 502568 384633
rect 502448 384233 502568 384599
rect 500568 383833 500688 384199
rect 500863 384195 502153 384201
rect 500863 384161 500879 384195
rect 500913 384161 500951 384195
rect 500985 384161 501023 384195
rect 501057 384161 501095 384195
rect 501129 384161 501167 384195
rect 501201 384161 501239 384195
rect 501273 384161 501311 384195
rect 501345 384161 501383 384195
rect 501417 384161 501455 384195
rect 501489 384161 501527 384195
rect 501561 384161 501599 384195
rect 501633 384161 501671 384195
rect 501705 384161 501743 384195
rect 501777 384161 501815 384195
rect 501849 384161 501887 384195
rect 501921 384161 501959 384195
rect 501993 384161 502031 384195
rect 502065 384161 502103 384195
rect 502137 384161 502153 384195
rect 500863 384155 502153 384161
rect 502448 384199 502491 384233
rect 502525 384199 502568 384233
rect 500568 383799 500611 383833
rect 500645 383799 500688 383833
rect 500568 383433 500688 383799
rect 502448 383833 502568 384199
rect 502448 383799 502491 383833
rect 502525 383799 502568 383833
rect 500863 383737 502153 383743
rect 500863 383703 500879 383737
rect 500913 383703 500951 383737
rect 500985 383703 501023 383737
rect 501057 383703 501095 383737
rect 501129 383703 501167 383737
rect 501201 383703 501239 383737
rect 501273 383703 501311 383737
rect 501345 383703 501383 383737
rect 501417 383703 501455 383737
rect 501489 383703 501527 383737
rect 501561 383703 501599 383737
rect 501633 383703 501671 383737
rect 501705 383703 501743 383737
rect 501777 383703 501815 383737
rect 501849 383703 501887 383737
rect 501921 383703 501959 383737
rect 501993 383703 502031 383737
rect 502065 383703 502103 383737
rect 502137 383703 502153 383737
rect 500863 383697 502153 383703
rect 500568 383399 500611 383433
rect 500645 383399 500688 383433
rect 500568 383033 500688 383399
rect 502448 383433 502568 383799
rect 502448 383399 502491 383433
rect 502525 383399 502568 383433
rect 500863 383279 502153 383285
rect 500863 383245 500879 383279
rect 500913 383245 500951 383279
rect 500985 383245 501023 383279
rect 501057 383245 501095 383279
rect 501129 383245 501167 383279
rect 501201 383245 501239 383279
rect 501273 383245 501311 383279
rect 501345 383245 501383 383279
rect 501417 383245 501455 383279
rect 501489 383245 501527 383279
rect 501561 383245 501599 383279
rect 501633 383245 501671 383279
rect 501705 383245 501743 383279
rect 501777 383245 501815 383279
rect 501849 383245 501887 383279
rect 501921 383245 501959 383279
rect 501993 383245 502031 383279
rect 502065 383245 502103 383279
rect 502137 383245 502153 383279
rect 500863 383239 502153 383245
rect 500568 382999 500611 383033
rect 500645 382999 500688 383033
rect 500568 382633 500688 382999
rect 502448 383033 502568 383399
rect 502448 382999 502491 383033
rect 502525 382999 502568 383033
rect 500863 382821 502153 382827
rect 500863 382787 500879 382821
rect 500913 382787 500951 382821
rect 500985 382787 501023 382821
rect 501057 382787 501095 382821
rect 501129 382787 501167 382821
rect 501201 382787 501239 382821
rect 501273 382787 501311 382821
rect 501345 382787 501383 382821
rect 501417 382787 501455 382821
rect 501489 382787 501527 382821
rect 501561 382787 501599 382821
rect 501633 382787 501671 382821
rect 501705 382787 501743 382821
rect 501777 382787 501815 382821
rect 501849 382787 501887 382821
rect 501921 382787 501959 382821
rect 501993 382787 502031 382821
rect 502065 382787 502103 382821
rect 502137 382787 502153 382821
rect 500863 382781 502153 382787
rect 500568 382599 500611 382633
rect 500645 382599 500688 382633
rect 500568 382354 500688 382599
rect 502448 382633 502568 382999
rect 502448 382599 502491 382633
rect 502525 382599 502568 382633
rect 500863 382363 502153 382369
rect 500863 382354 500879 382363
rect 500568 382329 500879 382354
rect 500913 382329 500951 382363
rect 500985 382329 501023 382363
rect 501057 382329 501095 382363
rect 501129 382329 501167 382363
rect 501201 382329 501239 382363
rect 501273 382329 501311 382363
rect 501345 382329 501383 382363
rect 501417 382329 501455 382363
rect 501489 382329 501527 382363
rect 501561 382329 501599 382363
rect 501633 382329 501671 382363
rect 501705 382329 501743 382363
rect 501777 382329 501815 382363
rect 501849 382329 501887 382363
rect 501921 382329 501959 382363
rect 501993 382329 502031 382363
rect 502065 382329 502103 382363
rect 502137 382329 502153 382363
rect 500568 382326 502153 382329
rect 500568 382233 500688 382326
rect 500863 382323 502153 382326
rect 500568 382199 500611 382233
rect 500645 382199 500688 382233
rect 500568 381833 500688 382199
rect 502448 382233 502568 382599
rect 502448 382199 502491 382233
rect 502525 382199 502568 382233
rect 500863 381905 502153 381911
rect 500863 381871 500879 381905
rect 500913 381871 500951 381905
rect 500985 381871 501023 381905
rect 501057 381871 501095 381905
rect 501129 381871 501167 381905
rect 501201 381871 501239 381905
rect 501273 381871 501311 381905
rect 501345 381871 501383 381905
rect 501417 381871 501455 381905
rect 501489 381871 501527 381905
rect 501561 381871 501599 381905
rect 501633 381871 501671 381905
rect 501705 381871 501743 381905
rect 501777 381871 501815 381905
rect 501849 381871 501887 381905
rect 501921 381871 501959 381905
rect 501993 381871 502031 381905
rect 502065 381871 502103 381905
rect 502137 381871 502153 381905
rect 500863 381865 502153 381871
rect 500568 381799 500611 381833
rect 500645 381799 500688 381833
rect 500568 381433 500688 381799
rect 502448 381833 502568 382199
rect 502448 381799 502491 381833
rect 502525 381799 502568 381833
rect 500568 381399 500611 381433
rect 500645 381399 500688 381433
rect 500863 381447 502153 381453
rect 500863 381413 500879 381447
rect 500913 381413 500951 381447
rect 500985 381413 501023 381447
rect 501057 381413 501095 381447
rect 501129 381413 501167 381447
rect 501201 381413 501239 381447
rect 501273 381413 501311 381447
rect 501345 381413 501383 381447
rect 501417 381413 501455 381447
rect 501489 381413 501527 381447
rect 501561 381413 501599 381447
rect 501633 381413 501671 381447
rect 501705 381413 501743 381447
rect 501777 381413 501815 381447
rect 501849 381413 501887 381447
rect 501921 381413 501959 381447
rect 501993 381413 502031 381447
rect 502065 381413 502103 381447
rect 502137 381413 502153 381447
rect 500863 381407 502153 381413
rect 502448 381433 502568 381799
rect 500568 381033 500688 381399
rect 500568 380999 500611 381033
rect 500645 380999 500688 381033
rect 500568 380633 500688 380999
rect 502448 381399 502491 381433
rect 502525 381399 502568 381433
rect 502448 381033 502568 381399
rect 502448 380999 502491 381033
rect 502525 380999 502568 381033
rect 500863 380989 502153 380995
rect 500863 380955 500879 380989
rect 500913 380955 500951 380989
rect 500985 380955 501023 380989
rect 501057 380955 501095 380989
rect 501129 380955 501167 380989
rect 501201 380955 501239 380989
rect 501273 380955 501311 380989
rect 501345 380955 501383 380989
rect 501417 380955 501455 380989
rect 501489 380955 501527 380989
rect 501561 380955 501599 380989
rect 501633 380955 501671 380989
rect 501705 380955 501743 380989
rect 501777 380955 501815 380989
rect 501849 380955 501887 380989
rect 501921 380955 501959 380989
rect 501993 380955 502031 380989
rect 502065 380955 502103 380989
rect 502137 380955 502153 380989
rect 500863 380949 502153 380955
rect 500568 380599 500611 380633
rect 500645 380599 500688 380633
rect 500568 380233 500688 380599
rect 502448 380633 502568 380999
rect 502448 380599 502491 380633
rect 502525 380599 502568 380633
rect 500863 380531 502153 380537
rect 500863 380497 500879 380531
rect 500913 380497 500951 380531
rect 500985 380497 501023 380531
rect 501057 380497 501095 380531
rect 501129 380497 501167 380531
rect 501201 380497 501239 380531
rect 501273 380497 501311 380531
rect 501345 380497 501383 380531
rect 501417 380497 501455 380531
rect 501489 380497 501527 380531
rect 501561 380497 501599 380531
rect 501633 380497 501671 380531
rect 501705 380497 501743 380531
rect 501777 380497 501815 380531
rect 501849 380497 501887 380531
rect 501921 380497 501959 380531
rect 501993 380497 502031 380531
rect 502065 380497 502103 380531
rect 502137 380497 502153 380531
rect 500863 380491 502153 380497
rect 500568 380199 500611 380233
rect 500645 380199 500688 380233
rect 500568 377495 500688 380199
rect 502448 380233 502568 380599
rect 504328 388953 504448 389319
rect 506208 389353 506328 390239
rect 506208 389319 506251 389353
rect 506285 389319 506328 389353
rect 504872 389174 504924 389180
rect 504872 389116 504924 389122
rect 504884 389072 504912 389116
rect 504868 389066 505668 389072
rect 504868 389032 504891 389066
rect 504925 389032 504963 389066
rect 504997 389032 505035 389066
rect 505069 389032 505107 389066
rect 505141 389032 505179 389066
rect 505213 389032 505251 389066
rect 505285 389032 505323 389066
rect 505357 389032 505395 389066
rect 505429 389032 505467 389066
rect 505501 389032 505539 389066
rect 505573 389032 505611 389066
rect 505645 389032 505668 389066
rect 504868 389026 505668 389032
rect 504328 388919 504371 388953
rect 504405 388919 504448 388953
rect 504328 388553 504448 388919
rect 506208 388953 506328 389319
rect 506208 388919 506251 388953
rect 506285 388919 506328 388953
rect 504868 388608 505668 388614
rect 504868 388574 504891 388608
rect 504925 388574 504963 388608
rect 504997 388574 505035 388608
rect 505069 388574 505107 388608
rect 505141 388574 505179 388608
rect 505213 388574 505251 388608
rect 505285 388574 505323 388608
rect 505357 388574 505395 388608
rect 505429 388574 505467 388608
rect 505501 388574 505539 388608
rect 505573 388574 505611 388608
rect 505645 388574 505668 388608
rect 504868 388568 505668 388574
rect 504328 388519 504371 388553
rect 504405 388519 504448 388553
rect 504328 388153 504448 388519
rect 506208 388553 506328 388919
rect 506208 388519 506251 388553
rect 506285 388519 506328 388553
rect 504328 388119 504371 388153
rect 504405 388119 504448 388153
rect 504328 387753 504448 388119
rect 504868 388150 505668 388156
rect 504868 388116 504891 388150
rect 504925 388116 504963 388150
rect 504997 388116 505035 388150
rect 505069 388116 505107 388150
rect 505141 388116 505179 388150
rect 505213 388116 505251 388150
rect 505285 388116 505323 388150
rect 505357 388116 505395 388150
rect 505429 388116 505467 388150
rect 505501 388116 505539 388150
rect 505573 388116 505611 388150
rect 505645 388116 505668 388150
rect 504868 388110 505668 388116
rect 506208 388153 506328 388519
rect 506208 388119 506251 388153
rect 506285 388119 506328 388153
rect 504328 387719 504371 387753
rect 504405 387719 504448 387753
rect 504328 387353 504448 387719
rect 506208 387753 506328 388119
rect 506208 387719 506251 387753
rect 506285 387719 506328 387753
rect 504868 387692 505668 387698
rect 504868 387658 504891 387692
rect 504925 387658 504963 387692
rect 504997 387658 505035 387692
rect 505069 387658 505107 387692
rect 505141 387658 505179 387692
rect 505213 387658 505251 387692
rect 505285 387658 505323 387692
rect 505357 387658 505395 387692
rect 505429 387658 505467 387692
rect 505501 387658 505539 387692
rect 505573 387658 505611 387692
rect 505645 387658 505668 387692
rect 504868 387652 505668 387658
rect 504328 387319 504371 387353
rect 504405 387319 504448 387353
rect 504328 386953 504448 387319
rect 506208 387353 506328 387719
rect 506208 387319 506251 387353
rect 506285 387319 506328 387353
rect 504868 387234 505668 387240
rect 504868 387200 504891 387234
rect 504925 387200 504963 387234
rect 504997 387200 505035 387234
rect 505069 387200 505107 387234
rect 505141 387200 505179 387234
rect 505213 387200 505251 387234
rect 505285 387200 505323 387234
rect 505357 387200 505395 387234
rect 505429 387200 505467 387234
rect 505501 387200 505539 387234
rect 505573 387200 505611 387234
rect 505645 387200 505668 387234
rect 504868 387194 505668 387200
rect 504328 386919 504371 386953
rect 504405 386919 504448 386953
rect 506208 386953 506328 387319
rect 504328 386553 504448 386919
rect 505904 386880 505932 386935
rect 506208 386919 506251 386953
rect 506285 386919 506328 386953
rect 505892 386874 505944 386880
rect 505892 386816 505944 386822
rect 504868 386776 505668 386782
rect 504868 386742 504891 386776
rect 504925 386742 504963 386776
rect 504997 386742 505035 386776
rect 505069 386742 505107 386776
rect 505141 386742 505179 386776
rect 505213 386742 505251 386776
rect 505285 386742 505323 386776
rect 505357 386742 505395 386776
rect 505429 386742 505467 386776
rect 505501 386742 505539 386776
rect 505573 386742 505611 386776
rect 505645 386742 505668 386776
rect 504868 386736 505668 386742
rect 504328 386519 504371 386553
rect 504405 386519 504448 386553
rect 504328 386153 504448 386519
rect 506208 386553 506328 386919
rect 506208 386519 506251 386553
rect 506285 386519 506328 386553
rect 504868 386318 505668 386324
rect 504868 386284 504891 386318
rect 504925 386284 504963 386318
rect 504997 386284 505035 386318
rect 505069 386284 505107 386318
rect 505141 386284 505179 386318
rect 505213 386284 505251 386318
rect 505285 386284 505323 386318
rect 505357 386284 505395 386318
rect 505429 386284 505467 386318
rect 505501 386284 505539 386318
rect 505573 386284 505611 386318
rect 505645 386284 505668 386318
rect 504868 386278 505668 386284
rect 504328 386119 504371 386153
rect 504405 386119 504448 386153
rect 504328 385753 504448 386119
rect 506208 386153 506328 386519
rect 506208 386119 506251 386153
rect 506285 386119 506328 386153
rect 504868 385860 505668 385866
rect 504868 385826 504891 385860
rect 504925 385826 504963 385860
rect 504997 385826 505035 385860
rect 505069 385826 505107 385860
rect 505141 385826 505179 385860
rect 505213 385826 505251 385860
rect 505285 385826 505323 385860
rect 505357 385826 505395 385860
rect 505429 385826 505467 385860
rect 505501 385826 505539 385860
rect 505573 385826 505611 385860
rect 505645 385826 505668 385860
rect 504868 385820 505668 385826
rect 504328 385719 504371 385753
rect 504405 385719 504448 385753
rect 504328 384843 504448 385719
rect 505088 385500 505116 385820
rect 506208 385753 506328 386119
rect 506208 385719 506251 385753
rect 506285 385719 506328 385753
rect 505076 385494 505128 385500
rect 505076 385436 505128 385442
rect 504868 385402 505668 385408
rect 504868 385368 504891 385402
rect 504925 385368 504963 385402
rect 504997 385368 505035 385402
rect 505069 385368 505107 385402
rect 505141 385368 505179 385402
rect 505213 385368 505251 385402
rect 505285 385368 505323 385402
rect 505357 385368 505395 385402
rect 505429 385368 505467 385402
rect 505501 385368 505539 385402
rect 505573 385368 505611 385402
rect 505645 385368 505668 385402
rect 504868 385362 505668 385368
rect 504328 384809 504371 384843
rect 504405 384809 504448 384843
rect 504328 384443 504448 384809
rect 504328 384409 504371 384443
rect 504405 384409 504448 384443
rect 504328 384043 504448 384409
rect 504328 384009 504371 384043
rect 504405 384009 504448 384043
rect 504328 383643 504448 384009
rect 504328 383609 504371 383643
rect 504405 383609 504448 383643
rect 504328 383243 504448 383609
rect 504328 383209 504371 383243
rect 504405 383209 504448 383243
rect 504328 382843 504448 383209
rect 504328 382809 504371 382843
rect 504405 382809 504448 382843
rect 504328 382443 504448 382809
rect 504328 382409 504371 382443
rect 504405 382409 504448 382443
rect 504328 382043 504448 382409
rect 504328 382009 504371 382043
rect 504405 382009 504448 382043
rect 504328 381643 504448 382009
rect 504328 381609 504371 381643
rect 504405 381609 504448 381643
rect 504328 381538 504448 381609
rect 504328 381486 504396 381538
rect 504328 381243 504448 381486
rect 504328 381209 504371 381243
rect 504405 381209 504448 381243
rect 504328 380843 504448 381209
rect 504328 380809 504371 380843
rect 504405 380809 504448 380843
rect 504056 380526 504108 380532
rect 504056 380468 504108 380474
rect 502448 380199 502491 380233
rect 502525 380199 502568 380233
rect 500863 380073 502153 380079
rect 500863 380039 500879 380073
rect 500913 380039 500951 380073
rect 500985 380039 501023 380073
rect 501057 380039 501095 380073
rect 501129 380039 501167 380073
rect 501201 380039 501239 380073
rect 501273 380039 501311 380073
rect 501345 380039 501383 380073
rect 501417 380039 501455 380073
rect 501489 380039 501527 380073
rect 501561 380039 501599 380073
rect 501633 380039 501671 380073
rect 501705 380039 501743 380073
rect 501777 380039 501815 380073
rect 501849 380039 501887 380073
rect 501921 380039 501959 380073
rect 501993 380039 502031 380073
rect 502065 380039 502103 380073
rect 502137 380039 502153 380073
rect 500863 380033 502153 380039
rect 501948 379146 502000 379152
rect 501948 379088 502000 379094
rect 501108 377666 501908 377672
rect 501108 377632 501131 377666
rect 501165 377632 501203 377666
rect 501237 377632 501275 377666
rect 501309 377632 501347 377666
rect 501381 377632 501419 377666
rect 501453 377632 501491 377666
rect 501525 377632 501563 377666
rect 501597 377632 501635 377666
rect 501669 377632 501707 377666
rect 501741 377632 501779 377666
rect 501813 377632 501851 377666
rect 501885 377632 501908 377666
rect 501108 377626 501908 377632
rect 500568 377461 500611 377495
rect 500645 377461 500688 377495
rect 500568 377095 500688 377461
rect 501108 377208 501908 377214
rect 501108 377174 501131 377208
rect 501165 377174 501203 377208
rect 501237 377174 501275 377208
rect 501309 377174 501347 377208
rect 501381 377174 501419 377208
rect 501453 377174 501491 377208
rect 501525 377174 501563 377208
rect 501597 377174 501635 377208
rect 501669 377174 501707 377208
rect 501741 377174 501779 377208
rect 501813 377174 501851 377208
rect 501885 377202 501908 377208
rect 501960 377202 501988 379088
rect 501885 377174 501988 377202
rect 502448 377495 502568 380199
rect 504068 379152 504096 380468
rect 504328 380443 504448 380809
rect 504884 380532 504912 385362
rect 506208 384843 506328 385719
rect 506208 384809 506251 384843
rect 506285 384809 506328 384843
rect 506208 384443 506328 384809
rect 506208 384409 506251 384443
rect 506285 384409 506328 384443
rect 506208 384043 506328 384409
rect 506208 384009 506251 384043
rect 506285 384009 506328 384043
rect 506208 383643 506328 384009
rect 506208 383609 506251 383643
rect 506285 383609 506328 383643
rect 506208 383243 506328 383609
rect 506208 383209 506251 383243
rect 506285 383209 506328 383243
rect 506208 382843 506328 383209
rect 506208 382809 506251 382843
rect 506285 382809 506328 382843
rect 506208 382443 506328 382809
rect 506208 382409 506251 382443
rect 506285 382409 506328 382443
rect 506208 382043 506328 382409
rect 506208 382009 506251 382043
rect 506285 382009 506328 382043
rect 506208 381643 506328 382009
rect 506208 381609 506251 381643
rect 506285 381609 506328 381643
rect 506208 381243 506328 381609
rect 506208 381209 506251 381243
rect 506285 381209 506328 381243
rect 506208 380843 506328 381209
rect 506208 380809 506251 380843
rect 506285 380809 506328 380843
rect 504872 380526 504924 380532
rect 504872 380468 504924 380474
rect 504328 380409 504371 380443
rect 504405 380409 504448 380443
rect 504328 380043 504448 380409
rect 504328 380009 504371 380043
rect 504405 380009 504448 380043
rect 504328 379643 504448 380009
rect 504328 379609 504371 379643
rect 504405 379609 504448 379643
rect 504328 379243 504448 379609
rect 504328 379209 504371 379243
rect 504405 379209 504448 379243
rect 504056 379146 504108 379152
rect 504056 379088 504108 379094
rect 502448 377461 502491 377495
rect 502525 377461 502568 377495
rect 501108 377168 501908 377174
rect 500568 377061 500611 377095
rect 500645 377061 500688 377095
rect 500568 376695 500688 377061
rect 502448 377095 502568 377461
rect 502448 377061 502491 377095
rect 502525 377061 502568 377095
rect 501108 376750 501908 376756
rect 501108 376716 501131 376750
rect 501165 376716 501203 376750
rect 501237 376716 501275 376750
rect 501309 376716 501347 376750
rect 501381 376716 501419 376750
rect 501453 376716 501491 376750
rect 501525 376716 501563 376750
rect 501597 376716 501635 376750
rect 501669 376716 501707 376750
rect 501741 376716 501779 376750
rect 501813 376716 501851 376750
rect 501885 376716 501908 376750
rect 501108 376710 501908 376716
rect 500568 376661 500611 376695
rect 500645 376661 500688 376695
rect 500568 376295 500688 376661
rect 501824 376392 501852 376710
rect 502448 376695 502568 377061
rect 502448 376661 502491 376695
rect 502525 376661 502568 376695
rect 501812 376386 501864 376392
rect 501812 376328 501864 376334
rect 500568 376261 500611 376295
rect 500645 376261 500688 376295
rect 500568 375895 500688 376261
rect 501108 376292 501908 376298
rect 501108 376258 501131 376292
rect 501165 376258 501203 376292
rect 501237 376258 501275 376292
rect 501309 376258 501347 376292
rect 501381 376258 501419 376292
rect 501453 376258 501491 376292
rect 501525 376258 501563 376292
rect 501597 376258 501635 376292
rect 501669 376258 501707 376292
rect 501741 376258 501779 376292
rect 501813 376258 501851 376292
rect 501885 376258 501908 376292
rect 501108 376252 501908 376258
rect 502448 376295 502568 376661
rect 502448 376261 502491 376295
rect 502525 376261 502568 376295
rect 500568 375861 500611 375895
rect 500645 375861 500688 375895
rect 500568 375495 500688 375861
rect 502448 375895 502568 376261
rect 502448 375861 502491 375895
rect 502525 375861 502568 375895
rect 501108 375834 501908 375840
rect 501108 375800 501131 375834
rect 501165 375800 501203 375834
rect 501237 375800 501275 375834
rect 501309 375800 501347 375834
rect 501381 375800 501419 375834
rect 501453 375800 501491 375834
rect 501525 375800 501563 375834
rect 501597 375800 501635 375834
rect 501669 375800 501707 375834
rect 501741 375800 501779 375834
rect 501813 375800 501851 375834
rect 501885 375800 501908 375834
rect 501108 375794 501908 375800
rect 500568 375461 500611 375495
rect 500645 375461 500688 375495
rect 500568 375095 500688 375461
rect 502448 375495 502568 375861
rect 502448 375461 502491 375495
rect 502525 375461 502568 375495
rect 501108 375376 501908 375382
rect 501108 375342 501131 375376
rect 501165 375342 501203 375376
rect 501237 375342 501275 375376
rect 501309 375342 501347 375376
rect 501381 375342 501419 375376
rect 501453 375342 501491 375376
rect 501525 375342 501563 375376
rect 501597 375342 501635 375376
rect 501669 375342 501707 375376
rect 501741 375342 501779 375376
rect 501813 375342 501851 375376
rect 501885 375342 501908 375376
rect 501108 375336 501908 375342
rect 500568 375061 500611 375095
rect 500645 375061 500688 375095
rect 500568 374695 500688 375061
rect 502448 375095 502568 375461
rect 502448 375061 502491 375095
rect 502525 375061 502568 375095
rect 501108 374918 501908 374924
rect 501108 374884 501131 374918
rect 501165 374884 501203 374918
rect 501237 374884 501275 374918
rect 501309 374884 501347 374918
rect 501381 374884 501419 374918
rect 501453 374884 501491 374918
rect 501525 374884 501563 374918
rect 501597 374884 501635 374918
rect 501669 374884 501707 374918
rect 501741 374884 501779 374918
rect 501813 374884 501851 374918
rect 501885 374884 501908 374918
rect 501108 374878 501908 374884
rect 500568 374661 500611 374695
rect 500645 374661 500688 374695
rect 500568 374295 500688 374661
rect 502448 374695 502568 375061
rect 502448 374661 502491 374695
rect 502525 374661 502568 374695
rect 501108 374460 501908 374466
rect 501108 374426 501131 374460
rect 501165 374426 501203 374460
rect 501237 374426 501275 374460
rect 501309 374426 501347 374460
rect 501381 374426 501419 374460
rect 501453 374426 501491 374460
rect 501525 374426 501563 374460
rect 501597 374426 501635 374460
rect 501669 374426 501707 374460
rect 501741 374426 501779 374460
rect 501813 374426 501851 374460
rect 501885 374426 501908 374460
rect 501108 374420 501908 374426
rect 500568 374261 500611 374295
rect 500645 374261 500688 374295
rect 500568 373895 500688 374261
rect 502448 374295 502568 374661
rect 502448 374261 502491 374295
rect 502525 374261 502568 374295
rect 501108 374002 501908 374008
rect 501108 373968 501131 374002
rect 501165 373968 501203 374002
rect 501237 373968 501275 374002
rect 501309 373968 501347 374002
rect 501381 373968 501419 374002
rect 501453 373968 501491 374002
rect 501525 373968 501563 374002
rect 501597 373968 501635 374002
rect 501669 373968 501707 374002
rect 501741 373968 501779 374002
rect 501813 373968 501851 374002
rect 501885 373968 501908 374002
rect 501108 373962 501908 373968
rect 500568 373861 500611 373895
rect 500645 373861 500688 373895
rect 500568 372987 500688 373861
rect 502448 373895 502568 374261
rect 502448 373861 502491 373895
rect 502525 373861 502568 373895
rect 501108 373544 501908 373550
rect 501108 373510 501131 373544
rect 501165 373510 501203 373544
rect 501237 373510 501275 373544
rect 501309 373510 501347 373544
rect 501381 373510 501419 373544
rect 501453 373510 501491 373544
rect 501525 373510 501563 373544
rect 501597 373510 501635 373544
rect 501669 373510 501707 373544
rect 501741 373510 501779 373544
rect 501813 373510 501851 373544
rect 501885 373510 501908 373544
rect 501108 373504 501908 373510
rect 502155 373525 502201 373537
rect 502155 373491 502161 373525
rect 502195 373491 502201 373525
rect 502155 373479 502201 373491
rect 500938 373124 501008 373144
rect 500938 373090 500944 373124
rect 500978 373090 501008 373124
rect 500938 373034 501008 373090
rect 500938 373000 500944 373034
rect 500978 373000 501008 373034
rect 500938 372988 501008 373000
rect 500568 372953 500611 372987
rect 500645 372953 500688 372987
rect 500568 372787 500688 372953
rect 500928 372982 501008 372988
rect 500980 372930 501008 372982
rect 501132 372982 501184 372988
rect 500928 372924 500944 372930
rect 500568 372753 500611 372787
rect 500645 372753 500688 372787
rect 500568 372587 500688 372753
rect 500568 372553 500611 372587
rect 500645 372553 500688 372587
rect 500568 372387 500688 372553
rect 500568 372353 500611 372387
rect 500645 372353 500688 372387
rect 500568 372187 500688 372353
rect 500568 372153 500611 372187
rect 500645 372153 500688 372187
rect 500568 371987 500688 372153
rect 500568 371953 500611 371987
rect 500645 371953 500688 371987
rect 500568 371787 500688 371953
rect 500568 371753 500611 371787
rect 500645 371753 500688 371787
rect 500568 371587 500688 371753
rect 500568 371553 500611 371587
rect 500645 371553 500688 371587
rect 500568 371387 500688 371553
rect 500568 371353 500611 371387
rect 500645 371353 500688 371387
rect 500568 371187 500688 371353
rect 500568 371153 500611 371187
rect 500645 371153 500688 371187
rect 500568 370987 500688 371153
rect 500568 370953 500611 370987
rect 500645 370953 500688 370987
rect 500568 370787 500688 370953
rect 500568 370753 500611 370787
rect 500645 370753 500688 370787
rect 500568 370587 500688 370753
rect 500568 370553 500611 370587
rect 500645 370553 500688 370587
rect 500568 370387 500688 370553
rect 500568 370353 500611 370387
rect 500645 370353 500688 370387
rect 500568 370187 500688 370353
rect 500568 370153 500611 370187
rect 500645 370153 500688 370187
rect 500568 369987 500688 370153
rect 500568 369953 500611 369987
rect 500645 369953 500688 369987
rect 500568 369787 500688 369953
rect 500568 369753 500611 369787
rect 500645 369753 500688 369787
rect 500568 369587 500688 369753
rect 500568 369553 500611 369587
rect 500645 369553 500688 369587
rect 500568 369387 500688 369553
rect 500568 369353 500611 369387
rect 500645 369353 500688 369387
rect 500568 369187 500688 369353
rect 500568 369153 500611 369187
rect 500645 369153 500688 369187
rect 500568 368987 500688 369153
rect 500568 368953 500611 368987
rect 500645 368953 500688 368987
rect 500568 368787 500688 368953
rect 500568 368753 500611 368787
rect 500645 368753 500688 368787
rect 500568 368587 500688 368753
rect 500568 368553 500611 368587
rect 500645 368553 500688 368587
rect 500568 368387 500688 368553
rect 500568 368353 500611 368387
rect 500645 368353 500688 368387
rect 500568 368187 500688 368353
rect 500568 368153 500611 368187
rect 500645 368153 500688 368187
rect 500568 367987 500688 368153
rect 500568 367953 500611 367987
rect 500645 367953 500688 367987
rect 500568 367787 500688 367953
rect 500568 367753 500611 367787
rect 500645 367753 500688 367787
rect 500568 367587 500688 367753
rect 500568 367553 500611 367587
rect 500645 367553 500688 367587
rect 500568 367387 500688 367553
rect 500568 367353 500611 367387
rect 500645 367353 500688 367387
rect 500568 367187 500688 367353
rect 500568 367153 500611 367187
rect 500645 367153 500688 367187
rect 500568 366987 500688 367153
rect 500568 366953 500611 366987
rect 500645 366953 500688 366987
rect 500568 366787 500688 366953
rect 500568 366753 500611 366787
rect 500645 366753 500688 366787
rect 500568 366587 500688 366753
rect 500568 366553 500611 366587
rect 500645 366553 500688 366587
rect 500568 366387 500688 366553
rect 500568 366353 500611 366387
rect 500645 366353 500688 366387
rect 500568 366187 500688 366353
rect 500568 366153 500611 366187
rect 500645 366153 500688 366187
rect 500568 365987 500688 366153
rect 500568 365953 500611 365987
rect 500645 365953 500688 365987
rect 500568 365787 500688 365953
rect 500568 365753 500611 365787
rect 500645 365753 500688 365787
rect 500568 365587 500688 365753
rect 500568 365553 500611 365587
rect 500645 365553 500688 365587
rect 500568 365387 500688 365553
rect 500568 365353 500611 365387
rect 500645 365353 500688 365387
rect 500568 365187 500688 365353
rect 500568 365153 500611 365187
rect 500645 365153 500688 365187
rect 500568 364987 500688 365153
rect 500568 364953 500611 364987
rect 500645 364953 500688 364987
rect 500568 364787 500688 364953
rect 500568 364753 500611 364787
rect 500645 364753 500688 364787
rect 500568 364587 500688 364753
rect 500568 364553 500611 364587
rect 500645 364553 500688 364587
rect 500568 364387 500688 364553
rect 500568 364353 500611 364387
rect 500645 364353 500688 364387
rect 500568 364187 500688 364353
rect 500568 364153 500611 364187
rect 500645 364153 500688 364187
rect 500568 363987 500688 364153
rect 500568 363953 500611 363987
rect 500645 363953 500688 363987
rect 500568 363787 500688 363953
rect 500568 363753 500611 363787
rect 500645 363753 500688 363787
rect 500568 363587 500688 363753
rect 500568 363553 500611 363587
rect 500645 363553 500688 363587
rect 500568 363387 500688 363553
rect 500568 363353 500611 363387
rect 500645 363353 500688 363387
rect 500568 363187 500688 363353
rect 500568 363153 500611 363187
rect 500645 363153 500688 363187
rect 500568 362987 500688 363153
rect 500568 362953 500611 362987
rect 500645 362953 500688 362987
rect 500568 362787 500688 362953
rect 500568 362753 500611 362787
rect 500645 362753 500688 362787
rect 500568 362587 500688 362753
rect 500568 362553 500611 362587
rect 500645 362553 500688 362587
rect 500568 361476 500688 362553
rect 500938 372910 500944 372924
rect 500978 372910 501008 372930
rect 500938 372854 501008 372910
rect 500938 372820 500944 372854
rect 500978 372820 501008 372854
rect 500938 372764 501008 372820
rect 500938 372730 500944 372764
rect 500978 372730 501008 372764
rect 500938 372674 501008 372730
rect 500938 372640 500944 372674
rect 500978 372640 501008 372674
rect 500938 372584 501008 372640
rect 500938 372550 500944 372584
rect 500978 372550 501008 372584
rect 500938 372494 501008 372550
rect 500938 372460 500944 372494
rect 500978 372460 501008 372494
rect 500938 372404 501008 372460
rect 500938 372370 500944 372404
rect 500978 372370 501008 372404
rect 500938 372314 501008 372370
rect 500938 372280 500944 372314
rect 500978 372280 501008 372314
rect 500938 372224 501008 372280
rect 500938 372190 500944 372224
rect 500978 372190 501008 372224
rect 500938 372134 501008 372190
rect 500938 372100 500944 372134
rect 500978 372100 501008 372134
rect 500938 372044 501008 372100
rect 500938 372010 500944 372044
rect 500978 372010 501008 372044
rect 500938 371954 501008 372010
rect 500938 371920 500944 371954
rect 500978 371920 501008 371954
rect 500938 371784 501008 371920
rect 500938 371750 500944 371784
rect 500978 371750 501008 371784
rect 500938 371694 501008 371750
rect 500938 371660 500944 371694
rect 500978 371660 501008 371694
rect 500938 371604 501008 371660
rect 500938 371570 500944 371604
rect 500978 371570 501008 371604
rect 500938 371514 501008 371570
rect 500938 371480 500944 371514
rect 500978 371480 501008 371514
rect 500938 371424 501008 371480
rect 500938 371390 500944 371424
rect 500978 371390 501008 371424
rect 500938 371334 501008 371390
rect 500938 371300 500944 371334
rect 500978 371300 501008 371334
rect 500938 371244 501008 371300
rect 500938 371210 500944 371244
rect 500978 371210 501008 371244
rect 500938 371154 501008 371210
rect 500938 371120 500944 371154
rect 500978 371120 501008 371154
rect 500938 371064 501008 371120
rect 500938 371030 500944 371064
rect 500978 371030 501008 371064
rect 500938 370974 501008 371030
rect 500938 370940 500944 370974
rect 500978 370940 501008 370974
rect 500938 370884 501008 370940
rect 500938 370850 500944 370884
rect 500978 370850 501008 370884
rect 500938 370794 501008 370850
rect 500938 370760 500944 370794
rect 500978 370760 501008 370794
rect 500938 370704 501008 370760
rect 500938 370670 500944 370704
rect 500978 370670 501008 370704
rect 500938 370614 501008 370670
rect 500938 370580 500944 370614
rect 500978 370580 501008 370614
rect 500938 370444 501008 370580
rect 500938 370410 500944 370444
rect 500978 370410 501008 370444
rect 500938 370354 501008 370410
rect 500938 370320 500944 370354
rect 500978 370320 501008 370354
rect 500938 370264 501008 370320
rect 500938 370230 500944 370264
rect 500978 370230 501008 370264
rect 500938 370174 501008 370230
rect 500938 370140 500944 370174
rect 500978 370140 501008 370174
rect 500938 370084 501008 370140
rect 500938 370050 500944 370084
rect 500978 370050 501008 370084
rect 500938 369994 501008 370050
rect 500938 369960 500944 369994
rect 500978 369960 501008 369994
rect 500938 369904 501008 369960
rect 500938 369870 500944 369904
rect 500978 369870 501008 369904
rect 500938 369814 501008 369870
rect 500938 369780 500944 369814
rect 500978 369780 501008 369814
rect 500938 369724 501008 369780
rect 500938 369690 500944 369724
rect 500978 369690 501008 369724
rect 500938 369634 501008 369690
rect 500938 369600 500944 369634
rect 500978 369600 501008 369634
rect 500938 369544 501008 369600
rect 500938 369510 500944 369544
rect 500978 369510 501008 369544
rect 500938 369454 501008 369510
rect 500938 369420 500944 369454
rect 500978 369420 501008 369454
rect 500938 369364 501008 369420
rect 500938 369330 500944 369364
rect 500978 369330 501008 369364
rect 500938 369274 501008 369330
rect 500938 369240 500944 369274
rect 500978 369240 501008 369274
rect 500938 369104 501008 369240
rect 500938 369070 500944 369104
rect 500978 369070 501008 369104
rect 500938 369014 501008 369070
rect 500938 368980 500944 369014
rect 500978 368980 501008 369014
rect 500938 368924 501008 368980
rect 500938 368890 500944 368924
rect 500978 368890 501008 368924
rect 500938 368834 501008 368890
rect 500938 368800 500944 368834
rect 500978 368800 501008 368834
rect 500938 368744 501008 368800
rect 500938 368710 500944 368744
rect 500978 368710 501008 368744
rect 500938 368654 501008 368710
rect 500938 368620 500944 368654
rect 500978 368620 501008 368654
rect 500938 368564 501008 368620
rect 500938 368530 500944 368564
rect 500978 368530 501008 368564
rect 500938 368474 501008 368530
rect 500938 368440 500944 368474
rect 500978 368440 501008 368474
rect 500938 368384 501008 368440
rect 500938 368350 500944 368384
rect 500978 368350 501008 368384
rect 500938 368294 501008 368350
rect 500938 368260 500944 368294
rect 500978 368260 501008 368294
rect 500938 368204 501008 368260
rect 500938 368170 500944 368204
rect 500978 368170 501008 368204
rect 500938 368114 501008 368170
rect 500938 368080 500944 368114
rect 500978 368080 501008 368114
rect 500938 368024 501008 368080
rect 500938 367990 500944 368024
rect 500978 367990 501008 368024
rect 500938 367934 501008 367990
rect 500938 367900 500944 367934
rect 500978 367900 501008 367934
rect 500938 367764 501008 367900
rect 500938 367730 500944 367764
rect 500978 367730 501008 367764
rect 500938 367674 501008 367730
rect 500938 367640 500944 367674
rect 500978 367640 501008 367674
rect 500938 367584 501008 367640
rect 500938 367550 500944 367584
rect 500978 367550 501008 367584
rect 500938 367494 501008 367550
rect 500938 367460 500944 367494
rect 500978 367460 501008 367494
rect 500938 367404 501008 367460
rect 500938 367370 500944 367404
rect 500978 367370 501008 367404
rect 500938 367314 501008 367370
rect 500938 367280 500944 367314
rect 500978 367280 501008 367314
rect 500938 367224 501008 367280
rect 500938 367190 500944 367224
rect 500978 367190 501008 367224
rect 500938 367134 501008 367190
rect 500938 367100 500944 367134
rect 500978 367100 501008 367134
rect 500938 367044 501008 367100
rect 500938 367010 500944 367044
rect 500978 367010 501008 367044
rect 500938 366954 501008 367010
rect 500938 366920 500944 366954
rect 500978 366920 501008 366954
rect 500938 366864 501008 366920
rect 500938 366830 500944 366864
rect 500978 366830 501008 366864
rect 500938 366774 501008 366830
rect 500938 366740 500944 366774
rect 500978 366740 501008 366774
rect 500938 366684 501008 366740
rect 500938 366650 500944 366684
rect 500978 366650 501008 366684
rect 500938 366594 501008 366650
rect 500938 366560 500944 366594
rect 500978 366560 501008 366594
rect 500938 366424 501008 366560
rect 500938 366390 500944 366424
rect 500978 366390 501008 366424
rect 500938 366334 501008 366390
rect 500938 366300 500944 366334
rect 500978 366300 501008 366334
rect 500938 366244 501008 366300
rect 500938 366210 500944 366244
rect 500978 366210 501008 366244
rect 500938 366154 501008 366210
rect 500938 366120 500944 366154
rect 500978 366120 501008 366154
rect 500938 366064 501008 366120
rect 500938 366030 500944 366064
rect 500978 366030 501008 366064
rect 500938 365974 501008 366030
rect 500938 365940 500944 365974
rect 500978 365940 501008 365974
rect 500938 365884 501008 365940
rect 500938 365850 500944 365884
rect 500978 365850 501008 365884
rect 500938 365794 501008 365850
rect 500938 365760 500944 365794
rect 500978 365760 501008 365794
rect 500938 365704 501008 365760
rect 500938 365670 500944 365704
rect 500978 365670 501008 365704
rect 500938 365614 501008 365670
rect 500938 365580 500944 365614
rect 500978 365580 501008 365614
rect 500938 365524 501008 365580
rect 500938 365490 500944 365524
rect 500978 365490 501008 365524
rect 500938 365434 501008 365490
rect 500938 365400 500944 365434
rect 500978 365400 501008 365434
rect 500938 365344 501008 365400
rect 500938 365310 500944 365344
rect 500978 365310 501008 365344
rect 500938 365254 501008 365310
rect 500938 365220 500944 365254
rect 500978 365220 501008 365254
rect 500938 365084 501008 365220
rect 500938 365050 500944 365084
rect 500978 365050 501008 365084
rect 500938 364994 501008 365050
rect 500938 364960 500944 364994
rect 500978 364960 501008 364994
rect 500938 364904 501008 364960
rect 500938 364870 500944 364904
rect 500978 364870 501008 364904
rect 500938 364814 501008 364870
rect 500938 364780 500944 364814
rect 500978 364780 501008 364814
rect 500938 364724 501008 364780
rect 500938 364690 500944 364724
rect 500978 364690 501008 364724
rect 500938 364634 501008 364690
rect 500938 364600 500944 364634
rect 500978 364600 501008 364634
rect 500938 364544 501008 364600
rect 500938 364510 500944 364544
rect 500978 364510 501008 364544
rect 500938 364454 501008 364510
rect 500938 364420 500944 364454
rect 500978 364420 501008 364454
rect 500938 364364 501008 364420
rect 500938 364330 500944 364364
rect 500978 364330 501008 364364
rect 500938 364274 501008 364330
rect 500938 364240 500944 364274
rect 500978 364240 501008 364274
rect 500938 364184 501008 364240
rect 500938 364150 500944 364184
rect 500978 364150 501008 364184
rect 500938 364094 501008 364150
rect 500938 364060 500944 364094
rect 500978 364060 501008 364094
rect 500938 364004 501008 364060
rect 500938 363970 500944 364004
rect 500978 363970 501008 364004
rect 500938 363914 501008 363970
rect 500938 363880 500944 363914
rect 500978 363880 501008 363914
rect 500938 363744 501008 363880
rect 500938 363710 500944 363744
rect 500978 363710 501008 363744
rect 500938 363654 501008 363710
rect 500938 363620 500944 363654
rect 500978 363620 501008 363654
rect 500938 363564 501008 363620
rect 500938 363530 500944 363564
rect 500978 363530 501008 363564
rect 500938 363474 501008 363530
rect 500938 363440 500944 363474
rect 500978 363440 501008 363474
rect 500938 363384 501008 363440
rect 500938 363350 500944 363384
rect 500978 363350 501008 363384
rect 500938 363294 501008 363350
rect 500938 363260 500944 363294
rect 500978 363260 501008 363294
rect 500938 363204 501008 363260
rect 500938 363170 500944 363204
rect 500978 363170 501008 363204
rect 500938 363114 501008 363170
rect 500938 363080 500944 363114
rect 500978 363080 501008 363114
rect 500938 363024 501008 363080
rect 500938 362990 500944 363024
rect 500978 362990 501008 363024
rect 500938 362934 501008 362990
rect 500938 362900 500944 362934
rect 500978 362900 501008 362934
rect 500938 362844 501008 362900
rect 500938 362810 500944 362844
rect 500978 362810 501008 362844
rect 500938 362754 501008 362810
rect 500938 362720 500944 362754
rect 500978 362720 501008 362754
rect 500938 362664 501008 362720
rect 500938 362630 500944 362664
rect 500978 362630 501008 362664
rect 501088 372960 501132 372980
rect 501088 372926 501104 372960
rect 501138 372926 501184 372930
rect 501088 372924 501184 372926
rect 501088 372870 501158 372924
rect 501088 372836 501104 372870
rect 501138 372836 501158 372870
rect 501088 372780 501158 372836
rect 501088 372746 501104 372780
rect 501138 372746 501158 372780
rect 501088 372690 501158 372746
rect 501088 372656 501104 372690
rect 501138 372656 501158 372690
rect 501088 372600 501158 372656
rect 501088 372566 501104 372600
rect 501138 372566 501158 372600
rect 501088 372510 501158 372566
rect 501088 372476 501104 372510
rect 501138 372476 501158 372510
rect 501088 372420 501158 372476
rect 501088 372386 501104 372420
rect 501138 372386 501158 372420
rect 501088 372330 501158 372386
rect 501088 372296 501104 372330
rect 501138 372296 501158 372330
rect 501088 372240 501158 372296
rect 501088 372206 501104 372240
rect 501138 372206 501158 372240
rect 501088 372150 501158 372206
rect 501088 372116 501104 372150
rect 501138 372116 501158 372150
rect 501088 372060 501158 372116
rect 501088 372026 501104 372060
rect 501138 372026 501158 372060
rect 501088 371620 501158 372026
rect 501088 371586 501104 371620
rect 501138 371586 501158 371620
rect 501088 371530 501158 371586
rect 501088 371496 501104 371530
rect 501138 371496 501158 371530
rect 501088 371440 501158 371496
rect 501088 371406 501104 371440
rect 501138 371406 501158 371440
rect 501088 371350 501158 371406
rect 501088 371316 501104 371350
rect 501138 371316 501158 371350
rect 501088 371260 501158 371316
rect 501088 371226 501104 371260
rect 501138 371226 501158 371260
rect 501088 371170 501158 371226
rect 501088 371136 501104 371170
rect 501138 371136 501158 371170
rect 501088 371080 501158 371136
rect 501088 371046 501104 371080
rect 501138 371046 501158 371080
rect 501088 370990 501158 371046
rect 501088 370956 501104 370990
rect 501138 370956 501158 370990
rect 501088 370900 501158 370956
rect 501088 370866 501104 370900
rect 501138 370866 501158 370900
rect 501088 370810 501158 370866
rect 501088 370776 501104 370810
rect 501138 370776 501158 370810
rect 501088 370720 501158 370776
rect 501088 370686 501104 370720
rect 501138 370686 501158 370720
rect 501088 370280 501158 370686
rect 501088 370246 501104 370280
rect 501138 370246 501158 370280
rect 501088 370190 501158 370246
rect 501088 370156 501104 370190
rect 501138 370156 501158 370190
rect 501088 370100 501158 370156
rect 501088 370066 501104 370100
rect 501138 370066 501158 370100
rect 501088 370010 501158 370066
rect 501088 369976 501104 370010
rect 501138 369976 501158 370010
rect 501088 369920 501158 369976
rect 501088 369886 501104 369920
rect 501138 369886 501158 369920
rect 501088 369830 501158 369886
rect 501088 369796 501104 369830
rect 501138 369796 501158 369830
rect 501088 369740 501158 369796
rect 501088 369706 501104 369740
rect 501138 369706 501158 369740
rect 501088 369650 501158 369706
rect 501088 369616 501104 369650
rect 501138 369616 501158 369650
rect 501088 369560 501158 369616
rect 501088 369526 501104 369560
rect 501138 369526 501158 369560
rect 501088 369470 501158 369526
rect 501088 369436 501104 369470
rect 501138 369436 501158 369470
rect 501088 369380 501158 369436
rect 501088 369346 501104 369380
rect 501138 369346 501158 369380
rect 501088 368940 501158 369346
rect 501088 368906 501104 368940
rect 501138 368906 501158 368940
rect 501088 368850 501158 368906
rect 501088 368816 501104 368850
rect 501138 368816 501158 368850
rect 501088 368760 501158 368816
rect 501088 368726 501104 368760
rect 501138 368726 501158 368760
rect 501088 368670 501158 368726
rect 501088 368636 501104 368670
rect 501138 368636 501158 368670
rect 501088 368580 501158 368636
rect 501088 368546 501104 368580
rect 501138 368546 501158 368580
rect 501088 368490 501158 368546
rect 501088 368456 501104 368490
rect 501138 368456 501158 368490
rect 501088 368400 501158 368456
rect 501088 368366 501104 368400
rect 501138 368366 501158 368400
rect 501088 368310 501158 368366
rect 501088 368276 501104 368310
rect 501138 368276 501158 368310
rect 501088 368220 501158 368276
rect 501088 368186 501104 368220
rect 501138 368186 501158 368220
rect 501088 368130 501158 368186
rect 501088 368096 501104 368130
rect 501138 368096 501158 368130
rect 501088 368040 501158 368096
rect 501088 368006 501104 368040
rect 501138 368006 501158 368040
rect 501088 367600 501158 368006
rect 501088 367566 501104 367600
rect 501138 367566 501158 367600
rect 501088 367510 501158 367566
rect 501088 367476 501104 367510
rect 501138 367476 501158 367510
rect 501088 367420 501158 367476
rect 501088 367386 501104 367420
rect 501138 367386 501158 367420
rect 501088 367330 501158 367386
rect 501088 367296 501104 367330
rect 501138 367296 501158 367330
rect 501088 367240 501158 367296
rect 501088 367206 501104 367240
rect 501138 367206 501158 367240
rect 501088 367150 501158 367206
rect 501088 367116 501104 367150
rect 501138 367116 501158 367150
rect 501088 367060 501158 367116
rect 501088 367026 501104 367060
rect 501138 367026 501158 367060
rect 501088 366970 501158 367026
rect 501088 366936 501104 366970
rect 501138 366936 501158 366970
rect 501088 366880 501158 366936
rect 501088 366846 501104 366880
rect 501138 366846 501158 366880
rect 501088 366790 501158 366846
rect 501088 366756 501104 366790
rect 501138 366756 501158 366790
rect 501088 366700 501158 366756
rect 501088 366666 501104 366700
rect 501138 366666 501158 366700
rect 501088 366260 501158 366666
rect 501088 366226 501104 366260
rect 501138 366226 501158 366260
rect 501088 366170 501158 366226
rect 501088 366136 501104 366170
rect 501138 366136 501158 366170
rect 501088 366080 501158 366136
rect 501088 366046 501104 366080
rect 501138 366046 501158 366080
rect 501088 365990 501158 366046
rect 501088 365956 501104 365990
rect 501138 365956 501158 365990
rect 501088 365900 501158 365956
rect 501088 365866 501104 365900
rect 501138 365866 501158 365900
rect 501088 365810 501158 365866
rect 501088 365776 501104 365810
rect 501138 365776 501158 365810
rect 501088 365720 501158 365776
rect 501088 365686 501104 365720
rect 501138 365686 501158 365720
rect 501088 365630 501158 365686
rect 501088 365596 501104 365630
rect 501138 365596 501158 365630
rect 501088 365540 501158 365596
rect 501088 365506 501104 365540
rect 501138 365506 501158 365540
rect 501088 365450 501158 365506
rect 501088 365416 501104 365450
rect 501138 365416 501158 365450
rect 501088 365360 501158 365416
rect 501088 365326 501104 365360
rect 501138 365326 501158 365360
rect 501088 364920 501158 365326
rect 501088 364886 501104 364920
rect 501138 364886 501158 364920
rect 501088 364830 501158 364886
rect 501088 364796 501104 364830
rect 501138 364796 501158 364830
rect 501088 364740 501158 364796
rect 501088 364706 501104 364740
rect 501138 364706 501158 364740
rect 501088 364650 501158 364706
rect 501088 364616 501104 364650
rect 501138 364616 501158 364650
rect 501088 364560 501158 364616
rect 501088 364526 501104 364560
rect 501138 364526 501158 364560
rect 501088 364470 501158 364526
rect 501088 364436 501104 364470
rect 501138 364436 501158 364470
rect 501088 364380 501158 364436
rect 501088 364346 501104 364380
rect 501138 364346 501158 364380
rect 501088 364290 501158 364346
rect 501088 364256 501104 364290
rect 501138 364256 501158 364290
rect 501088 364200 501158 364256
rect 501088 364166 501104 364200
rect 501138 364166 501158 364200
rect 501088 364110 501158 364166
rect 501088 364076 501104 364110
rect 501138 364076 501158 364110
rect 501088 364020 501158 364076
rect 501088 363986 501104 364020
rect 501138 363986 501158 364020
rect 501088 363580 501158 363986
rect 501088 363546 501104 363580
rect 501138 363546 501158 363580
rect 501088 363490 501158 363546
rect 501088 363456 501104 363490
rect 501138 363456 501158 363490
rect 501088 363400 501158 363456
rect 501088 363366 501104 363400
rect 501138 363366 501158 363400
rect 501088 363310 501158 363366
rect 501088 363276 501104 363310
rect 501138 363276 501158 363310
rect 501088 363220 501158 363276
rect 501088 363186 501104 363220
rect 501138 363186 501158 363220
rect 501088 363130 501158 363186
rect 501088 363096 501104 363130
rect 501138 363096 501158 363130
rect 501088 363040 501158 363096
rect 501088 363006 501104 363040
rect 501138 363006 501158 363040
rect 501088 362950 501158 363006
rect 501088 362916 501104 362950
rect 501138 362916 501158 362950
rect 501088 362860 501158 362916
rect 501088 362826 501104 362860
rect 501138 362826 501158 362860
rect 501088 362770 501158 362826
rect 501262 372798 501874 372806
rect 501262 372774 501812 372798
rect 501262 372740 501308 372774
rect 501342 372740 501408 372774
rect 501442 372740 501508 372774
rect 501542 372740 501608 372774
rect 501642 372740 501708 372774
rect 501742 372740 501808 372774
rect 501864 372746 501874 372798
rect 501842 372740 501874 372746
rect 501262 372674 501874 372740
rect 501262 372640 501308 372674
rect 501342 372640 501408 372674
rect 501442 372640 501508 372674
rect 501542 372640 501608 372674
rect 501642 372640 501708 372674
rect 501742 372640 501808 372674
rect 501842 372640 501874 372674
rect 501262 372574 501874 372640
rect 501262 372540 501308 372574
rect 501342 372540 501408 372574
rect 501442 372540 501508 372574
rect 501542 372540 501608 372574
rect 501642 372540 501708 372574
rect 501742 372540 501808 372574
rect 501842 372540 501874 372574
rect 501262 372474 501874 372540
rect 501262 372440 501308 372474
rect 501342 372440 501408 372474
rect 501442 372440 501508 372474
rect 501542 372440 501608 372474
rect 501642 372440 501708 372474
rect 501742 372440 501808 372474
rect 501842 372440 501874 372474
rect 501262 372374 501874 372440
rect 501262 372340 501308 372374
rect 501342 372340 501408 372374
rect 501442 372340 501508 372374
rect 501542 372340 501608 372374
rect 501642 372340 501708 372374
rect 501742 372340 501808 372374
rect 501842 372340 501874 372374
rect 501262 372274 501874 372340
rect 501262 372240 501308 372274
rect 501342 372240 501408 372274
rect 501442 372240 501508 372274
rect 501542 372240 501608 372274
rect 501642 372240 501708 372274
rect 501742 372240 501808 372274
rect 501842 372240 501874 372274
rect 501262 371434 501874 372240
rect 501262 371400 501308 371434
rect 501342 371400 501408 371434
rect 501442 371400 501508 371434
rect 501542 371400 501608 371434
rect 501642 371400 501708 371434
rect 501742 371400 501808 371434
rect 501842 371400 501874 371434
rect 501262 371334 501874 371400
rect 501262 371300 501308 371334
rect 501342 371300 501408 371334
rect 501442 371300 501508 371334
rect 501542 371300 501608 371334
rect 501642 371300 501708 371334
rect 501742 371300 501808 371334
rect 501842 371300 501874 371334
rect 501262 371234 501874 371300
rect 501262 371200 501308 371234
rect 501342 371200 501408 371234
rect 501442 371200 501508 371234
rect 501542 371200 501608 371234
rect 501642 371200 501708 371234
rect 501742 371200 501808 371234
rect 501842 371200 501874 371234
rect 501262 371134 501874 371200
rect 501262 371100 501308 371134
rect 501342 371100 501408 371134
rect 501442 371100 501508 371134
rect 501542 371100 501608 371134
rect 501642 371100 501708 371134
rect 501742 371100 501808 371134
rect 501842 371100 501874 371134
rect 501262 371034 501874 371100
rect 501262 371000 501308 371034
rect 501342 371000 501408 371034
rect 501442 371000 501508 371034
rect 501542 371000 501608 371034
rect 501642 371000 501708 371034
rect 501742 371000 501808 371034
rect 501842 371000 501874 371034
rect 501262 370934 501874 371000
rect 501262 370900 501308 370934
rect 501342 370900 501408 370934
rect 501442 370900 501508 370934
rect 501542 370900 501608 370934
rect 501642 370900 501708 370934
rect 501742 370900 501808 370934
rect 501842 370900 501874 370934
rect 501262 370866 501874 370900
rect 501262 370814 501268 370866
rect 501320 370814 501874 370866
rect 501262 370094 501874 370814
rect 501262 370060 501308 370094
rect 501342 370060 501408 370094
rect 501442 370060 501508 370094
rect 501542 370060 501608 370094
rect 501642 370060 501708 370094
rect 501742 370060 501808 370094
rect 501842 370060 501874 370094
rect 501262 369994 501874 370060
rect 501262 369960 501308 369994
rect 501342 369960 501408 369994
rect 501442 369960 501508 369994
rect 501542 369960 501608 369994
rect 501642 369960 501708 369994
rect 501742 369960 501808 369994
rect 501842 369960 501874 369994
rect 501262 369894 501874 369960
rect 501262 369860 501308 369894
rect 501342 369860 501408 369894
rect 501442 369860 501508 369894
rect 501542 369860 501608 369894
rect 501642 369860 501708 369894
rect 501742 369860 501808 369894
rect 501842 369860 501874 369894
rect 501262 369794 501874 369860
rect 501262 369760 501308 369794
rect 501342 369760 501408 369794
rect 501442 369760 501508 369794
rect 501542 369760 501608 369794
rect 501642 369760 501708 369794
rect 501742 369760 501808 369794
rect 501842 369760 501874 369794
rect 501262 369694 501874 369760
rect 501262 369660 501308 369694
rect 501342 369660 501408 369694
rect 501442 369660 501508 369694
rect 501542 369660 501608 369694
rect 501642 369660 501708 369694
rect 501742 369660 501808 369694
rect 501842 369660 501874 369694
rect 501262 369594 501874 369660
rect 501262 369560 501308 369594
rect 501342 369560 501408 369594
rect 501442 369560 501508 369594
rect 501542 369560 501608 369594
rect 501642 369560 501708 369594
rect 501742 369560 501808 369594
rect 501842 369560 501874 369594
rect 501262 368754 501874 369560
rect 501262 368720 501308 368754
rect 501342 368720 501408 368754
rect 501442 368720 501508 368754
rect 501542 368720 501608 368754
rect 501642 368720 501708 368754
rect 501742 368720 501808 368754
rect 501842 368720 501874 368754
rect 501262 368654 501874 368720
rect 501262 368620 501308 368654
rect 501342 368620 501408 368654
rect 501442 368620 501508 368654
rect 501542 368620 501608 368654
rect 501642 368620 501708 368654
rect 501742 368620 501808 368654
rect 501842 368620 501874 368654
rect 501262 368554 501874 368620
rect 501262 368520 501308 368554
rect 501342 368520 501408 368554
rect 501442 368520 501508 368554
rect 501542 368520 501608 368554
rect 501642 368520 501708 368554
rect 501742 368520 501808 368554
rect 501842 368520 501874 368554
rect 501262 368454 501874 368520
rect 501262 368420 501308 368454
rect 501342 368420 501408 368454
rect 501442 368420 501508 368454
rect 501542 368420 501608 368454
rect 501642 368420 501708 368454
rect 501742 368420 501808 368454
rect 501842 368420 501874 368454
rect 501262 368354 501874 368420
rect 501262 368320 501308 368354
rect 501342 368320 501408 368354
rect 501442 368320 501508 368354
rect 501542 368320 501608 368354
rect 501642 368320 501708 368354
rect 501742 368320 501808 368354
rect 501842 368320 501874 368354
rect 501262 368254 501874 368320
rect 501262 368220 501308 368254
rect 501342 368220 501408 368254
rect 501442 368220 501508 368254
rect 501542 368220 501608 368254
rect 501642 368220 501708 368254
rect 501742 368220 501808 368254
rect 501842 368220 501874 368254
rect 501262 367414 501874 368220
rect 501262 367380 501308 367414
rect 501342 367380 501408 367414
rect 501442 367380 501508 367414
rect 501542 367380 501608 367414
rect 501642 367380 501708 367414
rect 501742 367380 501808 367414
rect 501842 367380 501874 367414
rect 501262 367314 501874 367380
rect 501262 367280 501308 367314
rect 501342 367280 501408 367314
rect 501442 367280 501508 367314
rect 501542 367280 501608 367314
rect 501642 367280 501708 367314
rect 501742 367280 501808 367314
rect 501842 367280 501874 367314
rect 501262 367214 501874 367280
rect 501262 367180 501308 367214
rect 501342 367180 501408 367214
rect 501442 367180 501508 367214
rect 501542 367180 501608 367214
rect 501642 367180 501708 367214
rect 501742 367180 501808 367214
rect 501842 367180 501874 367214
rect 501262 367114 501874 367180
rect 501262 367080 501308 367114
rect 501342 367080 501408 367114
rect 501442 367080 501508 367114
rect 501542 367080 501608 367114
rect 501642 367080 501708 367114
rect 501742 367080 501808 367114
rect 501842 367080 501874 367114
rect 501262 367014 501874 367080
rect 501262 366980 501308 367014
rect 501342 366980 501408 367014
rect 501442 366980 501508 367014
rect 501542 366980 501608 367014
rect 501642 366980 501708 367014
rect 501742 366980 501808 367014
rect 501842 366980 501874 367014
rect 501262 366914 501874 366980
rect 501262 366880 501308 366914
rect 501342 366880 501408 366914
rect 501442 366880 501508 366914
rect 501542 366880 501608 366914
rect 501642 366880 501708 366914
rect 501742 366880 501808 366914
rect 501842 366880 501874 366914
rect 501262 366074 501874 366880
rect 502164 366640 502192 373479
rect 502448 372987 502568 373861
rect 502448 372953 502491 372987
rect 502525 372982 502568 372987
rect 502448 372930 502492 372953
rect 502544 372930 502568 372982
rect 502448 372787 502568 372930
rect 502448 372753 502491 372787
rect 502525 372753 502568 372787
rect 502448 372587 502568 372753
rect 502448 372553 502491 372587
rect 502525 372553 502568 372587
rect 502448 372387 502568 372553
rect 502448 372353 502491 372387
rect 502525 372353 502568 372387
rect 502448 372187 502568 372353
rect 502448 372153 502491 372187
rect 502525 372153 502568 372187
rect 502448 371987 502568 372153
rect 502448 371953 502491 371987
rect 502525 371953 502568 371987
rect 502448 371787 502568 371953
rect 502448 371753 502491 371787
rect 502525 371753 502568 371787
rect 502448 371587 502568 371753
rect 502448 371553 502491 371587
rect 502525 371553 502568 371587
rect 502448 371387 502568 371553
rect 502448 371353 502491 371387
rect 502525 371353 502568 371387
rect 502448 371187 502568 371353
rect 502448 371153 502491 371187
rect 502525 371153 502568 371187
rect 502448 370987 502568 371153
rect 502448 370953 502491 370987
rect 502525 370953 502568 370987
rect 502448 370787 502568 370953
rect 502448 370753 502491 370787
rect 502525 370753 502568 370787
rect 502448 370587 502568 370753
rect 502448 370553 502491 370587
rect 502525 370553 502568 370587
rect 502448 370387 502568 370553
rect 502448 370353 502491 370387
rect 502525 370353 502568 370387
rect 502448 370187 502568 370353
rect 502448 370153 502491 370187
rect 502525 370153 502568 370187
rect 502448 369987 502568 370153
rect 502448 369953 502491 369987
rect 502525 369953 502568 369987
rect 502448 369787 502568 369953
rect 502448 369753 502491 369787
rect 502525 369753 502568 369787
rect 502448 369587 502568 369753
rect 502448 369553 502491 369587
rect 502525 369553 502568 369587
rect 502448 369387 502568 369553
rect 502448 369353 502491 369387
rect 502525 369353 502568 369387
rect 502448 369187 502568 369353
rect 502448 369153 502491 369187
rect 502525 369153 502568 369187
rect 502448 368987 502568 369153
rect 502448 368953 502491 368987
rect 502525 368953 502568 368987
rect 502448 368787 502568 368953
rect 502448 368753 502491 368787
rect 502525 368753 502568 368787
rect 502448 368587 502568 368753
rect 502448 368553 502491 368587
rect 502525 368553 502568 368587
rect 502448 368387 502568 368553
rect 502448 368353 502491 368387
rect 502525 368353 502568 368387
rect 502448 368187 502568 368353
rect 502448 368153 502491 368187
rect 502525 368153 502568 368187
rect 502448 367987 502568 368153
rect 502448 367953 502491 367987
rect 502525 367953 502568 367987
rect 502448 367787 502568 367953
rect 502448 367753 502491 367787
rect 502525 367753 502568 367787
rect 502448 367587 502568 367753
rect 502448 367553 502491 367587
rect 502525 367553 502568 367587
rect 502448 367387 502568 367553
rect 502448 367353 502491 367387
rect 502525 367353 502568 367387
rect 502448 367187 502568 367353
rect 502448 367153 502491 367187
rect 502525 367153 502568 367187
rect 502448 366987 502568 367153
rect 502448 366953 502491 366987
rect 502525 366953 502568 366987
rect 502448 366787 502568 366953
rect 502448 366753 502491 366787
rect 502525 366753 502568 366787
rect 502152 366634 502204 366640
rect 502152 366576 502204 366582
rect 502448 366587 502568 366753
rect 501262 366040 501308 366074
rect 501342 366040 501408 366074
rect 501442 366040 501508 366074
rect 501542 366040 501608 366074
rect 501642 366040 501708 366074
rect 501742 366040 501808 366074
rect 501842 366040 501874 366074
rect 501262 365974 501874 366040
rect 501262 365940 501308 365974
rect 501342 365940 501408 365974
rect 501442 365940 501508 365974
rect 501542 365940 501608 365974
rect 501642 365940 501708 365974
rect 501742 365940 501808 365974
rect 501842 365940 501874 365974
rect 501262 365874 501874 365940
rect 501262 365840 501308 365874
rect 501342 365840 501408 365874
rect 501442 365840 501508 365874
rect 501542 365840 501608 365874
rect 501642 365840 501708 365874
rect 501742 365840 501808 365874
rect 501842 365840 501874 365874
rect 501262 365774 501874 365840
rect 501262 365740 501308 365774
rect 501342 365740 501408 365774
rect 501442 365740 501508 365774
rect 501542 365740 501608 365774
rect 501642 365740 501708 365774
rect 501742 365740 501808 365774
rect 501842 365740 501874 365774
rect 501262 365674 501874 365740
rect 501262 365640 501308 365674
rect 501342 365640 501408 365674
rect 501442 365640 501508 365674
rect 501542 365640 501608 365674
rect 501642 365640 501708 365674
rect 501742 365640 501808 365674
rect 501842 365640 501874 365674
rect 501262 365574 501874 365640
rect 501262 365540 501308 365574
rect 501342 365540 501408 365574
rect 501442 365540 501508 365574
rect 501542 365540 501608 365574
rect 501642 365540 501708 365574
rect 501742 365540 501808 365574
rect 501842 365540 501874 365574
rect 501262 364734 501874 365540
rect 501262 364700 501308 364734
rect 501342 364700 501408 364734
rect 501442 364700 501508 364734
rect 501542 364700 501608 364734
rect 501642 364700 501708 364734
rect 501742 364700 501808 364734
rect 501842 364700 501874 364734
rect 501262 364634 501874 364700
rect 501262 364600 501308 364634
rect 501342 364600 501408 364634
rect 501442 364600 501508 364634
rect 501542 364600 501608 364634
rect 501642 364600 501708 364634
rect 501742 364600 501808 364634
rect 501842 364600 501874 364634
rect 501262 364534 501874 364600
rect 501262 364500 501308 364534
rect 501342 364500 501408 364534
rect 501442 364500 501508 364534
rect 501542 364500 501608 364534
rect 501642 364500 501708 364534
rect 501742 364500 501808 364534
rect 501842 364500 501874 364534
rect 501262 364434 501874 364500
rect 501262 364400 501308 364434
rect 501342 364400 501408 364434
rect 501442 364400 501508 364434
rect 501542 364400 501608 364434
rect 501642 364400 501708 364434
rect 501742 364400 501808 364434
rect 501842 364400 501874 364434
rect 501262 364334 501874 364400
rect 501262 364300 501308 364334
rect 501342 364300 501408 364334
rect 501442 364300 501508 364334
rect 501542 364300 501608 364334
rect 501642 364300 501708 364334
rect 501742 364300 501808 364334
rect 501842 364300 501874 364334
rect 501262 364234 501874 364300
rect 501262 364200 501308 364234
rect 501342 364200 501408 364234
rect 501442 364200 501508 364234
rect 501542 364200 501608 364234
rect 501642 364200 501708 364234
rect 501742 364200 501808 364234
rect 501842 364200 501874 364234
rect 501262 363394 501874 364200
rect 501262 363360 501308 363394
rect 501342 363360 501408 363394
rect 501442 363360 501508 363394
rect 501542 363360 501608 363394
rect 501642 363360 501708 363394
rect 501742 363360 501808 363394
rect 501842 363360 501874 363394
rect 501262 363294 501874 363360
rect 501262 363260 501308 363294
rect 501342 363260 501408 363294
rect 501442 363260 501508 363294
rect 501542 363260 501608 363294
rect 501642 363260 501708 363294
rect 501742 363260 501808 363294
rect 501842 363260 501874 363294
rect 501262 363194 501874 363260
rect 501262 363160 501308 363194
rect 501342 363160 501408 363194
rect 501442 363160 501508 363194
rect 501542 363160 501608 363194
rect 501642 363160 501708 363194
rect 501742 363160 501808 363194
rect 501842 363160 501874 363194
rect 501262 363094 501874 363160
rect 501262 363060 501308 363094
rect 501342 363060 501408 363094
rect 501442 363060 501508 363094
rect 501542 363060 501608 363094
rect 501642 363060 501708 363094
rect 501742 363060 501808 363094
rect 501842 363060 501874 363094
rect 501262 362994 501874 363060
rect 501262 362960 501308 362994
rect 501342 362960 501408 362994
rect 501442 362960 501508 362994
rect 501542 362960 501608 362994
rect 501642 362960 501708 362994
rect 501742 362960 501808 362994
rect 501842 362960 501874 362994
rect 501262 362894 501874 362960
rect 501262 362860 501308 362894
rect 501342 362860 501408 362894
rect 501442 362860 501508 362894
rect 501542 362860 501608 362894
rect 501642 362860 501708 362894
rect 501742 362860 501808 362894
rect 501842 362860 501874 362894
rect 501262 362814 501874 362860
rect 502448 366553 502491 366587
rect 502525 366553 502568 366587
rect 502448 366387 502568 366553
rect 502448 366353 502491 366387
rect 502525 366353 502568 366387
rect 502448 366187 502568 366353
rect 502448 366153 502491 366187
rect 502525 366153 502568 366187
rect 502448 365987 502568 366153
rect 502448 365953 502491 365987
rect 502525 365953 502568 365987
rect 502448 365787 502568 365953
rect 502448 365753 502491 365787
rect 502525 365753 502568 365787
rect 502448 365587 502568 365753
rect 502448 365553 502491 365587
rect 502525 365553 502568 365587
rect 502448 365387 502568 365553
rect 502448 365353 502491 365387
rect 502525 365353 502568 365387
rect 502448 365187 502568 365353
rect 502448 365153 502491 365187
rect 502525 365153 502568 365187
rect 502448 364987 502568 365153
rect 502448 364953 502491 364987
rect 502525 364953 502568 364987
rect 502448 364787 502568 364953
rect 502448 364753 502491 364787
rect 502525 364753 502568 364787
rect 502448 364587 502568 364753
rect 502448 364553 502491 364587
rect 502525 364553 502568 364587
rect 502448 364387 502568 364553
rect 502448 364353 502491 364387
rect 502525 364353 502568 364387
rect 502448 364187 502568 364353
rect 502448 364153 502491 364187
rect 502525 364153 502568 364187
rect 502448 363987 502568 364153
rect 502448 363953 502491 363987
rect 502525 363953 502568 363987
rect 502448 363787 502568 363953
rect 502448 363753 502491 363787
rect 502525 363753 502568 363787
rect 502448 363587 502568 363753
rect 502448 363553 502491 363587
rect 502525 363553 502568 363587
rect 502448 363387 502568 363553
rect 502448 363353 502491 363387
rect 502525 363353 502568 363387
rect 502448 363187 502568 363353
rect 502448 363153 502491 363187
rect 502525 363153 502568 363187
rect 502448 362987 502568 363153
rect 502448 362953 502491 362987
rect 502525 362953 502568 362987
rect 501088 362736 501104 362770
rect 501138 362736 501158 362770
rect 501088 362680 501158 362736
rect 501088 362646 501104 362680
rect 501138 362646 501158 362680
rect 501088 362640 501158 362646
rect 502448 362787 502568 362953
rect 502448 362753 502491 362787
rect 502525 362753 502568 362787
rect 500938 362574 501008 362630
rect 500938 362540 500944 362574
rect 500978 362540 501008 362574
rect 500938 362476 501008 362540
rect 502448 362587 502568 362753
rect 502448 362553 502491 362587
rect 502525 362553 502568 362587
rect 500568 359888 500570 361476
rect 500686 359888 500688 361476
rect 500568 359866 500688 359888
rect 498688 357440 498690 359028
rect 498806 357440 498808 359028
rect 498688 357418 498808 357440
rect 502448 359028 502568 362553
rect 504328 378843 504448 379209
rect 504328 378809 504371 378843
rect 504405 378809 504448 378843
rect 504328 378443 504448 378809
rect 504328 378409 504371 378443
rect 504405 378409 504448 378443
rect 504328 378043 504448 378409
rect 504328 378009 504371 378043
rect 504405 378009 504448 378043
rect 504328 377386 504448 378009
rect 506208 380443 506328 380809
rect 506208 380409 506251 380443
rect 506285 380409 506328 380443
rect 506208 380043 506328 380409
rect 506208 380009 506251 380043
rect 506285 380009 506328 380043
rect 506208 379643 506328 380009
rect 506208 379609 506251 379643
rect 506285 379609 506328 379643
rect 506208 379243 506328 379609
rect 506208 379209 506251 379243
rect 506285 379209 506328 379243
rect 506208 378843 506328 379209
rect 506208 378809 506251 378843
rect 506285 378809 506328 378843
rect 506208 378443 506328 378809
rect 506208 378409 506251 378443
rect 506285 378409 506328 378443
rect 506208 378043 506328 378409
rect 506208 378009 506251 378043
rect 506285 378009 506328 378043
rect 504623 377435 505913 377441
rect 504623 377401 504639 377435
rect 504673 377401 504711 377435
rect 504745 377401 504783 377435
rect 504817 377401 504855 377435
rect 504889 377401 504927 377435
rect 504961 377401 504999 377435
rect 505033 377401 505071 377435
rect 505105 377401 505143 377435
rect 505177 377401 505215 377435
rect 505249 377401 505287 377435
rect 505321 377401 505359 377435
rect 505393 377401 505431 377435
rect 505465 377401 505503 377435
rect 505537 377401 505575 377435
rect 505609 377401 505647 377435
rect 505681 377401 505719 377435
rect 505753 377401 505791 377435
rect 505825 377401 505863 377435
rect 505897 377401 505913 377435
rect 506028 377401 506080 377404
rect 504535 377389 504581 377401
rect 504623 377395 505913 377401
rect 505997 377398 506080 377401
rect 504535 377386 504541 377389
rect 504328 377358 504541 377386
rect 504328 377299 504448 377358
rect 504535 377355 504541 377358
rect 504575 377355 504581 377389
rect 504535 377343 504581 377355
rect 505997 377389 506028 377398
rect 505997 377355 506003 377389
rect 505997 377346 506028 377355
rect 505997 377343 506080 377346
rect 506028 377340 506080 377343
rect 504328 377265 504371 377299
rect 504405 377265 504448 377299
rect 504328 376899 504448 377265
rect 506208 377299 506328 378009
rect 506208 377265 506251 377299
rect 506285 377265 506328 377299
rect 504623 376977 505913 376983
rect 504623 376943 504639 376977
rect 504673 376943 504711 376977
rect 504745 376943 504783 376977
rect 504817 376943 504855 376977
rect 504889 376943 504927 376977
rect 504961 376943 504999 376977
rect 505033 376943 505071 376977
rect 505105 376943 505143 376977
rect 505177 376943 505215 376977
rect 505249 376943 505287 376977
rect 505321 376943 505359 376977
rect 505393 376943 505431 376977
rect 505465 376943 505503 376977
rect 505537 376943 505575 376977
rect 505609 376943 505647 376977
rect 505681 376943 505719 376977
rect 505753 376943 505791 376977
rect 505825 376943 505863 376977
rect 505897 376943 505913 376977
rect 504623 376937 505913 376943
rect 504328 376865 504371 376899
rect 504405 376865 504448 376899
rect 504328 376499 504448 376865
rect 506208 376899 506328 377265
rect 506208 376865 506251 376899
rect 506285 376865 506328 376899
rect 504328 376465 504371 376499
rect 504405 376465 504448 376499
rect 504623 376519 505913 376525
rect 504623 376485 504639 376519
rect 504673 376485 504711 376519
rect 504745 376485 504783 376519
rect 504817 376485 504855 376519
rect 504889 376485 504927 376519
rect 504961 376485 504999 376519
rect 505033 376485 505071 376519
rect 505105 376485 505143 376519
rect 505177 376485 505215 376519
rect 505249 376485 505287 376519
rect 505321 376485 505359 376519
rect 505393 376485 505431 376519
rect 505465 376485 505503 376519
rect 505537 376485 505575 376519
rect 505609 376485 505647 376519
rect 505681 376485 505719 376519
rect 505753 376485 505791 376519
rect 505825 376485 505863 376519
rect 505897 376485 505913 376519
rect 504623 376479 505913 376485
rect 506208 376499 506328 376865
rect 504328 376099 504448 376465
rect 506208 376465 506251 376499
rect 506285 376465 506328 376499
rect 506108 376392 506136 376447
rect 506096 376386 506148 376392
rect 506096 376328 506148 376334
rect 504328 376065 504371 376099
rect 504405 376065 504448 376099
rect 506208 376099 506328 376465
rect 504328 375699 504448 376065
rect 504623 376061 505913 376067
rect 504623 376027 504639 376061
rect 504673 376027 504711 376061
rect 504745 376027 504783 376061
rect 504817 376027 504855 376061
rect 504889 376027 504927 376061
rect 504961 376027 504999 376061
rect 505033 376027 505071 376061
rect 505105 376027 505143 376061
rect 505177 376027 505215 376061
rect 505249 376027 505287 376061
rect 505321 376027 505359 376061
rect 505393 376027 505431 376061
rect 505465 376027 505503 376061
rect 505537 376027 505575 376061
rect 505609 376027 505647 376061
rect 505681 376027 505719 376061
rect 505753 376027 505791 376061
rect 505825 376027 505863 376061
rect 505897 376027 505913 376061
rect 504623 376021 505913 376027
rect 506208 376065 506251 376099
rect 506285 376065 506328 376099
rect 504328 375665 504371 375699
rect 504405 375665 504448 375699
rect 504328 375299 504448 375665
rect 506208 375699 506328 376065
rect 506208 375665 506251 375699
rect 506285 375665 506328 375699
rect 504623 375603 505913 375609
rect 504623 375569 504639 375603
rect 504673 375569 504711 375603
rect 504745 375569 504783 375603
rect 504817 375569 504855 375603
rect 504889 375569 504927 375603
rect 504961 375569 504999 375603
rect 505033 375569 505071 375603
rect 505105 375569 505143 375603
rect 505177 375569 505215 375603
rect 505249 375569 505287 375603
rect 505321 375569 505359 375603
rect 505393 375569 505431 375603
rect 505465 375569 505503 375603
rect 505537 375569 505575 375603
rect 505609 375569 505647 375603
rect 505681 375569 505719 375603
rect 505753 375569 505791 375603
rect 505825 375569 505863 375603
rect 505897 375569 505913 375603
rect 504623 375563 505913 375569
rect 504328 375265 504371 375299
rect 504405 375265 504448 375299
rect 504328 374899 504448 375265
rect 506208 375299 506328 375665
rect 506208 375265 506251 375299
rect 506285 375265 506328 375299
rect 504623 375145 505913 375151
rect 504623 375111 504639 375145
rect 504673 375111 504711 375145
rect 504745 375111 504783 375145
rect 504817 375111 504855 375145
rect 504889 375111 504927 375145
rect 504961 375111 504999 375145
rect 505033 375111 505071 375145
rect 505105 375111 505143 375145
rect 505177 375111 505215 375145
rect 505249 375111 505287 375145
rect 505321 375111 505359 375145
rect 505393 375111 505431 375145
rect 505465 375111 505503 375145
rect 505537 375111 505575 375145
rect 505609 375111 505647 375145
rect 505681 375111 505719 375145
rect 505753 375111 505791 375145
rect 505825 375111 505863 375145
rect 505897 375111 505913 375145
rect 504623 375105 505913 375111
rect 504328 374865 504371 374899
rect 504405 374865 504448 374899
rect 504328 372987 504448 374865
rect 506208 374899 506328 375265
rect 506208 374865 506251 374899
rect 506285 374865 506328 374899
rect 504623 374687 505913 374693
rect 504623 374653 504639 374687
rect 504673 374653 504711 374687
rect 504745 374653 504783 374687
rect 504817 374653 504855 374687
rect 504889 374653 504927 374687
rect 504961 374653 504999 374687
rect 505033 374653 505071 374687
rect 505105 374653 505143 374687
rect 505177 374653 505215 374687
rect 505249 374653 505287 374687
rect 505321 374653 505359 374687
rect 505393 374653 505431 374687
rect 505465 374653 505503 374687
rect 505537 374653 505575 374687
rect 505609 374653 505647 374687
rect 505681 374653 505719 374687
rect 505753 374653 505791 374687
rect 505825 374653 505863 374687
rect 505897 374653 505913 374687
rect 504623 374647 505913 374653
rect 504328 372953 504371 372987
rect 504405 372953 504448 372987
rect 504328 372787 504448 372953
rect 504328 372753 504371 372787
rect 504405 372753 504448 372787
rect 504328 372587 504448 372753
rect 504328 372553 504371 372587
rect 504405 372553 504448 372587
rect 504328 372387 504448 372553
rect 504328 372353 504371 372387
rect 504405 372353 504448 372387
rect 504328 372187 504448 372353
rect 504328 372153 504371 372187
rect 504405 372153 504448 372187
rect 504328 371987 504448 372153
rect 504328 371953 504371 371987
rect 504405 371953 504448 371987
rect 504328 371787 504448 371953
rect 504328 371753 504371 371787
rect 504405 371753 504448 371787
rect 504328 371587 504448 371753
rect 504328 371553 504371 371587
rect 504405 371553 504448 371587
rect 504328 371387 504448 371553
rect 504328 371353 504371 371387
rect 504405 371353 504448 371387
rect 504328 371187 504448 371353
rect 504328 371153 504371 371187
rect 504405 371153 504448 371187
rect 504328 370987 504448 371153
rect 504328 370953 504371 370987
rect 504405 370953 504448 370987
rect 504328 370787 504448 370953
rect 504328 370753 504371 370787
rect 504405 370753 504448 370787
rect 504328 370587 504448 370753
rect 504328 370553 504371 370587
rect 504405 370553 504448 370587
rect 504328 370387 504448 370553
rect 504328 370353 504371 370387
rect 504405 370353 504448 370387
rect 504328 370187 504448 370353
rect 504328 370153 504371 370187
rect 504405 370153 504448 370187
rect 504328 369987 504448 370153
rect 504328 369953 504371 369987
rect 504405 369953 504448 369987
rect 504328 369787 504448 369953
rect 504328 369753 504371 369787
rect 504405 369753 504448 369787
rect 504328 369587 504448 369753
rect 504328 369553 504371 369587
rect 504405 369553 504448 369587
rect 504328 369387 504448 369553
rect 504328 369353 504371 369387
rect 504405 369353 504448 369387
rect 504328 369187 504448 369353
rect 504328 369153 504371 369187
rect 504405 369153 504448 369187
rect 504328 368987 504448 369153
rect 504328 368953 504371 368987
rect 504405 368953 504448 368987
rect 504328 368787 504448 368953
rect 504328 368753 504371 368787
rect 504405 368753 504448 368787
rect 504328 368587 504448 368753
rect 504328 368553 504371 368587
rect 504405 368553 504448 368587
rect 504328 368387 504448 368553
rect 504328 368353 504371 368387
rect 504405 368353 504448 368387
rect 504328 368187 504448 368353
rect 504328 368153 504371 368187
rect 504405 368153 504448 368187
rect 504328 367987 504448 368153
rect 504328 367953 504371 367987
rect 504405 367953 504448 367987
rect 504328 367787 504448 367953
rect 504328 367753 504371 367787
rect 504405 367753 504448 367787
rect 504328 367587 504448 367753
rect 504328 367553 504371 367587
rect 504405 367553 504448 367587
rect 504328 367387 504448 367553
rect 504328 367353 504371 367387
rect 504405 367353 504448 367387
rect 504328 367187 504448 367353
rect 504328 367153 504371 367187
rect 504405 367153 504448 367187
rect 504328 366987 504448 367153
rect 504328 366953 504371 366987
rect 504405 366953 504448 366987
rect 504328 366787 504448 366953
rect 504328 366753 504371 366787
rect 504405 366753 504448 366787
rect 504328 366587 504448 366753
rect 504328 366553 504371 366587
rect 504405 366553 504448 366587
rect 504328 366387 504448 366553
rect 504328 366353 504371 366387
rect 504405 366353 504448 366387
rect 504328 366187 504448 366353
rect 504328 366153 504371 366187
rect 504405 366153 504448 366187
rect 504328 365987 504448 366153
rect 504328 365953 504371 365987
rect 504405 365953 504448 365987
rect 504328 365787 504448 365953
rect 504328 365753 504371 365787
rect 504405 365753 504448 365787
rect 504328 365587 504448 365753
rect 504328 365553 504371 365587
rect 504405 365553 504448 365587
rect 504328 365387 504448 365553
rect 504328 365353 504371 365387
rect 504405 365353 504448 365387
rect 504328 365187 504448 365353
rect 504328 365153 504371 365187
rect 504405 365153 504448 365187
rect 504328 364987 504448 365153
rect 504328 364953 504371 364987
rect 504405 364953 504448 364987
rect 504328 364787 504448 364953
rect 504328 364753 504371 364787
rect 504405 364753 504448 364787
rect 504328 364587 504448 364753
rect 504328 364553 504371 364587
rect 504405 364553 504448 364587
rect 504328 364387 504448 364553
rect 504328 364353 504371 364387
rect 504405 364353 504448 364387
rect 504328 364187 504448 364353
rect 504328 364153 504371 364187
rect 504405 364153 504448 364187
rect 504328 363987 504448 364153
rect 504328 363953 504371 363987
rect 504405 363953 504448 363987
rect 504328 363787 504448 363953
rect 504328 363753 504371 363787
rect 504405 363753 504448 363787
rect 504328 363587 504448 363753
rect 504328 363553 504371 363587
rect 504405 363553 504448 363587
rect 504328 363387 504448 363553
rect 504328 363353 504371 363387
rect 504405 363353 504448 363387
rect 504328 363187 504448 363353
rect 504328 363153 504371 363187
rect 504405 363153 504448 363187
rect 504328 362987 504448 363153
rect 504328 362953 504371 362987
rect 504405 362953 504448 362987
rect 504328 362787 504448 362953
rect 504328 362753 504371 362787
rect 504405 362753 504448 362787
rect 504328 362587 504448 362753
rect 504328 362553 504371 362587
rect 504405 362553 504448 362587
rect 504328 361476 504448 362553
rect 504698 373124 504768 373144
rect 504698 373090 504704 373124
rect 504738 373090 504768 373124
rect 504698 373034 504768 373090
rect 504698 373000 504704 373034
rect 504738 373000 504768 373034
rect 504698 372970 504768 373000
rect 504872 372982 504924 372988
rect 504848 372970 504872 372980
rect 504698 372960 504872 372970
rect 504698 372944 504864 372960
rect 504698 372910 504704 372944
rect 504738 372942 504864 372944
rect 504738 372910 504768 372942
rect 504698 372854 504768 372910
rect 504698 372820 504704 372854
rect 504738 372820 504768 372854
rect 504698 372764 504768 372820
rect 504698 372730 504704 372764
rect 504738 372730 504768 372764
rect 504698 372674 504768 372730
rect 504698 372640 504704 372674
rect 504738 372640 504768 372674
rect 504698 372584 504768 372640
rect 504698 372550 504704 372584
rect 504738 372550 504768 372584
rect 504698 372494 504768 372550
rect 504698 372460 504704 372494
rect 504738 372460 504768 372494
rect 504698 372404 504768 372460
rect 504698 372370 504704 372404
rect 504738 372370 504768 372404
rect 504698 372314 504768 372370
rect 504698 372280 504704 372314
rect 504738 372280 504768 372314
rect 504698 372224 504768 372280
rect 504698 372190 504704 372224
rect 504738 372190 504768 372224
rect 504698 372134 504768 372190
rect 504698 372100 504704 372134
rect 504738 372100 504768 372134
rect 504698 372044 504768 372100
rect 504698 372010 504704 372044
rect 504738 372010 504768 372044
rect 504698 371954 504768 372010
rect 504698 371920 504704 371954
rect 504738 371920 504768 371954
rect 504698 371784 504768 371920
rect 504698 371750 504704 371784
rect 504738 371750 504768 371784
rect 504698 371694 504768 371750
rect 504698 371660 504704 371694
rect 504738 371660 504768 371694
rect 504698 371604 504768 371660
rect 504698 371570 504704 371604
rect 504738 371570 504768 371604
rect 504698 371514 504768 371570
rect 504698 371480 504704 371514
rect 504738 371480 504768 371514
rect 504698 371424 504768 371480
rect 504698 371390 504704 371424
rect 504738 371390 504768 371424
rect 504698 371334 504768 371390
rect 504698 371300 504704 371334
rect 504738 371300 504768 371334
rect 504698 371244 504768 371300
rect 504698 371210 504704 371244
rect 504738 371210 504768 371244
rect 504698 371154 504768 371210
rect 504698 371120 504704 371154
rect 504738 371120 504768 371154
rect 504698 371064 504768 371120
rect 504698 371030 504704 371064
rect 504738 371030 504768 371064
rect 504698 370974 504768 371030
rect 504698 370940 504704 370974
rect 504738 370940 504768 370974
rect 504698 370884 504768 370940
rect 504698 370850 504704 370884
rect 504738 370850 504768 370884
rect 504698 370794 504768 370850
rect 504698 370760 504704 370794
rect 504738 370760 504768 370794
rect 504698 370704 504768 370760
rect 504698 370670 504704 370704
rect 504738 370670 504768 370704
rect 504698 370614 504768 370670
rect 504698 370580 504704 370614
rect 504738 370580 504768 370614
rect 504698 370444 504768 370580
rect 504698 370410 504704 370444
rect 504738 370410 504768 370444
rect 504698 370354 504768 370410
rect 504698 370320 504704 370354
rect 504738 370320 504768 370354
rect 504698 370264 504768 370320
rect 504698 370230 504704 370264
rect 504738 370230 504768 370264
rect 504698 370174 504768 370230
rect 504698 370140 504704 370174
rect 504738 370140 504768 370174
rect 504698 370084 504768 370140
rect 504698 370050 504704 370084
rect 504738 370050 504768 370084
rect 504698 369994 504768 370050
rect 504698 369960 504704 369994
rect 504738 369960 504768 369994
rect 504698 369904 504768 369960
rect 504698 369870 504704 369904
rect 504738 369870 504768 369904
rect 504698 369814 504768 369870
rect 504698 369780 504704 369814
rect 504738 369780 504768 369814
rect 504698 369724 504768 369780
rect 504698 369690 504704 369724
rect 504738 369690 504768 369724
rect 504698 369634 504768 369690
rect 504698 369600 504704 369634
rect 504738 369600 504768 369634
rect 504698 369544 504768 369600
rect 504698 369510 504704 369544
rect 504738 369510 504768 369544
rect 504698 369454 504768 369510
rect 504698 369420 504704 369454
rect 504738 369420 504768 369454
rect 504698 369364 504768 369420
rect 504698 369330 504704 369364
rect 504738 369330 504768 369364
rect 504698 369274 504768 369330
rect 504698 369240 504704 369274
rect 504738 369240 504768 369274
rect 504698 369104 504768 369240
rect 504698 369070 504704 369104
rect 504738 369070 504768 369104
rect 504698 369014 504768 369070
rect 504698 368980 504704 369014
rect 504738 368980 504768 369014
rect 504698 368924 504768 368980
rect 504698 368890 504704 368924
rect 504738 368890 504768 368924
rect 504698 368834 504768 368890
rect 504698 368800 504704 368834
rect 504738 368800 504768 368834
rect 504698 368744 504768 368800
rect 504698 368710 504704 368744
rect 504738 368710 504768 368744
rect 504698 368654 504768 368710
rect 504698 368620 504704 368654
rect 504738 368620 504768 368654
rect 504698 368564 504768 368620
rect 504698 368530 504704 368564
rect 504738 368530 504768 368564
rect 504698 368474 504768 368530
rect 504698 368440 504704 368474
rect 504738 368440 504768 368474
rect 504698 368384 504768 368440
rect 504698 368350 504704 368384
rect 504738 368350 504768 368384
rect 504698 368294 504768 368350
rect 504698 368260 504704 368294
rect 504738 368260 504768 368294
rect 504698 368204 504768 368260
rect 504698 368170 504704 368204
rect 504738 368170 504768 368204
rect 504698 368114 504768 368170
rect 504698 368080 504704 368114
rect 504738 368080 504768 368114
rect 504698 368024 504768 368080
rect 504698 367990 504704 368024
rect 504738 367990 504768 368024
rect 504698 367934 504768 367990
rect 504698 367900 504704 367934
rect 504738 367900 504768 367934
rect 504698 367764 504768 367900
rect 504698 367730 504704 367764
rect 504738 367730 504768 367764
rect 504698 367674 504768 367730
rect 504698 367640 504704 367674
rect 504738 367640 504768 367674
rect 504698 367584 504768 367640
rect 504698 367550 504704 367584
rect 504738 367550 504768 367584
rect 504698 367494 504768 367550
rect 504698 367460 504704 367494
rect 504738 367460 504768 367494
rect 504698 367404 504768 367460
rect 504698 367370 504704 367404
rect 504738 367370 504768 367404
rect 504698 367314 504768 367370
rect 504698 367280 504704 367314
rect 504738 367280 504768 367314
rect 504698 367224 504768 367280
rect 504698 367190 504704 367224
rect 504738 367190 504768 367224
rect 504698 367134 504768 367190
rect 504698 367100 504704 367134
rect 504738 367100 504768 367134
rect 504698 367044 504768 367100
rect 504698 367010 504704 367044
rect 504738 367010 504768 367044
rect 504698 366954 504768 367010
rect 504698 366920 504704 366954
rect 504738 366920 504768 366954
rect 504698 366864 504768 366920
rect 504698 366830 504704 366864
rect 504738 366830 504768 366864
rect 504698 366774 504768 366830
rect 504698 366740 504704 366774
rect 504738 366740 504768 366774
rect 504698 366684 504768 366740
rect 504698 366650 504704 366684
rect 504738 366650 504768 366684
rect 504698 366594 504768 366650
rect 504698 366560 504704 366594
rect 504738 366560 504768 366594
rect 504698 366424 504768 366560
rect 504698 366390 504704 366424
rect 504738 366390 504768 366424
rect 504698 366334 504768 366390
rect 504698 366300 504704 366334
rect 504738 366300 504768 366334
rect 504698 366244 504768 366300
rect 504698 366210 504704 366244
rect 504738 366210 504768 366244
rect 504698 366154 504768 366210
rect 504698 366120 504704 366154
rect 504738 366120 504768 366154
rect 504698 366064 504768 366120
rect 504698 366030 504704 366064
rect 504738 366030 504768 366064
rect 504698 365974 504768 366030
rect 504698 365940 504704 365974
rect 504738 365940 504768 365974
rect 504698 365884 504768 365940
rect 504698 365850 504704 365884
rect 504738 365850 504768 365884
rect 504698 365794 504768 365850
rect 504698 365760 504704 365794
rect 504738 365760 504768 365794
rect 504698 365704 504768 365760
rect 504698 365670 504704 365704
rect 504738 365670 504768 365704
rect 504698 365614 504768 365670
rect 504698 365580 504704 365614
rect 504738 365580 504768 365614
rect 504698 365524 504768 365580
rect 504698 365490 504704 365524
rect 504738 365490 504768 365524
rect 504698 365434 504768 365490
rect 504698 365400 504704 365434
rect 504738 365400 504768 365434
rect 504698 365344 504768 365400
rect 504698 365310 504704 365344
rect 504738 365310 504768 365344
rect 504698 365254 504768 365310
rect 504698 365220 504704 365254
rect 504738 365220 504768 365254
rect 504698 365084 504768 365220
rect 504698 365050 504704 365084
rect 504738 365050 504768 365084
rect 504698 364994 504768 365050
rect 504698 364960 504704 364994
rect 504738 364960 504768 364994
rect 504698 364904 504768 364960
rect 504698 364870 504704 364904
rect 504738 364870 504768 364904
rect 504698 364814 504768 364870
rect 504698 364780 504704 364814
rect 504738 364780 504768 364814
rect 504698 364724 504768 364780
rect 504698 364690 504704 364724
rect 504738 364690 504768 364724
rect 504698 364634 504768 364690
rect 504698 364600 504704 364634
rect 504738 364600 504768 364634
rect 504698 364544 504768 364600
rect 504698 364510 504704 364544
rect 504738 364510 504768 364544
rect 504698 364454 504768 364510
rect 504698 364420 504704 364454
rect 504738 364420 504768 364454
rect 504698 364364 504768 364420
rect 504698 364330 504704 364364
rect 504738 364330 504768 364364
rect 504698 364274 504768 364330
rect 504698 364240 504704 364274
rect 504738 364240 504768 364274
rect 504698 364184 504768 364240
rect 504698 364150 504704 364184
rect 504738 364150 504768 364184
rect 504698 364094 504768 364150
rect 504698 364060 504704 364094
rect 504738 364060 504768 364094
rect 504698 364004 504768 364060
rect 504698 363970 504704 364004
rect 504738 363970 504768 364004
rect 504698 363914 504768 363970
rect 504698 363880 504704 363914
rect 504738 363880 504768 363914
rect 504698 363744 504768 363880
rect 504698 363710 504704 363744
rect 504738 363710 504768 363744
rect 504698 363654 504768 363710
rect 504698 363620 504704 363654
rect 504738 363620 504768 363654
rect 504698 363564 504768 363620
rect 504698 363530 504704 363564
rect 504738 363530 504768 363564
rect 504698 363474 504768 363530
rect 504698 363440 504704 363474
rect 504738 363440 504768 363474
rect 504698 363384 504768 363440
rect 504698 363350 504704 363384
rect 504738 363350 504768 363384
rect 504698 363294 504768 363350
rect 504698 363260 504704 363294
rect 504738 363260 504768 363294
rect 504698 363204 504768 363260
rect 504698 363170 504704 363204
rect 504738 363170 504768 363204
rect 504698 363114 504768 363170
rect 504698 363080 504704 363114
rect 504738 363080 504768 363114
rect 504698 363024 504768 363080
rect 504698 362990 504704 363024
rect 504738 362990 504768 363024
rect 504698 362934 504768 362990
rect 504698 362900 504704 362934
rect 504738 362900 504768 362934
rect 504698 362844 504768 362900
rect 504698 362810 504704 362844
rect 504738 362810 504768 362844
rect 504698 362754 504768 362810
rect 504698 362720 504704 362754
rect 504738 362720 504768 362754
rect 504698 362664 504768 362720
rect 504698 362630 504704 362664
rect 504738 362630 504768 362664
rect 504848 372926 504864 372942
rect 504898 372926 504924 372930
rect 504848 372924 504924 372926
rect 506208 372987 506328 374865
rect 506208 372982 506251 372987
rect 506208 372930 506232 372982
rect 506285 372953 506328 372987
rect 506284 372930 506328 372953
rect 504848 372870 504918 372924
rect 504848 372836 504864 372870
rect 504898 372836 504918 372870
rect 504848 372780 504918 372836
rect 504848 372746 504864 372780
rect 504898 372746 504918 372780
rect 504848 372690 504918 372746
rect 504848 372656 504864 372690
rect 504898 372656 504918 372690
rect 504848 372600 504918 372656
rect 504848 372566 504864 372600
rect 504898 372566 504918 372600
rect 504848 372510 504918 372566
rect 504848 372476 504864 372510
rect 504898 372476 504918 372510
rect 504848 372420 504918 372476
rect 504848 372386 504864 372420
rect 504898 372386 504918 372420
rect 504848 372330 504918 372386
rect 504848 372296 504864 372330
rect 504898 372296 504918 372330
rect 504848 372240 504918 372296
rect 504848 372206 504864 372240
rect 504898 372206 504918 372240
rect 504848 372150 504918 372206
rect 504848 372116 504864 372150
rect 504898 372116 504918 372150
rect 504848 372060 504918 372116
rect 504848 372026 504864 372060
rect 504898 372026 504918 372060
rect 504848 371620 504918 372026
rect 504848 371586 504864 371620
rect 504898 371586 504918 371620
rect 504848 371530 504918 371586
rect 504848 371496 504864 371530
rect 504898 371496 504918 371530
rect 504848 371440 504918 371496
rect 504848 371406 504864 371440
rect 504898 371406 504918 371440
rect 504848 371350 504918 371406
rect 504848 371316 504864 371350
rect 504898 371316 504918 371350
rect 504848 371260 504918 371316
rect 504848 371226 504864 371260
rect 504898 371226 504918 371260
rect 504848 371170 504918 371226
rect 504848 371136 504864 371170
rect 504898 371136 504918 371170
rect 504848 371080 504918 371136
rect 504848 371046 504864 371080
rect 504898 371046 504918 371080
rect 504848 370990 504918 371046
rect 504848 370956 504864 370990
rect 504898 370956 504918 370990
rect 504848 370900 504918 370956
rect 504848 370866 504864 370900
rect 504898 370866 504918 370900
rect 504848 370810 504918 370866
rect 504848 370776 504864 370810
rect 504898 370776 504918 370810
rect 504848 370720 504918 370776
rect 504848 370686 504864 370720
rect 504898 370686 504918 370720
rect 504848 370280 504918 370686
rect 504848 370246 504864 370280
rect 504898 370246 504918 370280
rect 504848 370190 504918 370246
rect 504848 370156 504864 370190
rect 504898 370156 504918 370190
rect 504848 370100 504918 370156
rect 504848 370066 504864 370100
rect 504898 370066 504918 370100
rect 504848 370010 504918 370066
rect 504848 369976 504864 370010
rect 504898 369976 504918 370010
rect 504848 369920 504918 369976
rect 504848 369886 504864 369920
rect 504898 369886 504918 369920
rect 504848 369830 504918 369886
rect 504848 369796 504864 369830
rect 504898 369796 504918 369830
rect 504848 369740 504918 369796
rect 504848 369706 504864 369740
rect 504898 369706 504918 369740
rect 504848 369650 504918 369706
rect 504848 369616 504864 369650
rect 504898 369616 504918 369650
rect 504848 369560 504918 369616
rect 504848 369526 504864 369560
rect 504898 369526 504918 369560
rect 504848 369470 504918 369526
rect 504848 369436 504864 369470
rect 504898 369436 504918 369470
rect 504848 369380 504918 369436
rect 504848 369346 504864 369380
rect 504898 369346 504918 369380
rect 504848 368940 504918 369346
rect 504848 368906 504864 368940
rect 504898 368906 504918 368940
rect 504848 368850 504918 368906
rect 504848 368816 504864 368850
rect 504898 368816 504918 368850
rect 504848 368760 504918 368816
rect 504848 368726 504864 368760
rect 504898 368726 504918 368760
rect 504848 368670 504918 368726
rect 504848 368636 504864 368670
rect 504898 368636 504918 368670
rect 504848 368580 504918 368636
rect 504848 368546 504864 368580
rect 504898 368546 504918 368580
rect 504848 368490 504918 368546
rect 504848 368456 504864 368490
rect 504898 368456 504918 368490
rect 504848 368400 504918 368456
rect 504848 368366 504864 368400
rect 504898 368366 504918 368400
rect 504848 368310 504918 368366
rect 504848 368276 504864 368310
rect 504898 368276 504918 368310
rect 504848 368220 504918 368276
rect 504848 368186 504864 368220
rect 504898 368186 504918 368220
rect 504848 368130 504918 368186
rect 504848 368096 504864 368130
rect 504898 368096 504918 368130
rect 504848 368040 504918 368096
rect 504848 368006 504864 368040
rect 504898 368006 504918 368040
rect 504848 367600 504918 368006
rect 504848 367566 504864 367600
rect 504898 367566 504918 367600
rect 504848 367510 504918 367566
rect 504848 367476 504864 367510
rect 504898 367476 504918 367510
rect 504848 367420 504918 367476
rect 504848 367386 504864 367420
rect 504898 367386 504918 367420
rect 504848 367330 504918 367386
rect 504848 367296 504864 367330
rect 504898 367296 504918 367330
rect 504848 367240 504918 367296
rect 504848 367206 504864 367240
rect 504898 367206 504918 367240
rect 504848 367150 504918 367206
rect 504848 367116 504864 367150
rect 504898 367116 504918 367150
rect 504848 367060 504918 367116
rect 504848 367026 504864 367060
rect 504898 367026 504918 367060
rect 504848 366970 504918 367026
rect 504848 366936 504864 366970
rect 504898 366936 504918 366970
rect 504848 366880 504918 366936
rect 504848 366846 504864 366880
rect 504898 366846 504918 366880
rect 504848 366790 504918 366846
rect 504848 366756 504864 366790
rect 504898 366756 504918 366790
rect 504848 366700 504918 366756
rect 504848 366666 504864 366700
rect 504898 366666 504918 366700
rect 504848 366260 504918 366666
rect 504848 366226 504864 366260
rect 504898 366226 504918 366260
rect 504848 366170 504918 366226
rect 504848 366136 504864 366170
rect 504898 366136 504918 366170
rect 504848 366080 504918 366136
rect 504848 366046 504864 366080
rect 504898 366046 504918 366080
rect 504848 365990 504918 366046
rect 504848 365956 504864 365990
rect 504898 365956 504918 365990
rect 504848 365900 504918 365956
rect 504848 365866 504864 365900
rect 504898 365866 504918 365900
rect 504848 365810 504918 365866
rect 504848 365776 504864 365810
rect 504898 365776 504918 365810
rect 504848 365720 504918 365776
rect 504848 365686 504864 365720
rect 504898 365686 504918 365720
rect 504848 365630 504918 365686
rect 504848 365596 504864 365630
rect 504898 365596 504918 365630
rect 504848 365540 504918 365596
rect 504848 365506 504864 365540
rect 504898 365506 504918 365540
rect 504848 365450 504918 365506
rect 504848 365416 504864 365450
rect 504898 365416 504918 365450
rect 504848 365360 504918 365416
rect 504848 365326 504864 365360
rect 504898 365326 504918 365360
rect 504848 364920 504918 365326
rect 504848 364886 504864 364920
rect 504898 364886 504918 364920
rect 504848 364830 504918 364886
rect 504848 364796 504864 364830
rect 504898 364796 504918 364830
rect 504848 364740 504918 364796
rect 504848 364706 504864 364740
rect 504898 364706 504918 364740
rect 504848 364650 504918 364706
rect 504848 364616 504864 364650
rect 504898 364616 504918 364650
rect 504848 364560 504918 364616
rect 504848 364526 504864 364560
rect 504898 364526 504918 364560
rect 504848 364470 504918 364526
rect 504848 364436 504864 364470
rect 504898 364436 504918 364470
rect 504848 364380 504918 364436
rect 504848 364346 504864 364380
rect 504898 364346 504918 364380
rect 504848 364290 504918 364346
rect 504848 364256 504864 364290
rect 504898 364256 504918 364290
rect 504848 364200 504918 364256
rect 504848 364166 504864 364200
rect 504898 364166 504918 364200
rect 504848 364110 504918 364166
rect 504848 364076 504864 364110
rect 504898 364076 504918 364110
rect 504848 364020 504918 364076
rect 504848 363986 504864 364020
rect 504898 363986 504918 364020
rect 504848 363580 504918 363986
rect 504848 363546 504864 363580
rect 504898 363546 504918 363580
rect 504848 363490 504918 363546
rect 504848 363456 504864 363490
rect 504898 363456 504918 363490
rect 504848 363400 504918 363456
rect 504848 363366 504864 363400
rect 504898 363366 504918 363400
rect 504848 363310 504918 363366
rect 504848 363276 504864 363310
rect 504898 363276 504918 363310
rect 504848 363220 504918 363276
rect 504848 363186 504864 363220
rect 504898 363186 504918 363220
rect 504848 363130 504918 363186
rect 504848 363096 504864 363130
rect 504898 363096 504918 363130
rect 504848 363040 504918 363096
rect 504848 363006 504864 363040
rect 504898 363006 504918 363040
rect 504848 362950 504918 363006
rect 504848 362916 504864 362950
rect 504898 362916 504918 362950
rect 504848 362860 504918 362916
rect 504848 362826 504864 362860
rect 504898 362826 504918 362860
rect 504848 362770 504918 362826
rect 505022 372798 505634 372806
rect 505022 372774 505552 372798
rect 505022 372740 505068 372774
rect 505102 372740 505168 372774
rect 505202 372740 505268 372774
rect 505302 372740 505368 372774
rect 505402 372740 505468 372774
rect 505502 372746 505552 372774
rect 505604 372746 505634 372798
rect 505502 372740 505568 372746
rect 505602 372740 505634 372746
rect 505022 372674 505634 372740
rect 505022 372640 505068 372674
rect 505102 372640 505168 372674
rect 505202 372640 505268 372674
rect 505302 372640 505368 372674
rect 505402 372640 505468 372674
rect 505502 372640 505568 372674
rect 505602 372640 505634 372674
rect 505022 372574 505634 372640
rect 505022 372540 505068 372574
rect 505102 372540 505168 372574
rect 505202 372540 505268 372574
rect 505302 372540 505368 372574
rect 505402 372540 505468 372574
rect 505502 372540 505568 372574
rect 505602 372540 505634 372574
rect 505022 372474 505634 372540
rect 505022 372440 505068 372474
rect 505102 372440 505168 372474
rect 505202 372440 505268 372474
rect 505302 372440 505368 372474
rect 505402 372440 505468 372474
rect 505502 372440 505568 372474
rect 505602 372440 505634 372474
rect 505022 372374 505634 372440
rect 505022 372340 505068 372374
rect 505102 372340 505168 372374
rect 505202 372340 505268 372374
rect 505302 372340 505368 372374
rect 505402 372340 505468 372374
rect 505502 372340 505568 372374
rect 505602 372340 505634 372374
rect 505022 372274 505634 372340
rect 505022 372240 505068 372274
rect 505102 372240 505168 372274
rect 505202 372240 505268 372274
rect 505302 372240 505368 372274
rect 505402 372240 505468 372274
rect 505502 372240 505568 372274
rect 505602 372240 505634 372274
rect 505022 371434 505634 372240
rect 505022 371400 505068 371434
rect 505102 371400 505168 371434
rect 505202 371400 505268 371434
rect 505302 371400 505368 371434
rect 505402 371400 505468 371434
rect 505502 371400 505568 371434
rect 505602 371400 505634 371434
rect 505022 371334 505634 371400
rect 505022 371300 505068 371334
rect 505102 371300 505168 371334
rect 505202 371300 505268 371334
rect 505302 371300 505368 371334
rect 505402 371300 505468 371334
rect 505502 371300 505568 371334
rect 505602 371300 505634 371334
rect 505022 371234 505634 371300
rect 505022 371200 505068 371234
rect 505102 371200 505168 371234
rect 505202 371200 505268 371234
rect 505302 371200 505368 371234
rect 505402 371200 505468 371234
rect 505502 371200 505568 371234
rect 505602 371200 505634 371234
rect 505022 371134 505634 371200
rect 505022 371100 505068 371134
rect 505102 371100 505168 371134
rect 505202 371100 505268 371134
rect 505302 371100 505368 371134
rect 505402 371100 505468 371134
rect 505502 371100 505568 371134
rect 505602 371100 505634 371134
rect 505022 371034 505634 371100
rect 505022 371000 505068 371034
rect 505102 371000 505168 371034
rect 505202 371000 505268 371034
rect 505302 371000 505368 371034
rect 505402 371000 505468 371034
rect 505502 371000 505568 371034
rect 505602 371000 505634 371034
rect 505022 370934 505634 371000
rect 505022 370900 505068 370934
rect 505102 370900 505168 370934
rect 505202 370900 505268 370934
rect 505302 370900 505368 370934
rect 505402 370900 505468 370934
rect 505502 370900 505568 370934
rect 505602 370900 505634 370934
rect 505022 370094 505634 370900
rect 505022 370060 505068 370094
rect 505102 370060 505168 370094
rect 505202 370060 505268 370094
rect 505302 370060 505368 370094
rect 505402 370060 505468 370094
rect 505502 370060 505568 370094
rect 505602 370060 505634 370094
rect 505022 369994 505634 370060
rect 505022 369960 505068 369994
rect 505102 369960 505168 369994
rect 505202 369960 505268 369994
rect 505302 369960 505368 369994
rect 505402 369960 505468 369994
rect 505502 369960 505568 369994
rect 505602 369960 505634 369994
rect 505022 369894 505634 369960
rect 505022 369860 505068 369894
rect 505102 369860 505168 369894
rect 505202 369860 505268 369894
rect 505302 369860 505368 369894
rect 505402 369860 505468 369894
rect 505502 369860 505568 369894
rect 505602 369860 505634 369894
rect 505022 369794 505634 369860
rect 505022 369760 505068 369794
rect 505102 369760 505168 369794
rect 505202 369760 505268 369794
rect 505302 369760 505368 369794
rect 505402 369760 505468 369794
rect 505502 369760 505568 369794
rect 505602 369760 505634 369794
rect 505022 369694 505634 369760
rect 505022 369660 505068 369694
rect 505102 369660 505168 369694
rect 505202 369660 505268 369694
rect 505302 369660 505368 369694
rect 505402 369660 505468 369694
rect 505502 369660 505568 369694
rect 505602 369660 505634 369694
rect 505022 369594 505634 369660
rect 505022 369560 505068 369594
rect 505102 369560 505168 369594
rect 505202 369560 505268 369594
rect 505302 369560 505368 369594
rect 505402 369560 505468 369594
rect 505502 369560 505568 369594
rect 505602 369560 505634 369594
rect 505022 368754 505634 369560
rect 505022 368720 505068 368754
rect 505102 368720 505168 368754
rect 505202 368720 505268 368754
rect 505302 368720 505368 368754
rect 505402 368720 505468 368754
rect 505502 368720 505568 368754
rect 505602 368720 505634 368754
rect 505022 368654 505634 368720
rect 505022 368620 505068 368654
rect 505102 368620 505168 368654
rect 505202 368620 505268 368654
rect 505302 368620 505368 368654
rect 505402 368620 505468 368654
rect 505502 368620 505568 368654
rect 505602 368620 505634 368654
rect 505022 368554 505634 368620
rect 505022 368520 505068 368554
rect 505102 368520 505168 368554
rect 505202 368520 505268 368554
rect 505302 368520 505368 368554
rect 505402 368520 505468 368554
rect 505502 368520 505568 368554
rect 505602 368520 505634 368554
rect 505022 368454 505634 368520
rect 505022 368420 505068 368454
rect 505102 368420 505168 368454
rect 505202 368420 505268 368454
rect 505302 368420 505368 368454
rect 505402 368420 505468 368454
rect 505502 368420 505568 368454
rect 505602 368420 505634 368454
rect 505022 368354 505634 368420
rect 505022 368320 505068 368354
rect 505102 368320 505168 368354
rect 505202 368320 505268 368354
rect 505302 368320 505368 368354
rect 505402 368320 505468 368354
rect 505502 368320 505568 368354
rect 505602 368320 505634 368354
rect 505022 368254 505634 368320
rect 505022 368220 505068 368254
rect 505102 368220 505168 368254
rect 505202 368220 505268 368254
rect 505302 368220 505368 368254
rect 505402 368220 505468 368254
rect 505502 368220 505568 368254
rect 505602 368220 505634 368254
rect 505022 367414 505634 368220
rect 505022 367380 505068 367414
rect 505102 367380 505168 367414
rect 505202 367380 505268 367414
rect 505302 367380 505368 367414
rect 505402 367380 505468 367414
rect 505502 367380 505568 367414
rect 505602 367380 505634 367414
rect 505022 367314 505634 367380
rect 505022 367280 505068 367314
rect 505102 367280 505168 367314
rect 505202 367280 505268 367314
rect 505302 367280 505368 367314
rect 505402 367280 505468 367314
rect 505502 367280 505568 367314
rect 505602 367280 505634 367314
rect 505022 367214 505634 367280
rect 505022 367180 505068 367214
rect 505102 367180 505168 367214
rect 505202 367180 505268 367214
rect 505302 367180 505368 367214
rect 505402 367180 505468 367214
rect 505502 367180 505568 367214
rect 505602 367180 505634 367214
rect 505022 367114 505634 367180
rect 505022 367080 505068 367114
rect 505102 367080 505168 367114
rect 505202 367080 505268 367114
rect 505302 367080 505368 367114
rect 505402 367080 505468 367114
rect 505502 367080 505568 367114
rect 505602 367080 505634 367114
rect 505022 367014 505634 367080
rect 505022 366980 505068 367014
rect 505102 366980 505168 367014
rect 505202 366980 505268 367014
rect 505302 366980 505368 367014
rect 505402 366980 505468 367014
rect 505502 366980 505568 367014
rect 505602 366980 505634 367014
rect 505022 366914 505634 366980
rect 505022 366880 505068 366914
rect 505102 366880 505168 366914
rect 505202 366880 505268 366914
rect 505302 366880 505368 366914
rect 505402 366880 505468 366914
rect 505502 366880 505568 366914
rect 505602 366880 505634 366914
rect 505022 366074 505634 366880
rect 505022 366040 505068 366074
rect 505102 366040 505168 366074
rect 505202 366040 505268 366074
rect 505302 366040 505368 366074
rect 505402 366040 505468 366074
rect 505502 366040 505568 366074
rect 505602 366040 505634 366074
rect 505022 365974 505634 366040
rect 505022 365940 505068 365974
rect 505102 365940 505168 365974
rect 505202 365940 505268 365974
rect 505302 365940 505368 365974
rect 505402 365940 505468 365974
rect 505502 365940 505568 365974
rect 505602 365940 505634 365974
rect 505022 365874 505634 365940
rect 505022 365840 505068 365874
rect 505102 365840 505168 365874
rect 505202 365840 505268 365874
rect 505302 365840 505368 365874
rect 505402 365840 505468 365874
rect 505502 365840 505568 365874
rect 505602 365840 505634 365874
rect 505022 365774 505634 365840
rect 505022 365740 505068 365774
rect 505102 365740 505168 365774
rect 505202 365740 505268 365774
rect 505302 365740 505368 365774
rect 505402 365740 505468 365774
rect 505502 365740 505568 365774
rect 505602 365740 505634 365774
rect 505022 365674 505634 365740
rect 505022 365640 505068 365674
rect 505102 365640 505168 365674
rect 505202 365640 505268 365674
rect 505302 365640 505368 365674
rect 505402 365640 505468 365674
rect 505502 365640 505568 365674
rect 505602 365640 505634 365674
rect 505022 365574 505634 365640
rect 505022 365540 505068 365574
rect 505102 365540 505168 365574
rect 505202 365540 505268 365574
rect 505302 365540 505368 365574
rect 505402 365540 505468 365574
rect 505502 365540 505568 365574
rect 505602 365540 505634 365574
rect 505022 364734 505634 365540
rect 505022 364700 505068 364734
rect 505102 364700 505168 364734
rect 505202 364700 505268 364734
rect 505302 364700 505368 364734
rect 505402 364700 505468 364734
rect 505502 364700 505568 364734
rect 505602 364700 505634 364734
rect 505022 364634 505634 364700
rect 505022 364600 505068 364634
rect 505102 364600 505168 364634
rect 505202 364600 505268 364634
rect 505302 364600 505368 364634
rect 505402 364600 505468 364634
rect 505502 364600 505568 364634
rect 505602 364600 505634 364634
rect 505022 364534 505634 364600
rect 505022 364500 505068 364534
rect 505102 364500 505168 364534
rect 505202 364500 505268 364534
rect 505302 364500 505368 364534
rect 505402 364500 505468 364534
rect 505502 364500 505568 364534
rect 505602 364500 505634 364534
rect 505022 364434 505634 364500
rect 505022 364400 505068 364434
rect 505102 364400 505168 364434
rect 505202 364400 505268 364434
rect 505302 364400 505368 364434
rect 505402 364400 505468 364434
rect 505502 364400 505568 364434
rect 505602 364400 505634 364434
rect 505022 364334 505634 364400
rect 505022 364300 505068 364334
rect 505102 364300 505168 364334
rect 505202 364300 505268 364334
rect 505302 364300 505368 364334
rect 505402 364300 505468 364334
rect 505502 364300 505568 364334
rect 505602 364300 505634 364334
rect 505022 364234 505634 364300
rect 505022 364200 505068 364234
rect 505102 364200 505168 364234
rect 505202 364200 505268 364234
rect 505302 364200 505368 364234
rect 505402 364200 505468 364234
rect 505502 364200 505568 364234
rect 505602 364200 505634 364234
rect 505022 363394 505634 364200
rect 505022 363360 505068 363394
rect 505102 363360 505168 363394
rect 505202 363360 505268 363394
rect 505302 363360 505368 363394
rect 505402 363360 505468 363394
rect 505502 363360 505568 363394
rect 505602 363360 505634 363394
rect 505022 363294 505634 363360
rect 505022 363260 505068 363294
rect 505102 363260 505168 363294
rect 505202 363260 505268 363294
rect 505302 363260 505368 363294
rect 505402 363260 505468 363294
rect 505502 363260 505568 363294
rect 505602 363260 505634 363294
rect 505022 363194 505634 363260
rect 505022 363160 505068 363194
rect 505102 363160 505168 363194
rect 505202 363160 505268 363194
rect 505302 363160 505368 363194
rect 505402 363160 505468 363194
rect 505502 363160 505568 363194
rect 505602 363160 505634 363194
rect 505022 363094 505634 363160
rect 505022 363060 505068 363094
rect 505102 363060 505168 363094
rect 505202 363060 505268 363094
rect 505302 363060 505368 363094
rect 505402 363060 505468 363094
rect 505502 363060 505568 363094
rect 505602 363060 505634 363094
rect 505022 362994 505634 363060
rect 505022 362960 505068 362994
rect 505102 362960 505168 362994
rect 505202 362960 505268 362994
rect 505302 362960 505368 362994
rect 505402 362960 505468 362994
rect 505502 362960 505568 362994
rect 505602 362960 505634 362994
rect 505022 362894 505634 362960
rect 505022 362860 505068 362894
rect 505102 362860 505168 362894
rect 505202 362860 505268 362894
rect 505302 362860 505368 362894
rect 505402 362860 505468 362894
rect 505502 362860 505568 362894
rect 505602 362860 505634 362894
rect 505022 362814 505634 362860
rect 506208 372787 506328 372930
rect 506208 372753 506251 372787
rect 506285 372753 506328 372787
rect 506208 372587 506328 372753
rect 506208 372553 506251 372587
rect 506285 372553 506328 372587
rect 506208 372387 506328 372553
rect 506208 372353 506251 372387
rect 506285 372353 506328 372387
rect 506208 372187 506328 372353
rect 506208 372153 506251 372187
rect 506285 372153 506328 372187
rect 506208 371987 506328 372153
rect 506208 371953 506251 371987
rect 506285 371953 506328 371987
rect 506208 371787 506328 371953
rect 506208 371753 506251 371787
rect 506285 371753 506328 371787
rect 506208 371587 506328 371753
rect 506208 371553 506251 371587
rect 506285 371553 506328 371587
rect 506208 371387 506328 371553
rect 506208 371353 506251 371387
rect 506285 371353 506328 371387
rect 506208 371187 506328 371353
rect 506208 371153 506251 371187
rect 506285 371153 506328 371187
rect 506208 370987 506328 371153
rect 506208 370953 506251 370987
rect 506285 370953 506328 370987
rect 506208 370787 506328 370953
rect 506208 370753 506251 370787
rect 506285 370753 506328 370787
rect 506208 370587 506328 370753
rect 506208 370553 506251 370587
rect 506285 370553 506328 370587
rect 506208 370387 506328 370553
rect 506208 370353 506251 370387
rect 506285 370353 506328 370387
rect 506208 370187 506328 370353
rect 506208 370153 506251 370187
rect 506285 370153 506328 370187
rect 506208 369987 506328 370153
rect 506208 369953 506251 369987
rect 506285 369953 506328 369987
rect 506208 369787 506328 369953
rect 506208 369753 506251 369787
rect 506285 369753 506328 369787
rect 506208 369587 506328 369753
rect 506208 369553 506251 369587
rect 506285 369553 506328 369587
rect 506208 369387 506328 369553
rect 506208 369353 506251 369387
rect 506285 369353 506328 369387
rect 506208 369187 506328 369353
rect 506208 369153 506251 369187
rect 506285 369153 506328 369187
rect 506208 368987 506328 369153
rect 506208 368953 506251 368987
rect 506285 368953 506328 368987
rect 506208 368787 506328 368953
rect 506208 368753 506251 368787
rect 506285 368753 506328 368787
rect 506208 368587 506328 368753
rect 506208 368553 506251 368587
rect 506285 368553 506328 368587
rect 506208 368387 506328 368553
rect 506208 368353 506251 368387
rect 506285 368353 506328 368387
rect 506208 368187 506328 368353
rect 506208 368153 506251 368187
rect 506285 368153 506328 368187
rect 506208 367987 506328 368153
rect 506208 367953 506251 367987
rect 506285 367953 506328 367987
rect 506208 367787 506328 367953
rect 506208 367753 506251 367787
rect 506285 367753 506328 367787
rect 506208 367587 506328 367753
rect 506208 367553 506251 367587
rect 506285 367553 506328 367587
rect 506208 367387 506328 367553
rect 506208 367353 506251 367387
rect 506285 367353 506328 367387
rect 506208 367187 506328 367353
rect 506208 367153 506251 367187
rect 506285 367153 506328 367187
rect 506208 366987 506328 367153
rect 506208 366953 506251 366987
rect 506285 366953 506328 366987
rect 506208 366787 506328 366953
rect 506208 366753 506251 366787
rect 506285 366753 506328 366787
rect 506208 366587 506328 366753
rect 506208 366553 506251 366587
rect 506285 366553 506328 366587
rect 506208 366387 506328 366553
rect 506208 366353 506251 366387
rect 506285 366353 506328 366387
rect 506208 366187 506328 366353
rect 506208 366153 506251 366187
rect 506285 366153 506328 366187
rect 506208 365987 506328 366153
rect 506208 365953 506251 365987
rect 506285 365953 506328 365987
rect 506208 365787 506328 365953
rect 506208 365753 506251 365787
rect 506285 365753 506328 365787
rect 506208 365587 506328 365753
rect 506208 365553 506251 365587
rect 506285 365553 506328 365587
rect 506208 365387 506328 365553
rect 506208 365353 506251 365387
rect 506285 365353 506328 365387
rect 506208 365187 506328 365353
rect 506208 365153 506251 365187
rect 506285 365153 506328 365187
rect 506208 364987 506328 365153
rect 506208 364953 506251 364987
rect 506285 364953 506328 364987
rect 506208 364787 506328 364953
rect 506208 364753 506251 364787
rect 506285 364753 506328 364787
rect 506208 364587 506328 364753
rect 506208 364553 506251 364587
rect 506285 364553 506328 364587
rect 506208 364387 506328 364553
rect 506208 364353 506251 364387
rect 506285 364353 506328 364387
rect 506208 364187 506328 364353
rect 506208 364153 506251 364187
rect 506285 364153 506328 364187
rect 506208 363987 506328 364153
rect 506208 363953 506251 363987
rect 506285 363953 506328 363987
rect 506208 363787 506328 363953
rect 506208 363753 506251 363787
rect 506285 363753 506328 363787
rect 506208 363587 506328 363753
rect 506208 363553 506251 363587
rect 506285 363553 506328 363587
rect 506208 363387 506328 363553
rect 506208 363353 506251 363387
rect 506285 363353 506328 363387
rect 506208 363187 506328 363353
rect 506208 363153 506251 363187
rect 506285 363153 506328 363187
rect 506208 362987 506328 363153
rect 506208 362953 506251 362987
rect 506285 362953 506328 362987
rect 504848 362736 504864 362770
rect 504898 362736 504918 362770
rect 504848 362680 504918 362736
rect 504848 362646 504864 362680
rect 504898 362646 504918 362680
rect 504848 362640 504918 362646
rect 506208 362787 506328 362953
rect 506208 362753 506251 362787
rect 506285 362753 506328 362787
rect 504698 362574 504768 362630
rect 504698 362540 504704 362574
rect 504738 362540 504768 362574
rect 504698 362476 504768 362540
rect 506208 362587 506328 362753
rect 506208 362553 506251 362587
rect 506285 362553 506328 362587
rect 504328 359888 504330 361476
rect 504446 359888 504448 361476
rect 504328 359866 504448 359888
rect 502448 357440 502450 359028
rect 502566 357440 502568 359028
rect 502448 357418 502568 357440
rect 506208 359028 506328 362553
rect 508088 411584 508208 411606
rect 508088 409996 508090 411584
rect 508206 409996 508208 411584
rect 508088 395507 508208 409996
rect 509360 398374 509412 398380
rect 509360 398316 509412 398322
rect 509372 395679 509400 398316
rect 508088 395473 508131 395507
rect 508165 395473 508208 395507
rect 508088 395307 508208 395473
rect 508088 395273 508131 395307
rect 508165 395273 508208 395307
rect 508088 395107 508208 395273
rect 508387 395671 508949 395679
rect 508387 395277 508399 395671
rect 508937 395277 508949 395671
rect 508387 395269 508949 395277
rect 509347 395671 509909 395679
rect 509347 395277 509359 395671
rect 509897 395277 509909 395671
rect 509347 395269 509909 395277
rect 509968 395507 510088 412444
rect 513728 414032 513848 414054
rect 513728 412444 513730 414032
rect 513846 412444 513848 414032
rect 509968 395473 510011 395507
rect 510045 395473 510088 395507
rect 509968 395307 510088 395473
rect 509968 395273 510011 395307
rect 510045 395273 510088 395307
rect 508088 395073 508131 395107
rect 508165 395073 508208 395107
rect 508088 394907 508208 395073
rect 508088 394873 508131 394907
rect 508165 394873 508208 394907
rect 508088 394707 508208 394873
rect 508088 394673 508131 394707
rect 508165 394673 508208 394707
rect 508088 394507 508208 394673
rect 508088 394473 508131 394507
rect 508165 394473 508208 394507
rect 508088 394307 508208 394473
rect 508088 394273 508131 394307
rect 508165 394273 508208 394307
rect 508088 394107 508208 394273
rect 508088 394073 508131 394107
rect 508165 394073 508208 394107
rect 508088 393907 508208 394073
rect 508088 393873 508131 393907
rect 508165 393873 508208 393907
rect 508088 393707 508208 393873
rect 508088 393673 508131 393707
rect 508165 393673 508208 393707
rect 509968 395107 510088 395273
rect 509968 395073 510011 395107
rect 510045 395073 510088 395107
rect 509968 394907 510088 395073
rect 509968 394873 510011 394907
rect 510045 394873 510088 394907
rect 509968 394707 510088 394873
rect 509968 394673 510011 394707
rect 510045 394673 510088 394707
rect 509968 394507 510088 394673
rect 509968 394473 510011 394507
rect 510045 394473 510088 394507
rect 509968 394307 510088 394473
rect 509968 394273 510011 394307
rect 510045 394273 510088 394307
rect 509968 394107 510088 394273
rect 509968 394073 510011 394107
rect 510045 394073 510088 394107
rect 509968 393907 510088 394073
rect 509968 393873 510011 393907
rect 510045 393873 510088 393907
rect 509968 393707 510088 393873
rect 508088 393507 508208 393673
rect 508949 393671 509913 393682
rect 508088 393473 508131 393507
rect 508165 393473 508208 393507
rect 508088 392761 508208 393473
rect 508387 393664 509913 393671
rect 508387 393270 508399 393664
rect 508937 393270 509359 393664
rect 509897 393270 509913 393664
rect 508387 393261 509913 393270
rect 508949 393250 509913 393261
rect 509968 393673 510011 393707
rect 510045 393673 510088 393707
rect 509968 393507 510088 393673
rect 509968 393473 510011 393507
rect 510045 393473 510088 393507
rect 508088 392727 508131 392761
rect 508165 392727 508208 392761
rect 508088 392561 508208 392727
rect 508088 392527 508131 392561
rect 508165 392527 508208 392561
rect 508088 392361 508208 392527
rect 508387 392926 508949 392934
rect 508387 392532 508399 392926
rect 508937 392532 508949 392926
rect 508387 392524 508949 392532
rect 509347 392926 509909 392934
rect 509347 392532 509359 392926
rect 509897 392566 509909 392926
rect 509968 392761 510088 393473
rect 509968 392727 510011 392761
rect 510045 392727 510088 392761
rect 509968 392566 510088 392727
rect 509897 392561 510088 392566
rect 509897 392538 510011 392561
rect 509897 392532 509909 392538
rect 509347 392524 509909 392532
rect 509968 392527 510011 392538
rect 510045 392527 510088 392561
rect 508088 392327 508131 392361
rect 508165 392327 508208 392361
rect 508088 392161 508208 392327
rect 508088 392127 508131 392161
rect 508165 392127 508208 392161
rect 508088 391961 508208 392127
rect 508088 391927 508131 391961
rect 508165 391927 508208 391961
rect 508088 391761 508208 391927
rect 508088 391727 508131 391761
rect 508165 391727 508208 391761
rect 508088 391561 508208 391727
rect 508088 391527 508131 391561
rect 508165 391527 508208 391561
rect 508088 391361 508208 391527
rect 508088 391327 508131 391361
rect 508165 391327 508208 391361
rect 508088 391161 508208 391327
rect 508088 391127 508131 391161
rect 508165 391127 508208 391161
rect 508088 390961 508208 391127
rect 508088 390927 508131 390961
rect 508165 390927 508208 390961
rect 508088 390761 508208 390927
rect 508088 390727 508131 390761
rect 508165 390727 508208 390761
rect 508088 390561 508208 390727
rect 508088 390527 508131 390561
rect 508165 390527 508208 390561
rect 508088 390361 508208 390527
rect 508896 390468 508924 392524
rect 509968 392361 510088 392527
rect 509968 392327 510011 392361
rect 510045 392327 510088 392361
rect 509968 392161 510088 392327
rect 509968 392127 510011 392161
rect 510045 392127 510088 392161
rect 509968 391961 510088 392127
rect 509968 391927 510011 391961
rect 510045 391927 510088 391961
rect 509968 391761 510088 391927
rect 509968 391727 510011 391761
rect 510045 391727 510088 391761
rect 509968 391561 510088 391727
rect 509968 391527 510011 391561
rect 510045 391527 510088 391561
rect 509968 391361 510088 391527
rect 509968 391327 510011 391361
rect 510045 391327 510088 391361
rect 509968 391161 510088 391327
rect 509968 391127 510011 391161
rect 510045 391127 510088 391161
rect 509968 390961 510088 391127
rect 509968 390927 510011 390961
rect 510045 390927 510088 390961
rect 509968 390761 510088 390927
rect 509968 390727 510011 390761
rect 510045 390727 510088 390761
rect 509968 390561 510088 390727
rect 509968 390527 510011 390561
rect 510045 390527 510088 390561
rect 508884 390462 508936 390468
rect 508884 390404 508936 390410
rect 508088 390327 508131 390361
rect 508165 390327 508208 390361
rect 508949 390352 509913 390363
rect 508088 390161 508208 390327
rect 508088 390127 508131 390161
rect 508165 390127 508208 390161
rect 508088 388567 508208 390127
rect 508387 390345 509913 390352
rect 508387 389951 508399 390345
rect 508937 389951 509359 390345
rect 509897 389951 509913 390345
rect 508387 389942 509913 389951
rect 508949 389931 509913 389942
rect 509968 390361 510088 390527
rect 509968 390327 510011 390361
rect 510045 390327 510088 390361
rect 509968 390161 510088 390327
rect 509968 390127 510011 390161
rect 510045 390127 510088 390161
rect 508088 388533 508131 388567
rect 508165 388533 508208 388567
rect 508088 388167 508208 388533
rect 508088 388133 508131 388167
rect 508165 388133 508208 388167
rect 508088 387767 508208 388133
rect 508088 387733 508131 387767
rect 508165 387733 508208 387767
rect 508088 387367 508208 387733
rect 508088 387333 508131 387367
rect 508165 387333 508208 387367
rect 508088 386967 508208 387333
rect 508088 386933 508131 386967
rect 508165 386933 508208 386967
rect 508088 386567 508208 386933
rect 508088 386533 508131 386567
rect 508165 386533 508208 386567
rect 508088 386167 508208 386533
rect 508088 386133 508131 386167
rect 508165 386133 508208 386167
rect 508088 385767 508208 386133
rect 508088 385733 508131 385767
rect 508165 385733 508208 385767
rect 508088 385367 508208 385733
rect 508088 385333 508131 385367
rect 508165 385333 508208 385367
rect 508088 384967 508208 385333
rect 508088 384933 508131 384967
rect 508165 384933 508208 384967
rect 508088 384567 508208 384933
rect 508088 384533 508131 384567
rect 508165 384533 508208 384567
rect 508088 384167 508208 384533
rect 508088 384133 508131 384167
rect 508165 384133 508208 384167
rect 508088 383767 508208 384133
rect 508088 383733 508131 383767
rect 508165 383733 508208 383767
rect 508088 383367 508208 383733
rect 508088 383333 508131 383367
rect 508165 383333 508208 383367
rect 508088 382967 508208 383333
rect 508088 382933 508131 382967
rect 508165 382933 508208 382967
rect 508088 382567 508208 382933
rect 508088 382533 508131 382567
rect 508165 382533 508208 382567
rect 508088 382167 508208 382533
rect 508088 382133 508131 382167
rect 508165 382133 508208 382167
rect 508088 381767 508208 382133
rect 508088 381733 508131 381767
rect 508165 381733 508208 381767
rect 508088 381538 508208 381733
rect 508088 381486 508136 381538
rect 508188 381486 508208 381538
rect 508088 381119 508208 381486
rect 508088 381085 508131 381119
rect 508165 381085 508208 381119
rect 508088 380719 508208 381085
rect 508088 380685 508131 380719
rect 508165 380685 508208 380719
rect 508088 380319 508208 380685
rect 508088 380285 508131 380319
rect 508165 380285 508208 380319
rect 508088 379919 508208 380285
rect 508088 379885 508131 379919
rect 508165 379885 508208 379919
rect 508088 379519 508208 379885
rect 508088 379485 508131 379519
rect 508165 379485 508208 379519
rect 508088 379119 508208 379485
rect 508088 379085 508131 379119
rect 508165 379085 508208 379119
rect 508088 378719 508208 379085
rect 508088 378685 508131 378719
rect 508165 378685 508208 378719
rect 508088 378319 508208 378685
rect 508088 378285 508131 378319
rect 508165 378285 508208 378319
rect 508088 377919 508208 378285
rect 508088 377885 508131 377919
rect 508165 377885 508208 377919
rect 508088 377519 508208 377885
rect 508088 377485 508131 377519
rect 508165 377485 508208 377519
rect 508088 377119 508208 377485
rect 508088 377085 508131 377119
rect 508165 377085 508208 377119
rect 508088 376719 508208 377085
rect 508088 376685 508131 376719
rect 508165 376685 508208 376719
rect 508088 376319 508208 376685
rect 508088 376285 508131 376319
rect 508165 376285 508208 376319
rect 508088 375919 508208 376285
rect 508088 375885 508131 375919
rect 508165 375885 508208 375919
rect 508088 375519 508208 375885
rect 508088 375485 508131 375519
rect 508165 375485 508208 375519
rect 508088 375119 508208 375485
rect 508088 375085 508131 375119
rect 508165 375085 508208 375119
rect 508088 374719 508208 375085
rect 508088 374685 508131 374719
rect 508165 374685 508208 374719
rect 508088 374319 508208 374685
rect 508088 374285 508131 374319
rect 508165 374285 508208 374319
rect 508088 372987 508208 374285
rect 509968 388567 510088 390127
rect 509968 388533 510011 388567
rect 510045 388533 510088 388567
rect 509968 388167 510088 388533
rect 509968 388133 510011 388167
rect 510045 388133 510088 388167
rect 509968 387767 510088 388133
rect 509968 387733 510011 387767
rect 510045 387733 510088 387767
rect 509968 387367 510088 387733
rect 509968 387333 510011 387367
rect 510045 387333 510088 387367
rect 509968 386967 510088 387333
rect 509968 386933 510011 386967
rect 510045 386933 510088 386967
rect 509968 386567 510088 386933
rect 509968 386533 510011 386567
rect 510045 386533 510088 386567
rect 509968 386167 510088 386533
rect 509968 386133 510011 386167
rect 510045 386133 510088 386167
rect 509968 385767 510088 386133
rect 509968 385733 510011 385767
rect 510045 385733 510088 385767
rect 509968 385367 510088 385733
rect 509968 385333 510011 385367
rect 510045 385333 510088 385367
rect 509968 384967 510088 385333
rect 509968 384933 510011 384967
rect 510045 384933 510088 384967
rect 509968 384567 510088 384933
rect 509968 384533 510011 384567
rect 510045 384533 510088 384567
rect 509968 384167 510088 384533
rect 509968 384133 510011 384167
rect 510045 384133 510088 384167
rect 509968 383767 510088 384133
rect 509968 383733 510011 383767
rect 510045 383733 510088 383767
rect 509968 383367 510088 383733
rect 509968 383333 510011 383367
rect 510045 383333 510088 383367
rect 509968 382967 510088 383333
rect 509968 382933 510011 382967
rect 510045 382933 510088 382967
rect 509968 382567 510088 382933
rect 509968 382533 510011 382567
rect 510045 382533 510088 382567
rect 509968 382167 510088 382533
rect 509968 382133 510011 382167
rect 510045 382133 510088 382167
rect 509968 381767 510088 382133
rect 509968 381733 510011 381767
rect 510045 381733 510088 381767
rect 509968 381119 510088 381733
rect 509968 381085 510011 381119
rect 510045 381085 510088 381119
rect 509968 380719 510088 381085
rect 509968 380685 510011 380719
rect 510045 380685 510088 380719
rect 509968 380319 510088 380685
rect 509968 380285 510011 380319
rect 510045 380285 510088 380319
rect 509968 379919 510088 380285
rect 509968 379885 510011 379919
rect 510045 379885 510088 379919
rect 509968 379519 510088 379885
rect 509968 379485 510011 379519
rect 510045 379485 510088 379519
rect 509968 379119 510088 379485
rect 509968 379085 510011 379119
rect 510045 379085 510088 379119
rect 509968 378719 510088 379085
rect 509968 378685 510011 378719
rect 510045 378685 510088 378719
rect 509968 378319 510088 378685
rect 509968 378285 510011 378319
rect 510045 378285 510088 378319
rect 509968 377919 510088 378285
rect 509968 377885 510011 377919
rect 510045 377885 510088 377919
rect 509968 377519 510088 377885
rect 509968 377485 510011 377519
rect 510045 377485 510088 377519
rect 509968 377119 510088 377485
rect 509968 377085 510011 377119
rect 510045 377085 510088 377119
rect 509968 376719 510088 377085
rect 509968 376685 510011 376719
rect 510045 376685 510088 376719
rect 509968 376319 510088 376685
rect 509968 376285 510011 376319
rect 510045 376285 510088 376319
rect 509968 375919 510088 376285
rect 509968 375885 510011 375919
rect 510045 375885 510088 375919
rect 509968 375519 510088 375885
rect 509968 375485 510011 375519
rect 510045 375485 510088 375519
rect 509968 375119 510088 375485
rect 509968 375085 510011 375119
rect 510045 375085 510088 375119
rect 509968 374719 510088 375085
rect 509968 374685 510011 374719
rect 510045 374685 510088 374719
rect 509968 374319 510088 374685
rect 509968 374285 510011 374319
rect 510045 374285 510088 374319
rect 508088 372953 508131 372987
rect 508165 372953 508208 372987
rect 508088 372787 508208 372953
rect 508088 372753 508131 372787
rect 508165 372753 508208 372787
rect 508088 372587 508208 372753
rect 508088 372553 508131 372587
rect 508165 372553 508208 372587
rect 508088 372387 508208 372553
rect 508088 372353 508131 372387
rect 508165 372353 508208 372387
rect 508088 372187 508208 372353
rect 508088 372153 508131 372187
rect 508165 372153 508208 372187
rect 508088 371987 508208 372153
rect 508088 371953 508131 371987
rect 508165 371953 508208 371987
rect 508088 371787 508208 371953
rect 508088 371753 508131 371787
rect 508165 371753 508208 371787
rect 508088 371587 508208 371753
rect 508088 371553 508131 371587
rect 508165 371553 508208 371587
rect 508088 371387 508208 371553
rect 508088 371353 508131 371387
rect 508165 371353 508208 371387
rect 508088 371187 508208 371353
rect 508088 371153 508131 371187
rect 508165 371153 508208 371187
rect 508088 370987 508208 371153
rect 508088 370953 508131 370987
rect 508165 370953 508208 370987
rect 508088 370787 508208 370953
rect 508088 370753 508131 370787
rect 508165 370753 508208 370787
rect 508088 370587 508208 370753
rect 508088 370553 508131 370587
rect 508165 370553 508208 370587
rect 508088 370387 508208 370553
rect 508088 370353 508131 370387
rect 508165 370353 508208 370387
rect 508088 370187 508208 370353
rect 508088 370153 508131 370187
rect 508165 370153 508208 370187
rect 508088 369987 508208 370153
rect 508088 369953 508131 369987
rect 508165 369953 508208 369987
rect 508088 369787 508208 369953
rect 508088 369753 508131 369787
rect 508165 369753 508208 369787
rect 508088 369587 508208 369753
rect 508088 369553 508131 369587
rect 508165 369553 508208 369587
rect 508088 369387 508208 369553
rect 508088 369353 508131 369387
rect 508165 369353 508208 369387
rect 508088 369187 508208 369353
rect 508088 369153 508131 369187
rect 508165 369153 508208 369187
rect 508088 368987 508208 369153
rect 508088 368953 508131 368987
rect 508165 368953 508208 368987
rect 508088 368787 508208 368953
rect 508088 368753 508131 368787
rect 508165 368753 508208 368787
rect 508088 368587 508208 368753
rect 508088 368553 508131 368587
rect 508165 368553 508208 368587
rect 508088 368387 508208 368553
rect 508088 368353 508131 368387
rect 508165 368353 508208 368387
rect 508088 368187 508208 368353
rect 508088 368153 508131 368187
rect 508165 368153 508208 368187
rect 508088 367987 508208 368153
rect 508088 367953 508131 367987
rect 508165 367953 508208 367987
rect 508088 367787 508208 367953
rect 508088 367753 508131 367787
rect 508165 367753 508208 367787
rect 508088 367587 508208 367753
rect 508088 367553 508131 367587
rect 508165 367553 508208 367587
rect 508088 367387 508208 367553
rect 508088 367353 508131 367387
rect 508165 367353 508208 367387
rect 508088 367187 508208 367353
rect 508088 367153 508131 367187
rect 508165 367153 508208 367187
rect 508088 366987 508208 367153
rect 508088 366953 508131 366987
rect 508165 366953 508208 366987
rect 508088 366787 508208 366953
rect 508088 366753 508131 366787
rect 508165 366753 508208 366787
rect 508088 366587 508208 366753
rect 508088 366553 508131 366587
rect 508165 366553 508208 366587
rect 508088 366387 508208 366553
rect 508088 366353 508131 366387
rect 508165 366353 508208 366387
rect 508088 366187 508208 366353
rect 508458 373124 508528 373144
rect 508458 373090 508464 373124
rect 508498 373090 508528 373124
rect 508458 373074 508528 373090
rect 508458 373034 508476 373074
rect 508458 373000 508464 373034
rect 508498 373000 508528 373022
rect 508458 372944 508528 373000
rect 509968 372987 510088 374285
rect 508458 372910 508464 372944
rect 508498 372910 508528 372944
rect 508458 372854 508528 372910
rect 508458 372820 508464 372854
rect 508498 372820 508528 372854
rect 508458 372764 508528 372820
rect 508458 372730 508464 372764
rect 508498 372730 508528 372764
rect 508458 372674 508528 372730
rect 508458 372640 508464 372674
rect 508498 372640 508528 372674
rect 508458 372584 508528 372640
rect 508458 372550 508464 372584
rect 508498 372550 508528 372584
rect 508458 372494 508528 372550
rect 508458 372460 508464 372494
rect 508498 372460 508528 372494
rect 508458 372404 508528 372460
rect 508458 372370 508464 372404
rect 508498 372370 508528 372404
rect 508458 372314 508528 372370
rect 508458 372280 508464 372314
rect 508498 372280 508528 372314
rect 508458 372234 508528 372280
rect 508608 372960 508678 372980
rect 508608 372926 508624 372960
rect 508658 372926 508678 372960
rect 508608 372870 508678 372926
rect 508608 372836 508624 372870
rect 508658 372836 508678 372870
rect 508608 372780 508678 372836
rect 509968 372953 510011 372987
rect 510045 372953 510088 372987
rect 508608 372746 508624 372780
rect 508658 372746 508678 372780
rect 508608 372690 508678 372746
rect 508608 372656 508624 372690
rect 508658 372656 508678 372690
rect 508608 372600 508678 372656
rect 508608 372566 508624 372600
rect 508658 372566 508678 372600
rect 508608 372510 508678 372566
rect 508608 372476 508624 372510
rect 508658 372476 508678 372510
rect 508608 372420 508678 372476
rect 508608 372386 508624 372420
rect 508658 372386 508678 372420
rect 508608 372330 508678 372386
rect 508608 372296 508624 372330
rect 508658 372296 508678 372330
rect 508608 372240 508678 372296
rect 508608 372234 508624 372240
rect 508458 372224 508624 372234
rect 508458 372190 508464 372224
rect 508498 372206 508624 372224
rect 508658 372206 508678 372240
rect 508498 372190 508528 372206
rect 508458 372134 508528 372190
rect 508458 372100 508464 372134
rect 508498 372100 508528 372134
rect 508458 372044 508528 372100
rect 508458 372010 508464 372044
rect 508498 372010 508528 372044
rect 508458 371954 508528 372010
rect 508458 371920 508464 371954
rect 508498 371920 508528 371954
rect 508458 371784 508528 371920
rect 508458 371750 508464 371784
rect 508498 371750 508528 371784
rect 508458 371694 508528 371750
rect 508458 371660 508464 371694
rect 508498 371660 508528 371694
rect 508458 371604 508528 371660
rect 508458 371570 508464 371604
rect 508498 371570 508528 371604
rect 508458 371514 508528 371570
rect 508458 371480 508464 371514
rect 508498 371480 508528 371514
rect 508458 371424 508528 371480
rect 508458 371390 508464 371424
rect 508498 371390 508528 371424
rect 508458 371334 508528 371390
rect 508458 371300 508464 371334
rect 508498 371300 508528 371334
rect 508458 371244 508528 371300
rect 508458 371210 508464 371244
rect 508498 371210 508528 371244
rect 508458 371154 508528 371210
rect 508458 371120 508464 371154
rect 508498 371120 508528 371154
rect 508458 371064 508528 371120
rect 508458 371030 508464 371064
rect 508498 371030 508528 371064
rect 508458 370974 508528 371030
rect 508458 370940 508464 370974
rect 508498 370940 508528 370974
rect 508458 370884 508528 370940
rect 508458 370850 508464 370884
rect 508498 370850 508528 370884
rect 508458 370794 508528 370850
rect 508458 370760 508464 370794
rect 508498 370760 508528 370794
rect 508458 370704 508528 370760
rect 508458 370670 508464 370704
rect 508498 370670 508528 370704
rect 508458 370614 508528 370670
rect 508458 370580 508464 370614
rect 508498 370580 508528 370614
rect 508458 370444 508528 370580
rect 508458 370410 508464 370444
rect 508498 370410 508528 370444
rect 508458 370354 508528 370410
rect 508458 370320 508464 370354
rect 508498 370320 508528 370354
rect 508458 370264 508528 370320
rect 508458 370230 508464 370264
rect 508498 370230 508528 370264
rect 508458 370174 508528 370230
rect 508458 370140 508464 370174
rect 508498 370140 508528 370174
rect 508458 370084 508528 370140
rect 508458 370050 508464 370084
rect 508498 370050 508528 370084
rect 508458 369994 508528 370050
rect 508458 369960 508464 369994
rect 508498 369960 508528 369994
rect 508458 369904 508528 369960
rect 508458 369870 508464 369904
rect 508498 369870 508528 369904
rect 508458 369814 508528 369870
rect 508458 369780 508464 369814
rect 508498 369780 508528 369814
rect 508458 369724 508528 369780
rect 508458 369690 508464 369724
rect 508498 369690 508528 369724
rect 508458 369634 508528 369690
rect 508458 369600 508464 369634
rect 508498 369600 508528 369634
rect 508458 369544 508528 369600
rect 508458 369510 508464 369544
rect 508498 369510 508528 369544
rect 508458 369454 508528 369510
rect 508458 369420 508464 369454
rect 508498 369420 508528 369454
rect 508458 369364 508528 369420
rect 508458 369330 508464 369364
rect 508498 369330 508528 369364
rect 508458 369274 508528 369330
rect 508458 369240 508464 369274
rect 508498 369240 508528 369274
rect 508458 369104 508528 369240
rect 508458 369070 508464 369104
rect 508498 369070 508528 369104
rect 508458 369014 508528 369070
rect 508458 368980 508464 369014
rect 508498 368980 508528 369014
rect 508458 368924 508528 368980
rect 508458 368890 508464 368924
rect 508498 368890 508528 368924
rect 508458 368834 508528 368890
rect 508458 368800 508464 368834
rect 508498 368800 508528 368834
rect 508458 368744 508528 368800
rect 508458 368710 508464 368744
rect 508498 368710 508528 368744
rect 508458 368654 508528 368710
rect 508458 368620 508464 368654
rect 508498 368620 508528 368654
rect 508458 368564 508528 368620
rect 508458 368530 508464 368564
rect 508498 368530 508528 368564
rect 508458 368474 508528 368530
rect 508458 368440 508464 368474
rect 508498 368440 508528 368474
rect 508458 368384 508528 368440
rect 508458 368350 508464 368384
rect 508498 368350 508528 368384
rect 508458 368294 508528 368350
rect 508458 368260 508464 368294
rect 508498 368260 508528 368294
rect 508458 368204 508528 368260
rect 508458 368170 508464 368204
rect 508498 368170 508528 368204
rect 508458 368114 508528 368170
rect 508458 368080 508464 368114
rect 508498 368080 508528 368114
rect 508458 368024 508528 368080
rect 508458 367990 508464 368024
rect 508498 367990 508528 368024
rect 508458 367934 508528 367990
rect 508458 367900 508464 367934
rect 508498 367900 508528 367934
rect 508458 367764 508528 367900
rect 508458 367730 508464 367764
rect 508498 367730 508528 367764
rect 508458 367674 508528 367730
rect 508458 367640 508464 367674
rect 508498 367640 508528 367674
rect 508458 367584 508528 367640
rect 508458 367550 508464 367584
rect 508498 367550 508528 367584
rect 508458 367494 508528 367550
rect 508458 367460 508464 367494
rect 508498 367460 508528 367494
rect 508458 367404 508528 367460
rect 508458 367370 508464 367404
rect 508498 367370 508528 367404
rect 508458 367314 508528 367370
rect 508458 367280 508464 367314
rect 508498 367280 508528 367314
rect 508458 367224 508528 367280
rect 508458 367190 508464 367224
rect 508498 367190 508528 367224
rect 508458 367134 508528 367190
rect 508458 367100 508464 367134
rect 508498 367100 508528 367134
rect 508458 367044 508528 367100
rect 508458 367010 508464 367044
rect 508498 367010 508528 367044
rect 508458 366954 508528 367010
rect 508458 366920 508464 366954
rect 508498 366920 508528 366954
rect 508458 366864 508528 366920
rect 508458 366830 508464 366864
rect 508498 366830 508528 366864
rect 508458 366774 508528 366830
rect 508458 366740 508464 366774
rect 508498 366740 508528 366774
rect 508458 366684 508528 366740
rect 508458 366650 508464 366684
rect 508498 366650 508528 366684
rect 508458 366594 508528 366650
rect 508458 366560 508464 366594
rect 508498 366560 508528 366594
rect 508458 366424 508528 366560
rect 508458 366390 508464 366424
rect 508498 366390 508528 366424
rect 508458 366334 508528 366390
rect 508458 366300 508464 366334
rect 508498 366300 508528 366334
rect 508272 366266 508324 366272
rect 508324 366226 508380 366254
rect 508272 366208 508324 366214
rect 508088 366153 508131 366187
rect 508165 366153 508208 366187
rect 508088 365987 508208 366153
rect 508088 365953 508131 365987
rect 508165 365953 508208 365987
rect 508088 365787 508208 365953
rect 508088 365753 508131 365787
rect 508165 365753 508208 365787
rect 508088 365587 508208 365753
rect 508088 365553 508131 365587
rect 508165 365553 508208 365587
rect 508088 365387 508208 365553
rect 508088 365353 508131 365387
rect 508165 365353 508208 365387
rect 508088 365187 508208 365353
rect 508088 365153 508131 365187
rect 508165 365153 508208 365187
rect 508088 364987 508208 365153
rect 508088 364953 508131 364987
rect 508165 364953 508208 364987
rect 508088 364787 508208 364953
rect 508088 364753 508131 364787
rect 508165 364753 508208 364787
rect 508088 364587 508208 364753
rect 508088 364553 508131 364587
rect 508165 364553 508208 364587
rect 508088 364387 508208 364553
rect 508088 364353 508131 364387
rect 508165 364353 508208 364387
rect 508088 364187 508208 364353
rect 508088 364153 508131 364187
rect 508165 364153 508208 364187
rect 508088 363987 508208 364153
rect 508088 363953 508131 363987
rect 508165 363953 508208 363987
rect 508088 363787 508208 363953
rect 508088 363753 508131 363787
rect 508165 363753 508208 363787
rect 508088 363587 508208 363753
rect 508088 363553 508131 363587
rect 508165 363553 508208 363587
rect 508088 363387 508208 363553
rect 508088 363353 508131 363387
rect 508165 363353 508208 363387
rect 508088 363187 508208 363353
rect 508088 363153 508131 363187
rect 508165 363153 508208 363187
rect 508088 362987 508208 363153
rect 508088 362953 508131 362987
rect 508165 362953 508208 362987
rect 508088 362787 508208 362953
rect 508088 362753 508131 362787
rect 508165 362753 508208 362787
rect 508088 362587 508208 362753
rect 508088 362553 508131 362587
rect 508165 362553 508208 362587
rect 508088 361476 508208 362553
rect 508088 359888 508090 361476
rect 508206 359888 508208 361476
rect 508088 359866 508208 359888
rect 506208 357440 506210 359028
rect 506326 357440 506328 359028
rect 506208 357418 506328 357440
rect 508352 356582 508380 366226
rect 508458 366244 508528 366300
rect 508458 366210 508464 366244
rect 508498 366210 508528 366244
rect 508458 366154 508528 366210
rect 508458 366120 508464 366154
rect 508498 366120 508528 366154
rect 508458 366064 508528 366120
rect 508458 366030 508464 366064
rect 508498 366030 508528 366064
rect 508458 365974 508528 366030
rect 508458 365940 508464 365974
rect 508498 365940 508528 365974
rect 508458 365884 508528 365940
rect 508458 365850 508464 365884
rect 508498 365850 508528 365884
rect 508458 365794 508528 365850
rect 508458 365760 508464 365794
rect 508498 365760 508528 365794
rect 508458 365704 508528 365760
rect 508458 365670 508464 365704
rect 508498 365670 508528 365704
rect 508458 365614 508528 365670
rect 508458 365580 508464 365614
rect 508498 365580 508528 365614
rect 508458 365524 508528 365580
rect 508458 365490 508464 365524
rect 508498 365490 508528 365524
rect 508458 365434 508528 365490
rect 508458 365400 508464 365434
rect 508498 365400 508528 365434
rect 508458 365344 508528 365400
rect 508458 365310 508464 365344
rect 508498 365310 508528 365344
rect 508458 365254 508528 365310
rect 508458 365220 508464 365254
rect 508498 365220 508528 365254
rect 508458 365084 508528 365220
rect 508458 365050 508464 365084
rect 508498 365050 508528 365084
rect 508458 364994 508528 365050
rect 508458 364960 508464 364994
rect 508498 364960 508528 364994
rect 508458 364904 508528 364960
rect 508458 364870 508464 364904
rect 508498 364870 508528 364904
rect 508458 364814 508528 364870
rect 508458 364780 508464 364814
rect 508498 364780 508528 364814
rect 508458 364724 508528 364780
rect 508458 364690 508464 364724
rect 508498 364690 508528 364724
rect 508458 364634 508528 364690
rect 508458 364600 508464 364634
rect 508498 364600 508528 364634
rect 508458 364544 508528 364600
rect 508458 364510 508464 364544
rect 508498 364510 508528 364544
rect 508458 364454 508528 364510
rect 508458 364420 508464 364454
rect 508498 364420 508528 364454
rect 508458 364364 508528 364420
rect 508458 364330 508464 364364
rect 508498 364330 508528 364364
rect 508458 364274 508528 364330
rect 508458 364240 508464 364274
rect 508498 364240 508528 364274
rect 508458 364184 508528 364240
rect 508458 364150 508464 364184
rect 508498 364150 508528 364184
rect 508458 364094 508528 364150
rect 508458 364060 508464 364094
rect 508498 364060 508528 364094
rect 508458 364004 508528 364060
rect 508458 363970 508464 364004
rect 508498 363970 508528 364004
rect 508458 363914 508528 363970
rect 508458 363880 508464 363914
rect 508498 363880 508528 363914
rect 508458 363744 508528 363880
rect 508458 363710 508464 363744
rect 508498 363710 508528 363744
rect 508458 363654 508528 363710
rect 508458 363620 508464 363654
rect 508498 363620 508528 363654
rect 508458 363564 508528 363620
rect 508458 363530 508464 363564
rect 508498 363530 508528 363564
rect 508458 363474 508528 363530
rect 508458 363440 508464 363474
rect 508498 363440 508528 363474
rect 508458 363384 508528 363440
rect 508458 363350 508464 363384
rect 508498 363350 508528 363384
rect 508458 363294 508528 363350
rect 508458 363260 508464 363294
rect 508498 363260 508528 363294
rect 508458 363204 508528 363260
rect 508458 363170 508464 363204
rect 508498 363170 508528 363204
rect 508458 363114 508528 363170
rect 508458 363080 508464 363114
rect 508498 363080 508528 363114
rect 508458 363024 508528 363080
rect 508458 362990 508464 363024
rect 508498 362990 508528 363024
rect 508458 362934 508528 362990
rect 508458 362900 508464 362934
rect 508498 362900 508528 362934
rect 508458 362844 508528 362900
rect 508458 362810 508464 362844
rect 508498 362810 508528 362844
rect 508458 362754 508528 362810
rect 508458 362720 508464 362754
rect 508498 362720 508528 362754
rect 508458 362664 508528 362720
rect 508458 362630 508464 362664
rect 508498 362630 508528 362664
rect 508608 372150 508678 372206
rect 508608 372116 508624 372150
rect 508658 372116 508678 372150
rect 508608 372060 508678 372116
rect 508608 372026 508624 372060
rect 508658 372026 508678 372060
rect 508608 371620 508678 372026
rect 508608 371586 508624 371620
rect 508658 371586 508678 371620
rect 508608 371530 508678 371586
rect 508608 371496 508624 371530
rect 508658 371496 508678 371530
rect 508608 371440 508678 371496
rect 508608 371406 508624 371440
rect 508658 371406 508678 371440
rect 508608 371350 508678 371406
rect 508608 371316 508624 371350
rect 508658 371316 508678 371350
rect 508608 371260 508678 371316
rect 508608 371226 508624 371260
rect 508658 371226 508678 371260
rect 508608 371170 508678 371226
rect 508608 371136 508624 371170
rect 508658 371136 508678 371170
rect 508608 371080 508678 371136
rect 508608 371046 508624 371080
rect 508658 371046 508678 371080
rect 508608 370990 508678 371046
rect 508608 370956 508624 370990
rect 508658 370956 508678 370990
rect 508608 370900 508678 370956
rect 508608 370866 508624 370900
rect 508658 370866 508678 370900
rect 508608 370810 508678 370866
rect 508608 370776 508624 370810
rect 508658 370776 508678 370810
rect 508608 370720 508678 370776
rect 508608 370686 508624 370720
rect 508658 370686 508678 370720
rect 508608 370280 508678 370686
rect 508608 370246 508624 370280
rect 508658 370246 508678 370280
rect 508608 370190 508678 370246
rect 508608 370156 508624 370190
rect 508658 370156 508678 370190
rect 508608 370100 508678 370156
rect 508608 370066 508624 370100
rect 508658 370066 508678 370100
rect 508608 370010 508678 370066
rect 508608 369976 508624 370010
rect 508658 369976 508678 370010
rect 508608 369920 508678 369976
rect 508608 369886 508624 369920
rect 508658 369886 508678 369920
rect 508608 369830 508678 369886
rect 508608 369796 508624 369830
rect 508658 369796 508678 369830
rect 508608 369740 508678 369796
rect 508608 369706 508624 369740
rect 508658 369706 508678 369740
rect 508608 369650 508678 369706
rect 508608 369616 508624 369650
rect 508658 369616 508678 369650
rect 508608 369560 508678 369616
rect 508608 369526 508624 369560
rect 508658 369526 508678 369560
rect 508608 369470 508678 369526
rect 508608 369436 508624 369470
rect 508658 369436 508678 369470
rect 508608 369380 508678 369436
rect 508608 369346 508624 369380
rect 508658 369346 508678 369380
rect 508608 368940 508678 369346
rect 508608 368906 508624 368940
rect 508658 368906 508678 368940
rect 508608 368850 508678 368906
rect 508608 368816 508624 368850
rect 508658 368816 508678 368850
rect 508608 368760 508678 368816
rect 508608 368726 508624 368760
rect 508658 368726 508678 368760
rect 508608 368670 508678 368726
rect 508608 368636 508624 368670
rect 508658 368636 508678 368670
rect 508608 368580 508678 368636
rect 508608 368546 508624 368580
rect 508658 368546 508678 368580
rect 508608 368490 508678 368546
rect 508608 368456 508624 368490
rect 508658 368456 508678 368490
rect 508608 368400 508678 368456
rect 508608 368366 508624 368400
rect 508658 368366 508678 368400
rect 508608 368310 508678 368366
rect 508608 368276 508624 368310
rect 508658 368276 508678 368310
rect 508608 368220 508678 368276
rect 508608 368186 508624 368220
rect 508658 368186 508678 368220
rect 508608 368130 508678 368186
rect 508608 368096 508624 368130
rect 508658 368096 508678 368130
rect 508608 368040 508678 368096
rect 508608 368006 508624 368040
rect 508658 368006 508678 368040
rect 508608 367600 508678 368006
rect 508608 367566 508624 367600
rect 508658 367566 508678 367600
rect 508608 367510 508678 367566
rect 508608 367476 508624 367510
rect 508658 367476 508678 367510
rect 508608 367420 508678 367476
rect 508608 367386 508624 367420
rect 508658 367386 508678 367420
rect 508608 367330 508678 367386
rect 508608 367296 508624 367330
rect 508658 367296 508678 367330
rect 508608 367240 508678 367296
rect 508608 367206 508624 367240
rect 508658 367206 508678 367240
rect 508608 367150 508678 367206
rect 508608 367116 508624 367150
rect 508658 367116 508678 367150
rect 508608 367060 508678 367116
rect 508608 367026 508624 367060
rect 508658 367026 508678 367060
rect 508608 366970 508678 367026
rect 508608 366936 508624 366970
rect 508658 366936 508678 366970
rect 508608 366880 508678 366936
rect 508608 366846 508624 366880
rect 508658 366846 508678 366880
rect 508608 366790 508678 366846
rect 508608 366756 508624 366790
rect 508658 366756 508678 366790
rect 508608 366700 508678 366756
rect 508608 366666 508624 366700
rect 508658 366666 508678 366700
rect 508608 366260 508678 366666
rect 508608 366226 508624 366260
rect 508658 366226 508678 366260
rect 508608 366170 508678 366226
rect 508608 366136 508624 366170
rect 508658 366136 508678 366170
rect 508608 366080 508678 366136
rect 508608 366046 508624 366080
rect 508658 366046 508678 366080
rect 508608 365990 508678 366046
rect 508608 365956 508624 365990
rect 508658 365956 508678 365990
rect 508608 365900 508678 365956
rect 508608 365866 508624 365900
rect 508658 365866 508678 365900
rect 508608 365810 508678 365866
rect 508608 365776 508624 365810
rect 508658 365776 508678 365810
rect 508608 365720 508678 365776
rect 508608 365686 508624 365720
rect 508658 365686 508678 365720
rect 508608 365630 508678 365686
rect 508608 365596 508624 365630
rect 508658 365596 508678 365630
rect 508608 365540 508678 365596
rect 508608 365506 508624 365540
rect 508658 365506 508678 365540
rect 508608 365450 508678 365506
rect 508608 365416 508624 365450
rect 508658 365416 508678 365450
rect 508608 365360 508678 365416
rect 508608 365326 508624 365360
rect 508658 365326 508678 365360
rect 508608 364920 508678 365326
rect 508608 364886 508624 364920
rect 508658 364886 508678 364920
rect 508608 364830 508678 364886
rect 508608 364796 508624 364830
rect 508658 364796 508678 364830
rect 508608 364740 508678 364796
rect 508608 364706 508624 364740
rect 508658 364706 508678 364740
rect 508608 364650 508678 364706
rect 508608 364616 508624 364650
rect 508658 364616 508678 364650
rect 508608 364560 508678 364616
rect 508608 364526 508624 364560
rect 508658 364526 508678 364560
rect 508608 364470 508678 364526
rect 508608 364436 508624 364470
rect 508658 364436 508678 364470
rect 508608 364380 508678 364436
rect 508608 364346 508624 364380
rect 508658 364346 508678 364380
rect 508608 364290 508678 364346
rect 508608 364256 508624 364290
rect 508658 364256 508678 364290
rect 508608 364200 508678 364256
rect 508608 364166 508624 364200
rect 508658 364166 508678 364200
rect 508608 364110 508678 364166
rect 508608 364076 508624 364110
rect 508658 364076 508678 364110
rect 508608 364020 508678 364076
rect 508608 363986 508624 364020
rect 508658 363986 508678 364020
rect 508608 363580 508678 363986
rect 508608 363546 508624 363580
rect 508658 363546 508678 363580
rect 508608 363490 508678 363546
rect 508608 363456 508624 363490
rect 508658 363456 508678 363490
rect 508608 363400 508678 363456
rect 508608 363366 508624 363400
rect 508658 363366 508678 363400
rect 508608 363310 508678 363366
rect 508608 363276 508624 363310
rect 508658 363276 508678 363310
rect 508608 363220 508678 363276
rect 508608 363186 508624 363220
rect 508658 363186 508678 363220
rect 508608 363130 508678 363186
rect 508608 363096 508624 363130
rect 508658 363096 508678 363130
rect 508608 363040 508678 363096
rect 508608 363006 508624 363040
rect 508658 363006 508678 363040
rect 508608 362950 508678 363006
rect 508608 362916 508624 362950
rect 508658 362916 508678 362950
rect 508608 362860 508678 362916
rect 508608 362826 508624 362860
rect 508658 362826 508678 362860
rect 508608 362770 508678 362826
rect 508782 372798 509394 372806
rect 508782 372746 508816 372798
rect 508868 372774 509394 372798
rect 508868 372746 508928 372774
rect 508782 372740 508828 372746
rect 508862 372740 508928 372746
rect 508962 372740 509028 372774
rect 509062 372740 509128 372774
rect 509162 372740 509228 372774
rect 509262 372740 509328 372774
rect 509362 372740 509394 372774
rect 508782 372712 509394 372740
rect 509968 372787 510088 372953
rect 509968 372753 510011 372787
rect 510045 372753 510088 372787
rect 508782 372706 509412 372712
rect 508782 372674 509360 372706
rect 508782 372640 508828 372674
rect 508862 372640 508928 372674
rect 508962 372640 509028 372674
rect 509062 372640 509128 372674
rect 509162 372640 509228 372674
rect 509262 372640 509328 372674
rect 509362 372648 509412 372654
rect 509362 372640 509394 372648
rect 508782 372574 509394 372640
rect 508782 372540 508828 372574
rect 508862 372540 508928 372574
rect 508962 372540 509028 372574
rect 509062 372540 509128 372574
rect 509162 372540 509228 372574
rect 509262 372540 509328 372574
rect 509362 372540 509394 372574
rect 508782 372474 509394 372540
rect 508782 372440 508828 372474
rect 508862 372440 508928 372474
rect 508962 372440 509028 372474
rect 509062 372440 509128 372474
rect 509162 372440 509228 372474
rect 509262 372440 509328 372474
rect 509362 372440 509394 372474
rect 508782 372374 509394 372440
rect 508782 372340 508828 372374
rect 508862 372340 508928 372374
rect 508962 372340 509028 372374
rect 509062 372340 509128 372374
rect 509162 372340 509228 372374
rect 509262 372340 509328 372374
rect 509362 372340 509394 372374
rect 508782 372274 509394 372340
rect 508782 372240 508828 372274
rect 508862 372240 508928 372274
rect 508962 372240 509028 372274
rect 509062 372240 509128 372274
rect 509162 372240 509228 372274
rect 509262 372240 509328 372274
rect 509362 372240 509394 372274
rect 508782 371434 509394 372240
rect 508782 371400 508828 371434
rect 508862 371400 508928 371434
rect 508962 371400 509028 371434
rect 509062 371400 509128 371434
rect 509162 371400 509228 371434
rect 509262 371400 509328 371434
rect 509362 371400 509394 371434
rect 508782 371334 509394 371400
rect 508782 371300 508828 371334
rect 508862 371300 508928 371334
rect 508962 371300 509028 371334
rect 509062 371300 509128 371334
rect 509162 371300 509228 371334
rect 509262 371300 509328 371334
rect 509362 371300 509394 371334
rect 508782 371234 509394 371300
rect 508782 371200 508828 371234
rect 508862 371200 508928 371234
rect 508962 371200 509028 371234
rect 509062 371200 509128 371234
rect 509162 371200 509228 371234
rect 509262 371200 509328 371234
rect 509362 371200 509394 371234
rect 508782 371134 509394 371200
rect 508782 371100 508828 371134
rect 508862 371100 508928 371134
rect 508962 371100 509028 371134
rect 509062 371100 509128 371134
rect 509162 371100 509228 371134
rect 509262 371100 509328 371134
rect 509362 371100 509394 371134
rect 508782 371034 509394 371100
rect 508782 371000 508828 371034
rect 508862 371000 508928 371034
rect 508962 371000 509028 371034
rect 509062 371000 509128 371034
rect 509162 371000 509228 371034
rect 509262 371000 509328 371034
rect 509362 371000 509394 371034
rect 508782 370934 509394 371000
rect 508782 370900 508828 370934
rect 508862 370900 508928 370934
rect 508962 370900 509028 370934
rect 509062 370900 509128 370934
rect 509162 370900 509228 370934
rect 509262 370900 509328 370934
rect 509362 370900 509394 370934
rect 508782 370094 509394 370900
rect 508782 370060 508828 370094
rect 508862 370060 508928 370094
rect 508962 370060 509028 370094
rect 509062 370060 509128 370094
rect 509162 370060 509228 370094
rect 509262 370060 509328 370094
rect 509362 370060 509394 370094
rect 508782 369994 509394 370060
rect 508782 369960 508828 369994
rect 508862 369960 508928 369994
rect 508962 369960 509028 369994
rect 509062 369960 509128 369994
rect 509162 369960 509228 369994
rect 509262 369960 509328 369994
rect 509362 369960 509394 369994
rect 508782 369894 509394 369960
rect 508782 369860 508828 369894
rect 508862 369860 508928 369894
rect 508962 369860 509028 369894
rect 509062 369860 509128 369894
rect 509162 369860 509228 369894
rect 509262 369860 509328 369894
rect 509362 369860 509394 369894
rect 508782 369794 509394 369860
rect 508782 369760 508828 369794
rect 508862 369760 508928 369794
rect 508962 369760 509028 369794
rect 509062 369760 509128 369794
rect 509162 369760 509228 369794
rect 509262 369760 509328 369794
rect 509362 369760 509394 369794
rect 508782 369694 509394 369760
rect 508782 369660 508828 369694
rect 508862 369660 508928 369694
rect 508962 369660 509028 369694
rect 509062 369660 509128 369694
rect 509162 369660 509228 369694
rect 509262 369660 509328 369694
rect 509362 369660 509394 369694
rect 508782 369594 509394 369660
rect 508782 369560 508828 369594
rect 508862 369560 508928 369594
rect 508962 369560 509028 369594
rect 509062 369560 509128 369594
rect 509162 369560 509228 369594
rect 509262 369560 509328 369594
rect 509362 369560 509394 369594
rect 508782 368754 509394 369560
rect 508782 368720 508828 368754
rect 508862 368720 508928 368754
rect 508962 368720 509028 368754
rect 509062 368720 509128 368754
rect 509162 368720 509228 368754
rect 509262 368720 509328 368754
rect 509362 368720 509394 368754
rect 508782 368654 509394 368720
rect 508782 368620 508828 368654
rect 508862 368620 508928 368654
rect 508962 368620 509028 368654
rect 509062 368620 509128 368654
rect 509162 368620 509228 368654
rect 509262 368620 509328 368654
rect 509362 368620 509394 368654
rect 508782 368554 509394 368620
rect 508782 368520 508828 368554
rect 508862 368520 508928 368554
rect 508962 368520 509028 368554
rect 509062 368520 509128 368554
rect 509162 368520 509228 368554
rect 509262 368520 509328 368554
rect 509362 368520 509394 368554
rect 508782 368454 509394 368520
rect 508782 368420 508828 368454
rect 508862 368420 508928 368454
rect 508962 368420 509028 368454
rect 509062 368420 509128 368454
rect 509162 368420 509228 368454
rect 509262 368420 509328 368454
rect 509362 368420 509394 368454
rect 508782 368354 509394 368420
rect 508782 368320 508828 368354
rect 508862 368320 508928 368354
rect 508962 368320 509028 368354
rect 509062 368320 509128 368354
rect 509162 368320 509228 368354
rect 509262 368320 509328 368354
rect 509362 368320 509394 368354
rect 508782 368254 509394 368320
rect 508782 368220 508828 368254
rect 508862 368220 508928 368254
rect 508962 368220 509028 368254
rect 509062 368220 509128 368254
rect 509162 368220 509228 368254
rect 509262 368220 509328 368254
rect 509362 368220 509394 368254
rect 508782 367414 509394 368220
rect 508782 367380 508828 367414
rect 508862 367380 508928 367414
rect 508962 367380 509028 367414
rect 509062 367380 509128 367414
rect 509162 367380 509228 367414
rect 509262 367380 509328 367414
rect 509362 367380 509394 367414
rect 508782 367314 509394 367380
rect 508782 367280 508828 367314
rect 508862 367280 508928 367314
rect 508962 367280 509028 367314
rect 509062 367280 509128 367314
rect 509162 367280 509228 367314
rect 509262 367280 509328 367314
rect 509362 367280 509394 367314
rect 508782 367214 509394 367280
rect 508782 367180 508828 367214
rect 508862 367180 508928 367214
rect 508962 367180 509028 367214
rect 509062 367180 509128 367214
rect 509162 367180 509228 367214
rect 509262 367180 509328 367214
rect 509362 367180 509394 367214
rect 508782 367114 509394 367180
rect 508782 367080 508828 367114
rect 508862 367080 508928 367114
rect 508962 367080 509028 367114
rect 509062 367080 509128 367114
rect 509162 367080 509228 367114
rect 509262 367080 509328 367114
rect 509362 367080 509394 367114
rect 508782 367014 509394 367080
rect 508782 366980 508828 367014
rect 508862 366980 508928 367014
rect 508962 366980 509028 367014
rect 509062 366980 509128 367014
rect 509162 366980 509228 367014
rect 509262 366980 509328 367014
rect 509362 366980 509394 367014
rect 508782 366914 509394 366980
rect 508782 366880 508828 366914
rect 508862 366880 508928 366914
rect 508962 366880 509028 366914
rect 509062 366880 509128 366914
rect 509162 366880 509228 366914
rect 509262 366880 509328 366914
rect 509362 366880 509394 366914
rect 508782 366074 509394 366880
rect 508782 366040 508828 366074
rect 508862 366040 508928 366074
rect 508962 366040 509028 366074
rect 509062 366040 509128 366074
rect 509162 366040 509228 366074
rect 509262 366040 509328 366074
rect 509362 366040 509394 366074
rect 508782 365974 509394 366040
rect 508782 365940 508828 365974
rect 508862 365940 508928 365974
rect 508962 365940 509028 365974
rect 509062 365940 509128 365974
rect 509162 365940 509228 365974
rect 509262 365940 509328 365974
rect 509362 365940 509394 365974
rect 508782 365874 509394 365940
rect 508782 365840 508828 365874
rect 508862 365840 508928 365874
rect 508962 365840 509028 365874
rect 509062 365840 509128 365874
rect 509162 365840 509228 365874
rect 509262 365840 509328 365874
rect 509362 365840 509394 365874
rect 508782 365774 509394 365840
rect 508782 365740 508828 365774
rect 508862 365740 508928 365774
rect 508962 365740 509028 365774
rect 509062 365740 509128 365774
rect 509162 365740 509228 365774
rect 509262 365740 509328 365774
rect 509362 365740 509394 365774
rect 508782 365674 509394 365740
rect 508782 365640 508828 365674
rect 508862 365640 508928 365674
rect 508962 365640 509028 365674
rect 509062 365640 509128 365674
rect 509162 365640 509228 365674
rect 509262 365640 509328 365674
rect 509362 365640 509394 365674
rect 508782 365574 509394 365640
rect 508782 365540 508828 365574
rect 508862 365540 508928 365574
rect 508962 365540 509028 365574
rect 509062 365540 509128 365574
rect 509162 365540 509228 365574
rect 509262 365540 509328 365574
rect 509362 365540 509394 365574
rect 508782 364734 509394 365540
rect 508782 364700 508828 364734
rect 508862 364700 508928 364734
rect 508962 364700 509028 364734
rect 509062 364700 509128 364734
rect 509162 364700 509228 364734
rect 509262 364700 509328 364734
rect 509362 364700 509394 364734
rect 508782 364634 509394 364700
rect 508782 364600 508828 364634
rect 508862 364600 508928 364634
rect 508962 364600 509028 364634
rect 509062 364600 509128 364634
rect 509162 364600 509228 364634
rect 509262 364600 509328 364634
rect 509362 364600 509394 364634
rect 508782 364534 509394 364600
rect 508782 364500 508828 364534
rect 508862 364500 508928 364534
rect 508962 364500 509028 364534
rect 509062 364500 509128 364534
rect 509162 364500 509228 364534
rect 509262 364500 509328 364534
rect 509362 364500 509394 364534
rect 508782 364434 509394 364500
rect 508782 364400 508828 364434
rect 508862 364400 508928 364434
rect 508962 364400 509028 364434
rect 509062 364400 509128 364434
rect 509162 364400 509228 364434
rect 509262 364400 509328 364434
rect 509362 364400 509394 364434
rect 508782 364334 509394 364400
rect 508782 364300 508828 364334
rect 508862 364300 508928 364334
rect 508962 364300 509028 364334
rect 509062 364300 509128 364334
rect 509162 364300 509228 364334
rect 509262 364300 509328 364334
rect 509362 364300 509394 364334
rect 508782 364234 509394 364300
rect 508782 364200 508828 364234
rect 508862 364200 508928 364234
rect 508962 364200 509028 364234
rect 509062 364200 509128 364234
rect 509162 364200 509228 364234
rect 509262 364200 509328 364234
rect 509362 364200 509394 364234
rect 508782 363394 509394 364200
rect 508782 363360 508828 363394
rect 508862 363360 508928 363394
rect 508962 363360 509028 363394
rect 509062 363360 509128 363394
rect 509162 363360 509228 363394
rect 509262 363360 509328 363394
rect 509362 363360 509394 363394
rect 508782 363294 509394 363360
rect 508782 363260 508828 363294
rect 508862 363260 508928 363294
rect 508962 363260 509028 363294
rect 509062 363260 509128 363294
rect 509162 363260 509228 363294
rect 509262 363260 509328 363294
rect 509362 363260 509394 363294
rect 508782 363194 509394 363260
rect 508782 363160 508828 363194
rect 508862 363160 508928 363194
rect 508962 363160 509028 363194
rect 509062 363160 509128 363194
rect 509162 363160 509228 363194
rect 509262 363160 509328 363194
rect 509362 363160 509394 363194
rect 508782 363094 509394 363160
rect 508782 363060 508828 363094
rect 508862 363060 508928 363094
rect 508962 363060 509028 363094
rect 509062 363060 509128 363094
rect 509162 363060 509228 363094
rect 509262 363060 509328 363094
rect 509362 363060 509394 363094
rect 508782 362994 509394 363060
rect 508782 362960 508828 362994
rect 508862 362960 508928 362994
rect 508962 362960 509028 362994
rect 509062 362960 509128 362994
rect 509162 362960 509228 362994
rect 509262 362960 509328 362994
rect 509362 362960 509394 362994
rect 508782 362894 509394 362960
rect 508782 362860 508828 362894
rect 508862 362860 508928 362894
rect 508962 362860 509028 362894
rect 509062 362860 509128 362894
rect 509162 362860 509228 362894
rect 509262 362860 509328 362894
rect 509362 362860 509394 362894
rect 508782 362814 509394 362860
rect 509968 372587 510088 372753
rect 509968 372553 510011 372587
rect 510045 372553 510088 372587
rect 509968 372387 510088 372553
rect 509968 372353 510011 372387
rect 510045 372353 510088 372387
rect 509968 372187 510088 372353
rect 509968 372153 510011 372187
rect 510045 372153 510088 372187
rect 509968 371987 510088 372153
rect 509968 371953 510011 371987
rect 510045 371953 510088 371987
rect 509968 371787 510088 371953
rect 509968 371753 510011 371787
rect 510045 371753 510088 371787
rect 509968 371587 510088 371753
rect 509968 371553 510011 371587
rect 510045 371553 510088 371587
rect 509968 371387 510088 371553
rect 509968 371353 510011 371387
rect 510045 371353 510088 371387
rect 509968 371187 510088 371353
rect 509968 371153 510011 371187
rect 510045 371153 510088 371187
rect 509968 370987 510088 371153
rect 509968 370953 510011 370987
rect 510045 370953 510088 370987
rect 509968 370787 510088 370953
rect 509968 370753 510011 370787
rect 510045 370753 510088 370787
rect 509968 370587 510088 370753
rect 509968 370553 510011 370587
rect 510045 370553 510088 370587
rect 509968 370387 510088 370553
rect 509968 370353 510011 370387
rect 510045 370353 510088 370387
rect 509968 370187 510088 370353
rect 509968 370153 510011 370187
rect 510045 370153 510088 370187
rect 509968 369987 510088 370153
rect 509968 369953 510011 369987
rect 510045 369953 510088 369987
rect 509968 369787 510088 369953
rect 509968 369753 510011 369787
rect 510045 369753 510088 369787
rect 509968 369587 510088 369753
rect 509968 369553 510011 369587
rect 510045 369553 510088 369587
rect 509968 369387 510088 369553
rect 509968 369353 510011 369387
rect 510045 369353 510088 369387
rect 509968 369187 510088 369353
rect 509968 369153 510011 369187
rect 510045 369153 510088 369187
rect 509968 368987 510088 369153
rect 509968 368953 510011 368987
rect 510045 368953 510088 368987
rect 509968 368787 510088 368953
rect 509968 368753 510011 368787
rect 510045 368753 510088 368787
rect 509968 368587 510088 368753
rect 509968 368553 510011 368587
rect 510045 368553 510088 368587
rect 509968 368387 510088 368553
rect 509968 368353 510011 368387
rect 510045 368353 510088 368387
rect 509968 368187 510088 368353
rect 509968 368153 510011 368187
rect 510045 368153 510088 368187
rect 509968 367987 510088 368153
rect 509968 367953 510011 367987
rect 510045 367953 510088 367987
rect 509968 367787 510088 367953
rect 509968 367753 510011 367787
rect 510045 367753 510088 367787
rect 509968 367587 510088 367753
rect 509968 367553 510011 367587
rect 510045 367553 510088 367587
rect 509968 367387 510088 367553
rect 509968 367353 510011 367387
rect 510045 367353 510088 367387
rect 509968 367187 510088 367353
rect 509968 367153 510011 367187
rect 510045 367153 510088 367187
rect 509968 366987 510088 367153
rect 509968 366953 510011 366987
rect 510045 366953 510088 366987
rect 509968 366787 510088 366953
rect 509968 366753 510011 366787
rect 510045 366753 510088 366787
rect 509968 366587 510088 366753
rect 509968 366553 510011 366587
rect 510045 366553 510088 366587
rect 509968 366387 510088 366553
rect 509968 366353 510011 366387
rect 510045 366353 510088 366387
rect 509968 366187 510088 366353
rect 509968 366153 510011 366187
rect 510045 366153 510088 366187
rect 509968 365987 510088 366153
rect 509968 365953 510011 365987
rect 510045 365953 510088 365987
rect 509968 365787 510088 365953
rect 509968 365753 510011 365787
rect 510045 365753 510088 365787
rect 509968 365587 510088 365753
rect 509968 365553 510011 365587
rect 510045 365553 510088 365587
rect 509968 365387 510088 365553
rect 509968 365353 510011 365387
rect 510045 365353 510088 365387
rect 509968 365187 510088 365353
rect 509968 365153 510011 365187
rect 510045 365153 510088 365187
rect 509968 364987 510088 365153
rect 509968 364953 510011 364987
rect 510045 364953 510088 364987
rect 509968 364787 510088 364953
rect 509968 364753 510011 364787
rect 510045 364753 510088 364787
rect 509968 364587 510088 364753
rect 509968 364553 510011 364587
rect 510045 364553 510088 364587
rect 509968 364387 510088 364553
rect 509968 364353 510011 364387
rect 510045 364353 510088 364387
rect 509968 364187 510088 364353
rect 509968 364153 510011 364187
rect 510045 364153 510088 364187
rect 509968 363987 510088 364153
rect 509968 363953 510011 363987
rect 510045 363953 510088 363987
rect 509968 363787 510088 363953
rect 509968 363753 510011 363787
rect 510045 363753 510088 363787
rect 509968 363587 510088 363753
rect 509968 363553 510011 363587
rect 510045 363553 510088 363587
rect 509968 363387 510088 363553
rect 509968 363353 510011 363387
rect 510045 363353 510088 363387
rect 509968 363187 510088 363353
rect 509968 363153 510011 363187
rect 510045 363153 510088 363187
rect 509968 362987 510088 363153
rect 509968 362953 510011 362987
rect 510045 362953 510088 362987
rect 508608 362736 508624 362770
rect 508658 362736 508678 362770
rect 508608 362680 508678 362736
rect 508608 362646 508624 362680
rect 508658 362646 508678 362680
rect 508608 362640 508678 362646
rect 509968 362787 510088 362953
rect 509968 362753 510011 362787
rect 510045 362753 510088 362787
rect 508458 362574 508528 362630
rect 508458 362540 508464 362574
rect 508498 362540 508528 362574
rect 508458 362476 508528 362540
rect 509968 362587 510088 362753
rect 509968 362553 510011 362587
rect 510045 362553 510088 362587
rect 509968 359028 510088 362553
rect 511848 411584 511968 411606
rect 511848 409996 511850 411584
rect 511966 409996 511968 411584
rect 511848 398251 511968 409996
rect 511848 398217 511891 398251
rect 511925 398217 511968 398251
rect 511848 398051 511968 398217
rect 511848 398017 511891 398051
rect 511925 398017 511968 398051
rect 511848 397851 511968 398017
rect 512147 398415 512709 398423
rect 512147 398021 512159 398415
rect 512697 398021 512709 398415
rect 512147 398013 512709 398021
rect 513107 398415 513669 398423
rect 513107 398021 513119 398415
rect 513657 398021 513669 398415
rect 513107 398013 513669 398021
rect 513728 398251 513848 412444
rect 517488 414032 517608 414054
rect 517488 412444 517490 414032
rect 517606 412444 517608 414032
rect 513728 398217 513771 398251
rect 513805 398217 513848 398251
rect 513728 398051 513848 398217
rect 513728 398017 513771 398051
rect 513805 398017 513848 398051
rect 511848 397817 511891 397851
rect 511925 397817 511968 397851
rect 511848 397651 511968 397817
rect 511848 397617 511891 397651
rect 511925 397617 511968 397651
rect 511848 397451 511968 397617
rect 511848 397417 511891 397451
rect 511925 397417 511968 397451
rect 511848 397251 511968 397417
rect 511848 397217 511891 397251
rect 511925 397217 511968 397251
rect 511848 397051 511968 397217
rect 511848 397017 511891 397051
rect 511925 397017 511968 397051
rect 511848 396851 511968 397017
rect 511848 396817 511891 396851
rect 511925 396817 511968 396851
rect 511848 396651 511968 396817
rect 511848 396617 511891 396651
rect 511925 396617 511968 396651
rect 511848 396451 511968 396617
rect 513112 396540 513140 398013
rect 513728 397851 513848 398017
rect 513728 397817 513771 397851
rect 513805 397817 513848 397851
rect 513728 397651 513848 397817
rect 513728 397617 513771 397651
rect 513805 397617 513848 397651
rect 513728 397451 513848 397617
rect 513728 397417 513771 397451
rect 513805 397417 513848 397451
rect 513728 397251 513848 397417
rect 513728 397217 513771 397251
rect 513805 397217 513848 397251
rect 513728 397051 513848 397217
rect 513728 397017 513771 397051
rect 513805 397017 513848 397051
rect 513728 396851 513848 397017
rect 513728 396817 513771 396851
rect 513805 396817 513848 396851
rect 513728 396651 513848 396817
rect 513728 396617 513771 396651
rect 513805 396617 513848 396651
rect 513100 396534 513152 396540
rect 513100 396476 513152 396482
rect 511848 396417 511891 396451
rect 511925 396417 511968 396451
rect 513728 396451 513848 396617
rect 511848 396251 511968 396417
rect 512709 396415 513673 396426
rect 511848 396217 511891 396251
rect 511925 396217 511968 396251
rect 511848 395507 511968 396217
rect 512147 396408 513673 396415
rect 512147 396014 512159 396408
rect 512697 396014 513119 396408
rect 513657 396014 513673 396408
rect 512147 396005 513673 396014
rect 512709 395994 513673 396005
rect 513728 396417 513771 396451
rect 513805 396417 513848 396451
rect 513728 396251 513848 396417
rect 513728 396217 513771 396251
rect 513805 396217 513848 396251
rect 512624 395890 512676 395896
rect 512624 395832 512676 395838
rect 512636 395679 512664 395832
rect 511848 395473 511891 395507
rect 511925 395473 511968 395507
rect 511848 395307 511968 395473
rect 511848 395273 511891 395307
rect 511925 395273 511968 395307
rect 511848 395107 511968 395273
rect 512147 395671 512709 395679
rect 512147 395277 512159 395671
rect 512697 395277 512709 395671
rect 512147 395269 512709 395277
rect 513107 395671 513669 395679
rect 513107 395277 513119 395671
rect 513657 395277 513669 395671
rect 513107 395269 513669 395277
rect 513728 395507 513848 396217
rect 513728 395473 513771 395507
rect 513805 395473 513848 395507
rect 513728 395307 513848 395473
rect 513728 395273 513771 395307
rect 513805 395273 513848 395307
rect 511848 395073 511891 395107
rect 511925 395073 511968 395107
rect 511848 394907 511968 395073
rect 511848 394873 511891 394907
rect 511925 394873 511968 394907
rect 511848 394707 511968 394873
rect 511848 394673 511891 394707
rect 511925 394673 511968 394707
rect 511848 394507 511968 394673
rect 511848 394473 511891 394507
rect 511925 394473 511968 394507
rect 511848 394307 511968 394473
rect 511848 394273 511891 394307
rect 511925 394273 511968 394307
rect 511848 394107 511968 394273
rect 511848 394073 511891 394107
rect 511925 394073 511968 394107
rect 511848 393907 511968 394073
rect 513112 394056 513140 395269
rect 513728 395107 513848 395273
rect 513728 395073 513771 395107
rect 513805 395073 513848 395107
rect 513728 394907 513848 395073
rect 513728 394873 513771 394907
rect 513805 394873 513848 394907
rect 513728 394707 513848 394873
rect 513728 394673 513771 394707
rect 513805 394673 513848 394707
rect 513728 394507 513848 394673
rect 513728 394473 513771 394507
rect 513805 394473 513848 394507
rect 513728 394307 513848 394473
rect 513728 394273 513771 394307
rect 513805 394273 513848 394307
rect 513728 394107 513848 394273
rect 513728 394073 513771 394107
rect 513805 394073 513848 394107
rect 512012 394050 512064 394056
rect 512012 393992 512064 393998
rect 513100 394050 513152 394056
rect 513100 393992 513152 393998
rect 511848 393873 511891 393907
rect 511925 393873 511968 393907
rect 511848 393707 511968 393873
rect 511848 393673 511891 393707
rect 511925 393673 511968 393707
rect 511848 393507 511968 393673
rect 511848 393473 511891 393507
rect 511925 393473 511968 393507
rect 511848 392763 511968 393473
rect 511848 392729 511891 392763
rect 511925 392729 511968 392763
rect 511848 392563 511968 392729
rect 512024 392584 512052 393992
rect 513728 393907 513848 394073
rect 513728 393873 513771 393907
rect 513805 393873 513848 393907
rect 513728 393707 513848 393873
rect 512709 393671 513673 393682
rect 512147 393664 513673 393671
rect 512147 393270 512159 393664
rect 512697 393270 513119 393664
rect 513657 393270 513673 393664
rect 512147 393261 513673 393270
rect 512709 393250 513673 393261
rect 513728 393673 513771 393707
rect 513805 393673 513848 393707
rect 513728 393507 513848 393673
rect 513728 393473 513771 393507
rect 513805 393473 513848 393507
rect 513094 393170 513100 393222
rect 513152 393170 513158 393222
rect 513112 392935 513140 393170
rect 512147 392927 512709 392935
rect 512147 392762 512159 392927
rect 512147 392710 512148 392762
rect 511848 392529 511891 392563
rect 511925 392529 511968 392563
rect 511848 392363 511968 392529
rect 512012 392578 512064 392584
rect 512012 392520 512064 392526
rect 512147 392533 512159 392710
rect 512697 392533 512709 392927
rect 512147 392525 512709 392533
rect 513107 392927 513669 392935
rect 513107 392533 513119 392927
rect 513657 392533 513669 392927
rect 513107 392525 513669 392533
rect 513728 392763 513848 393473
rect 513728 392729 513771 392763
rect 513805 392729 513848 392763
rect 513728 392563 513848 392729
rect 513728 392529 513771 392563
rect 513805 392529 513848 392563
rect 511848 392329 511891 392363
rect 511925 392329 511968 392363
rect 511848 392163 511968 392329
rect 511848 392129 511891 392163
rect 511925 392129 511968 392163
rect 511848 391963 511968 392129
rect 511848 391929 511891 391963
rect 511925 391929 511968 391963
rect 511848 391763 511968 391929
rect 511848 391729 511891 391763
rect 511925 391729 511968 391763
rect 511848 391563 511968 391729
rect 511848 391529 511891 391563
rect 511925 391529 511968 391563
rect 511848 391363 511968 391529
rect 511848 391329 511891 391363
rect 511925 391329 511968 391363
rect 511848 391163 511968 391329
rect 511848 391129 511891 391163
rect 511925 391129 511968 391163
rect 511848 390963 511968 391129
rect 511848 390929 511891 390963
rect 511925 390929 511968 390963
rect 513728 392363 513848 392529
rect 513728 392329 513771 392363
rect 513805 392329 513848 392363
rect 513728 392163 513848 392329
rect 513728 392129 513771 392163
rect 513805 392129 513848 392163
rect 513728 391963 513848 392129
rect 513728 391929 513771 391963
rect 513805 391929 513848 391963
rect 513728 391763 513848 391929
rect 513728 391729 513771 391763
rect 513805 391729 513848 391763
rect 513728 391563 513848 391729
rect 513728 391529 513771 391563
rect 513805 391529 513848 391563
rect 513728 391363 513848 391529
rect 513728 391329 513771 391363
rect 513805 391329 513848 391363
rect 513728 391163 513848 391329
rect 513728 391129 513771 391163
rect 513805 391129 513848 391163
rect 513728 390963 513848 391129
rect 511848 390763 511968 390929
rect 512709 390927 513673 390938
rect 511848 390729 511891 390763
rect 511925 390729 511968 390763
rect 511848 387569 511968 390729
rect 512147 390920 513673 390927
rect 512147 390526 512159 390920
rect 512697 390526 513119 390920
rect 513657 390526 513673 390920
rect 512147 390517 513673 390526
rect 512709 390506 513673 390517
rect 513728 390929 513771 390963
rect 513805 390929 513848 390963
rect 513728 390763 513848 390929
rect 513728 390729 513771 390763
rect 513805 390729 513848 390763
rect 513100 390462 513152 390468
rect 513100 390404 513152 390410
rect 513112 387741 513140 390404
rect 511848 387535 511891 387569
rect 511925 387535 511968 387569
rect 511848 387369 511968 387535
rect 511848 387335 511891 387369
rect 511925 387335 511968 387369
rect 511848 387169 511968 387335
rect 512147 387733 512709 387741
rect 512147 387339 512159 387733
rect 512697 387339 512709 387733
rect 512147 387331 512709 387339
rect 513107 387733 513669 387741
rect 513107 387339 513119 387733
rect 513657 387339 513669 387733
rect 513107 387331 513669 387339
rect 513728 387569 513848 390729
rect 513728 387535 513771 387569
rect 513805 387535 513848 387569
rect 513728 387369 513848 387535
rect 513728 387335 513771 387369
rect 513805 387335 513848 387369
rect 511848 387135 511891 387169
rect 511925 387135 511968 387169
rect 511848 386969 511968 387135
rect 511848 386935 511891 386969
rect 511925 386935 511968 386969
rect 511848 386769 511968 386935
rect 511848 386735 511891 386769
rect 511925 386735 511968 386769
rect 511848 386569 511968 386735
rect 511848 386535 511891 386569
rect 511925 386535 511968 386569
rect 511848 386369 511968 386535
rect 511848 386335 511891 386369
rect 511925 386335 511968 386369
rect 511848 386169 511968 386335
rect 511848 386135 511891 386169
rect 511925 386135 511968 386169
rect 511848 385969 511968 386135
rect 511848 385935 511891 385969
rect 511925 385935 511968 385969
rect 511848 385769 511968 385935
rect 511848 385735 511891 385769
rect 511925 385735 511968 385769
rect 513728 387169 513848 387335
rect 513728 387135 513771 387169
rect 513805 387135 513848 387169
rect 513728 386969 513848 387135
rect 513728 386935 513771 386969
rect 513805 386935 513848 386969
rect 513728 386769 513848 386935
rect 513728 386735 513771 386769
rect 513805 386735 513848 386769
rect 513728 386569 513848 386735
rect 513728 386535 513771 386569
rect 513805 386535 513848 386569
rect 513728 386369 513848 386535
rect 513728 386335 513771 386369
rect 513805 386335 513848 386369
rect 513728 386169 513848 386335
rect 513728 386135 513771 386169
rect 513805 386135 513848 386169
rect 513728 385969 513848 386135
rect 513728 385935 513771 385969
rect 513805 385935 513848 385969
rect 513728 385769 513848 385935
rect 511848 385569 511968 385735
rect 512709 385733 513673 385744
rect 511848 385535 511891 385569
rect 511925 385535 511968 385569
rect 511848 384843 511968 385535
rect 512147 385726 513673 385733
rect 512147 385332 512159 385726
rect 512697 385332 513119 385726
rect 513657 385332 513673 385726
rect 512147 385323 513673 385332
rect 512709 385312 513673 385323
rect 513728 385735 513771 385769
rect 513805 385735 513848 385769
rect 513728 385569 513848 385735
rect 513728 385535 513771 385569
rect 513805 385535 513848 385569
rect 511848 384809 511891 384843
rect 511925 384809 511968 384843
rect 511848 384443 511968 384809
rect 511848 384409 511891 384443
rect 511925 384409 511968 384443
rect 511848 384043 511968 384409
rect 511848 384009 511891 384043
rect 511925 384009 511968 384043
rect 511848 383643 511968 384009
rect 511848 383609 511891 383643
rect 511925 383609 511968 383643
rect 511848 383243 511968 383609
rect 511848 383209 511891 383243
rect 511925 383209 511968 383243
rect 511848 382843 511968 383209
rect 511848 382809 511891 382843
rect 511925 382809 511968 382843
rect 511848 382443 511968 382809
rect 511848 382409 511891 382443
rect 511925 382409 511968 382443
rect 511848 382043 511968 382409
rect 511848 382009 511891 382043
rect 511925 382009 511968 382043
rect 511848 381643 511968 382009
rect 511848 381609 511891 381643
rect 511925 381609 511968 381643
rect 511848 381538 511968 381609
rect 511848 381486 511876 381538
rect 511928 381486 511968 381538
rect 511848 381243 511968 381486
rect 511848 381209 511891 381243
rect 511925 381209 511968 381243
rect 511848 380843 511968 381209
rect 511848 380809 511891 380843
rect 511925 380809 511968 380843
rect 511848 380443 511968 380809
rect 511848 380409 511891 380443
rect 511925 380409 511968 380443
rect 511848 380043 511968 380409
rect 511848 380009 511891 380043
rect 511925 380009 511968 380043
rect 511848 379643 511968 380009
rect 511848 379609 511891 379643
rect 511925 379609 511968 379643
rect 511848 379243 511968 379609
rect 511848 379209 511891 379243
rect 511925 379209 511968 379243
rect 511848 378843 511968 379209
rect 511848 378809 511891 378843
rect 511925 378809 511968 378843
rect 511848 378443 511968 378809
rect 511848 378409 511891 378443
rect 511925 378409 511968 378443
rect 511848 378043 511968 378409
rect 511848 378009 511891 378043
rect 511925 378009 511968 378043
rect 511848 377299 511968 378009
rect 513728 384843 513848 385535
rect 513728 384809 513771 384843
rect 513805 384809 513848 384843
rect 513728 384443 513848 384809
rect 513728 384409 513771 384443
rect 513805 384409 513848 384443
rect 513728 384043 513848 384409
rect 513728 384009 513771 384043
rect 513805 384009 513848 384043
rect 513728 383643 513848 384009
rect 513728 383609 513771 383643
rect 513805 383609 513848 383643
rect 513728 383243 513848 383609
rect 513728 383209 513771 383243
rect 513805 383209 513848 383243
rect 513728 382843 513848 383209
rect 513728 382809 513771 382843
rect 513805 382809 513848 382843
rect 513728 382443 513848 382809
rect 513728 382409 513771 382443
rect 513805 382409 513848 382443
rect 513728 382043 513848 382409
rect 513728 382009 513771 382043
rect 513805 382009 513848 382043
rect 513728 381643 513848 382009
rect 513728 381609 513771 381643
rect 513805 381609 513848 381643
rect 513728 381243 513848 381609
rect 513728 381209 513771 381243
rect 513805 381209 513848 381243
rect 513728 380843 513848 381209
rect 513728 380809 513771 380843
rect 513805 380809 513848 380843
rect 513728 380443 513848 380809
rect 513728 380409 513771 380443
rect 513805 380409 513848 380443
rect 513728 380043 513848 380409
rect 513728 380009 513771 380043
rect 513805 380009 513848 380043
rect 513728 379643 513848 380009
rect 513728 379609 513771 379643
rect 513805 379609 513848 379643
rect 513728 379243 513848 379609
rect 513728 379209 513771 379243
rect 513805 379209 513848 379243
rect 513728 378843 513848 379209
rect 513728 378809 513771 378843
rect 513805 378809 513848 378843
rect 513728 378443 513848 378809
rect 513728 378409 513771 378443
rect 513805 378409 513848 378443
rect 513728 378043 513848 378409
rect 513728 378009 513771 378043
rect 513805 378009 513848 378043
rect 512143 377435 513433 377441
rect 512143 377401 512159 377435
rect 512193 377401 512231 377435
rect 512265 377401 512303 377435
rect 512337 377401 512375 377435
rect 512409 377401 512447 377435
rect 512481 377401 512519 377435
rect 512553 377401 512591 377435
rect 512625 377401 512663 377435
rect 512697 377401 512735 377435
rect 512769 377401 512807 377435
rect 512841 377401 512879 377435
rect 512913 377401 512951 377435
rect 512985 377401 513023 377435
rect 513057 377401 513095 377435
rect 513129 377401 513167 377435
rect 513201 377401 513239 377435
rect 513273 377401 513311 377435
rect 513345 377401 513383 377435
rect 513417 377401 513433 377435
rect 512143 377395 513433 377401
rect 511848 377265 511891 377299
rect 511925 377265 511968 377299
rect 511848 376899 511968 377265
rect 513728 377299 513848 378009
rect 513728 377265 513771 377299
rect 513805 377265 513848 377299
rect 512143 376977 513433 376983
rect 512143 376943 512159 376977
rect 512193 376943 512231 376977
rect 512265 376943 512303 376977
rect 512337 376943 512375 376977
rect 512409 376943 512447 376977
rect 512481 376943 512519 376977
rect 512553 376943 512591 376977
rect 512625 376943 512663 376977
rect 512697 376943 512735 376977
rect 512769 376943 512807 376977
rect 512841 376943 512879 376977
rect 512913 376943 512951 376977
rect 512985 376943 513023 376977
rect 513057 376943 513095 376977
rect 513129 376943 513167 376977
rect 513201 376943 513239 376977
rect 513273 376943 513311 376977
rect 513345 376943 513383 376977
rect 513417 376943 513433 376977
rect 512143 376937 513433 376943
rect 511848 376865 511891 376899
rect 511925 376865 511968 376899
rect 511848 376499 511968 376865
rect 513728 376899 513848 377265
rect 513728 376865 513771 376899
rect 513805 376865 513848 376899
rect 511848 376465 511891 376499
rect 511925 376465 511968 376499
rect 512143 376519 513433 376525
rect 512143 376485 512159 376519
rect 512193 376485 512231 376519
rect 512265 376485 512303 376519
rect 512337 376485 512375 376519
rect 512409 376485 512447 376519
rect 512481 376485 512519 376519
rect 512553 376485 512591 376519
rect 512625 376485 512663 376519
rect 512697 376485 512735 376519
rect 512769 376485 512807 376519
rect 512841 376485 512879 376519
rect 512913 376485 512951 376519
rect 512985 376485 513023 376519
rect 513057 376485 513095 376519
rect 513129 376485 513167 376519
rect 513201 376485 513239 376519
rect 513273 376485 513311 376519
rect 513345 376485 513383 376519
rect 513417 376485 513433 376519
rect 512143 376479 513433 376485
rect 513728 376499 513848 376865
rect 511848 376099 511968 376465
rect 513728 376465 513771 376499
rect 513805 376465 513848 376499
rect 513656 376392 513684 376447
rect 513511 376377 513557 376389
rect 513511 376343 513517 376377
rect 513551 376374 513557 376377
rect 513644 376386 513696 376392
rect 513551 376346 513644 376374
rect 513551 376343 513557 376346
rect 513511 376331 513557 376343
rect 513644 376328 513696 376334
rect 511848 376065 511891 376099
rect 511925 376065 511968 376099
rect 513728 376099 513848 376465
rect 511848 375699 511968 376065
rect 512143 376061 513433 376067
rect 512143 376027 512159 376061
rect 512193 376027 512231 376061
rect 512265 376027 512303 376061
rect 512337 376027 512375 376061
rect 512409 376027 512447 376061
rect 512481 376027 512519 376061
rect 512553 376027 512591 376061
rect 512625 376027 512663 376061
rect 512697 376027 512735 376061
rect 512769 376027 512807 376061
rect 512841 376027 512879 376061
rect 512913 376027 512951 376061
rect 512985 376027 513023 376061
rect 513057 376027 513095 376061
rect 513129 376027 513167 376061
rect 513201 376027 513239 376061
rect 513273 376027 513311 376061
rect 513345 376027 513383 376061
rect 513417 376027 513433 376061
rect 512143 376021 513433 376027
rect 513728 376065 513771 376099
rect 513805 376065 513848 376099
rect 511848 375665 511891 375699
rect 511925 375665 511968 375699
rect 511848 375299 511968 375665
rect 513728 375699 513848 376065
rect 513728 375665 513771 375699
rect 513805 375665 513848 375699
rect 512143 375603 513433 375609
rect 512143 375569 512159 375603
rect 512193 375569 512231 375603
rect 512265 375569 512303 375603
rect 512337 375569 512375 375603
rect 512409 375569 512447 375603
rect 512481 375569 512519 375603
rect 512553 375569 512591 375603
rect 512625 375569 512663 375603
rect 512697 375569 512735 375603
rect 512769 375569 512807 375603
rect 512841 375569 512879 375603
rect 512913 375569 512951 375603
rect 512985 375569 513023 375603
rect 513057 375569 513095 375603
rect 513129 375569 513167 375603
rect 513201 375569 513239 375603
rect 513273 375569 513311 375603
rect 513345 375569 513383 375603
rect 513417 375569 513433 375603
rect 512143 375563 513433 375569
rect 511848 375265 511891 375299
rect 511925 375265 511968 375299
rect 511848 374899 511968 375265
rect 513728 375299 513848 375665
rect 513728 375265 513771 375299
rect 513805 375265 513848 375299
rect 512143 375145 513433 375151
rect 512143 375111 512159 375145
rect 512193 375111 512231 375145
rect 512265 375111 512303 375145
rect 512337 375111 512375 375145
rect 512409 375111 512447 375145
rect 512481 375111 512519 375145
rect 512553 375111 512591 375145
rect 512625 375111 512663 375145
rect 512697 375111 512735 375145
rect 512769 375111 512807 375145
rect 512841 375111 512879 375145
rect 512913 375111 512951 375145
rect 512985 375111 513023 375145
rect 513057 375111 513095 375145
rect 513129 375111 513167 375145
rect 513201 375111 513239 375145
rect 513273 375111 513311 375145
rect 513345 375111 513383 375145
rect 513417 375111 513433 375145
rect 512143 375105 513433 375111
rect 511848 374865 511891 374899
rect 511925 374865 511968 374899
rect 511848 374626 511968 374865
rect 513728 374899 513848 375265
rect 513728 374865 513771 374899
rect 513805 374865 513848 374899
rect 512143 374687 513433 374693
rect 512143 374653 512159 374687
rect 512193 374653 512231 374687
rect 512265 374653 512303 374687
rect 512337 374653 512375 374687
rect 512409 374653 512447 374687
rect 512481 374653 512519 374687
rect 512553 374653 512591 374687
rect 512625 374653 512663 374687
rect 512697 374653 512735 374687
rect 512769 374653 512807 374687
rect 512841 374653 512879 374687
rect 512913 374653 512951 374687
rect 512985 374653 513023 374687
rect 513057 374653 513095 374687
rect 513129 374653 513167 374687
rect 513201 374653 513239 374687
rect 513273 374653 513311 374687
rect 513345 374653 513383 374687
rect 513417 374653 513433 374687
rect 512143 374647 513433 374653
rect 512055 374629 512101 374641
rect 512055 374626 512061 374629
rect 511848 374598 512061 374626
rect 511848 372987 511968 374598
rect 512055 374595 512061 374598
rect 512095 374595 512101 374629
rect 512055 374583 512101 374595
rect 511848 372953 511891 372987
rect 511925 372953 511968 372987
rect 511848 372787 511968 372953
rect 511848 372753 511891 372787
rect 511925 372753 511968 372787
rect 511848 372587 511968 372753
rect 511848 372553 511891 372587
rect 511925 372553 511968 372587
rect 511848 372387 511968 372553
rect 511848 372353 511891 372387
rect 511925 372353 511968 372387
rect 511848 372187 511968 372353
rect 511848 372153 511891 372187
rect 511925 372153 511968 372187
rect 511848 371987 511968 372153
rect 511848 371953 511891 371987
rect 511925 371953 511968 371987
rect 511848 371787 511968 371953
rect 511848 371753 511891 371787
rect 511925 371753 511968 371787
rect 511848 371587 511968 371753
rect 511848 371553 511891 371587
rect 511925 371553 511968 371587
rect 511848 371387 511968 371553
rect 511848 371353 511891 371387
rect 511925 371353 511968 371387
rect 511848 371187 511968 371353
rect 511848 371153 511891 371187
rect 511925 371153 511968 371187
rect 511848 370987 511968 371153
rect 511848 370953 511891 370987
rect 511925 370953 511968 370987
rect 511848 370787 511968 370953
rect 511848 370753 511891 370787
rect 511925 370753 511968 370787
rect 511848 370587 511968 370753
rect 511848 370553 511891 370587
rect 511925 370553 511968 370587
rect 511848 370387 511968 370553
rect 511848 370353 511891 370387
rect 511925 370353 511968 370387
rect 511848 370187 511968 370353
rect 511848 370153 511891 370187
rect 511925 370153 511968 370187
rect 511848 369987 511968 370153
rect 511848 369953 511891 369987
rect 511925 369953 511968 369987
rect 511848 369787 511968 369953
rect 511848 369753 511891 369787
rect 511925 369753 511968 369787
rect 511848 369587 511968 369753
rect 511848 369553 511891 369587
rect 511925 369553 511968 369587
rect 511848 369387 511968 369553
rect 511848 369353 511891 369387
rect 511925 369353 511968 369387
rect 511848 369187 511968 369353
rect 511848 369153 511891 369187
rect 511925 369153 511968 369187
rect 511848 368987 511968 369153
rect 511848 368953 511891 368987
rect 511925 368953 511968 368987
rect 511848 368787 511968 368953
rect 511848 368753 511891 368787
rect 511925 368753 511968 368787
rect 511848 368587 511968 368753
rect 511848 368553 511891 368587
rect 511925 368553 511968 368587
rect 511848 368387 511968 368553
rect 511848 368353 511891 368387
rect 511925 368353 511968 368387
rect 511848 368187 511968 368353
rect 511848 368153 511891 368187
rect 511925 368153 511968 368187
rect 511848 367987 511968 368153
rect 511848 367953 511891 367987
rect 511925 367953 511968 367987
rect 511848 367787 511968 367953
rect 511848 367753 511891 367787
rect 511925 367753 511968 367787
rect 511848 367587 511968 367753
rect 511848 367553 511891 367587
rect 511925 367553 511968 367587
rect 511848 367387 511968 367553
rect 511848 367353 511891 367387
rect 511925 367353 511968 367387
rect 511848 367187 511968 367353
rect 511848 367153 511891 367187
rect 511925 367153 511968 367187
rect 511848 366987 511968 367153
rect 511848 366953 511891 366987
rect 511925 366953 511968 366987
rect 511848 366787 511968 366953
rect 511848 366753 511891 366787
rect 511925 366753 511968 366787
rect 511848 366587 511968 366753
rect 511848 366553 511891 366587
rect 511925 366553 511968 366587
rect 511848 366387 511968 366553
rect 511848 366353 511891 366387
rect 511925 366353 511968 366387
rect 511848 366187 511968 366353
rect 511848 366153 511891 366187
rect 511925 366153 511968 366187
rect 511848 365987 511968 366153
rect 511848 365953 511891 365987
rect 511925 365953 511968 365987
rect 511848 365787 511968 365953
rect 511848 365753 511891 365787
rect 511925 365753 511968 365787
rect 511848 365587 511968 365753
rect 511848 365553 511891 365587
rect 511925 365553 511968 365587
rect 511848 365387 511968 365553
rect 511848 365353 511891 365387
rect 511925 365353 511968 365387
rect 511848 365187 511968 365353
rect 511848 365153 511891 365187
rect 511925 365153 511968 365187
rect 511848 364987 511968 365153
rect 511848 364953 511891 364987
rect 511925 364953 511968 364987
rect 511848 364787 511968 364953
rect 511848 364753 511891 364787
rect 511925 364753 511968 364787
rect 511848 364587 511968 364753
rect 511848 364553 511891 364587
rect 511925 364553 511968 364587
rect 511848 364387 511968 364553
rect 511848 364353 511891 364387
rect 511925 364353 511968 364387
rect 511848 364187 511968 364353
rect 511848 364153 511891 364187
rect 511925 364153 511968 364187
rect 511848 363987 511968 364153
rect 511848 363953 511891 363987
rect 511925 363953 511968 363987
rect 511848 363787 511968 363953
rect 511848 363753 511891 363787
rect 511925 363753 511968 363787
rect 511848 363587 511968 363753
rect 511848 363553 511891 363587
rect 511925 363553 511968 363587
rect 511848 363387 511968 363553
rect 511848 363353 511891 363387
rect 511925 363353 511968 363387
rect 511848 363187 511968 363353
rect 511848 363153 511891 363187
rect 511925 363153 511968 363187
rect 511848 362987 511968 363153
rect 511848 362953 511891 362987
rect 511925 362953 511968 362987
rect 511848 362787 511968 362953
rect 511848 362753 511891 362787
rect 511925 362753 511968 362787
rect 511848 362587 511968 362753
rect 511848 362553 511891 362587
rect 511925 362553 511968 362587
rect 511848 361476 511968 362553
rect 512218 373124 512288 373144
rect 512218 373090 512224 373124
rect 512258 373090 512288 373124
rect 512218 373034 512288 373090
rect 512218 373000 512224 373034
rect 512258 373000 512288 373034
rect 512218 372944 512288 373000
rect 513728 372987 513848 374865
rect 512218 372910 512224 372944
rect 512258 372910 512288 372944
rect 512218 372854 512288 372910
rect 512218 372820 512224 372854
rect 512258 372820 512288 372854
rect 512218 372786 512288 372820
rect 512368 372960 512438 372980
rect 512368 372926 512384 372960
rect 512418 372926 512438 372960
rect 512368 372870 512438 372926
rect 512368 372836 512384 372870
rect 512418 372836 512438 372870
rect 512368 372804 512438 372836
rect 513728 372953 513771 372987
rect 513805 372953 513848 372987
rect 512352 372798 512438 372804
rect 512218 372764 512352 372786
rect 512404 372780 512438 372798
rect 512218 372730 512224 372764
rect 512258 372758 512352 372764
rect 512258 372730 512288 372758
rect 512418 372746 512438 372780
rect 512352 372740 512438 372746
rect 512218 372674 512288 372730
rect 512218 372640 512224 372674
rect 512258 372640 512288 372674
rect 512218 372584 512288 372640
rect 512218 372550 512224 372584
rect 512258 372550 512288 372584
rect 512218 372494 512288 372550
rect 512218 372460 512224 372494
rect 512258 372460 512288 372494
rect 512218 372404 512288 372460
rect 512218 372370 512224 372404
rect 512258 372370 512288 372404
rect 512218 372314 512288 372370
rect 512218 372280 512224 372314
rect 512258 372280 512288 372314
rect 512218 372224 512288 372280
rect 512218 372190 512224 372224
rect 512258 372190 512288 372224
rect 512218 372134 512288 372190
rect 512218 372100 512224 372134
rect 512258 372100 512288 372134
rect 512218 372044 512288 372100
rect 512218 372010 512224 372044
rect 512258 372010 512288 372044
rect 512218 371954 512288 372010
rect 512218 371920 512224 371954
rect 512258 371920 512288 371954
rect 512218 371784 512288 371920
rect 512218 371750 512224 371784
rect 512258 371750 512288 371784
rect 512218 371694 512288 371750
rect 512218 371660 512224 371694
rect 512258 371660 512288 371694
rect 512218 371604 512288 371660
rect 512218 371570 512224 371604
rect 512258 371570 512288 371604
rect 512218 371514 512288 371570
rect 512218 371480 512224 371514
rect 512258 371480 512288 371514
rect 512218 371424 512288 371480
rect 512218 371390 512224 371424
rect 512258 371390 512288 371424
rect 512218 371334 512288 371390
rect 512218 371300 512224 371334
rect 512258 371300 512288 371334
rect 512218 371244 512288 371300
rect 512218 371210 512224 371244
rect 512258 371210 512288 371244
rect 512218 371154 512288 371210
rect 512218 371120 512224 371154
rect 512258 371120 512288 371154
rect 512218 371064 512288 371120
rect 512218 371030 512224 371064
rect 512258 371030 512288 371064
rect 512218 370974 512288 371030
rect 512218 370940 512224 370974
rect 512258 370940 512288 370974
rect 512218 370884 512288 370940
rect 512218 370850 512224 370884
rect 512258 370850 512288 370884
rect 512218 370794 512288 370850
rect 512218 370760 512224 370794
rect 512258 370760 512288 370794
rect 512218 370704 512288 370760
rect 512218 370670 512224 370704
rect 512258 370670 512288 370704
rect 512218 370614 512288 370670
rect 512218 370580 512224 370614
rect 512258 370580 512288 370614
rect 512218 370444 512288 370580
rect 512218 370410 512224 370444
rect 512258 370410 512288 370444
rect 512218 370354 512288 370410
rect 512218 370320 512224 370354
rect 512258 370320 512288 370354
rect 512218 370264 512288 370320
rect 512218 370230 512224 370264
rect 512258 370230 512288 370264
rect 512218 370174 512288 370230
rect 512218 370140 512224 370174
rect 512258 370140 512288 370174
rect 512218 370084 512288 370140
rect 512218 370050 512224 370084
rect 512258 370050 512288 370084
rect 512218 369994 512288 370050
rect 512218 369960 512224 369994
rect 512258 369960 512288 369994
rect 512218 369904 512288 369960
rect 512218 369870 512224 369904
rect 512258 369870 512288 369904
rect 512218 369814 512288 369870
rect 512218 369780 512224 369814
rect 512258 369780 512288 369814
rect 512218 369724 512288 369780
rect 512218 369690 512224 369724
rect 512258 369690 512288 369724
rect 512218 369634 512288 369690
rect 512218 369600 512224 369634
rect 512258 369600 512288 369634
rect 512218 369544 512288 369600
rect 512218 369510 512224 369544
rect 512258 369510 512288 369544
rect 512218 369454 512288 369510
rect 512218 369420 512224 369454
rect 512258 369420 512288 369454
rect 512218 369364 512288 369420
rect 512218 369330 512224 369364
rect 512258 369330 512288 369364
rect 512218 369274 512288 369330
rect 512218 369240 512224 369274
rect 512258 369240 512288 369274
rect 512218 369104 512288 369240
rect 512218 369070 512224 369104
rect 512258 369070 512288 369104
rect 512218 369014 512288 369070
rect 512218 368980 512224 369014
rect 512258 368980 512288 369014
rect 512218 368924 512288 368980
rect 512218 368890 512224 368924
rect 512258 368890 512288 368924
rect 512218 368834 512288 368890
rect 512218 368800 512224 368834
rect 512258 368800 512288 368834
rect 512218 368744 512288 368800
rect 512218 368710 512224 368744
rect 512258 368710 512288 368744
rect 512218 368654 512288 368710
rect 512218 368620 512224 368654
rect 512258 368620 512288 368654
rect 512218 368564 512288 368620
rect 512218 368530 512224 368564
rect 512258 368530 512288 368564
rect 512218 368474 512288 368530
rect 512218 368440 512224 368474
rect 512258 368440 512288 368474
rect 512218 368384 512288 368440
rect 512218 368350 512224 368384
rect 512258 368350 512288 368384
rect 512218 368294 512288 368350
rect 512218 368260 512224 368294
rect 512258 368260 512288 368294
rect 512218 368204 512288 368260
rect 512218 368170 512224 368204
rect 512258 368170 512288 368204
rect 512218 368114 512288 368170
rect 512218 368080 512224 368114
rect 512258 368080 512288 368114
rect 512218 368024 512288 368080
rect 512218 367990 512224 368024
rect 512258 367990 512288 368024
rect 512218 367934 512288 367990
rect 512218 367900 512224 367934
rect 512258 367900 512288 367934
rect 512218 367764 512288 367900
rect 512218 367730 512224 367764
rect 512258 367730 512288 367764
rect 512218 367674 512288 367730
rect 512218 367640 512224 367674
rect 512258 367640 512288 367674
rect 512218 367584 512288 367640
rect 512218 367550 512224 367584
rect 512258 367550 512288 367584
rect 512218 367494 512288 367550
rect 512218 367460 512224 367494
rect 512258 367460 512288 367494
rect 512218 367404 512288 367460
rect 512218 367370 512224 367404
rect 512258 367370 512288 367404
rect 512218 367314 512288 367370
rect 512218 367280 512224 367314
rect 512258 367280 512288 367314
rect 512218 367224 512288 367280
rect 512218 367190 512224 367224
rect 512258 367190 512288 367224
rect 512218 367134 512288 367190
rect 512218 367100 512224 367134
rect 512258 367100 512288 367134
rect 512218 367044 512288 367100
rect 512218 367010 512224 367044
rect 512258 367010 512288 367044
rect 512218 366954 512288 367010
rect 512218 366920 512224 366954
rect 512258 366920 512288 366954
rect 512218 366864 512288 366920
rect 512218 366830 512224 366864
rect 512258 366830 512288 366864
rect 512218 366774 512288 366830
rect 512218 366740 512224 366774
rect 512258 366740 512288 366774
rect 512218 366684 512288 366740
rect 512218 366650 512224 366684
rect 512258 366650 512288 366684
rect 512218 366594 512288 366650
rect 512218 366560 512224 366594
rect 512258 366560 512288 366594
rect 512218 366424 512288 366560
rect 512218 366390 512224 366424
rect 512258 366390 512288 366424
rect 512218 366334 512288 366390
rect 512218 366300 512224 366334
rect 512258 366300 512288 366334
rect 512218 366244 512288 366300
rect 512218 366210 512224 366244
rect 512258 366210 512288 366244
rect 512218 366154 512288 366210
rect 512218 366120 512224 366154
rect 512258 366120 512288 366154
rect 512218 366064 512288 366120
rect 512218 366030 512224 366064
rect 512258 366030 512288 366064
rect 512218 365974 512288 366030
rect 512218 365940 512224 365974
rect 512258 365940 512288 365974
rect 512218 365884 512288 365940
rect 512218 365850 512224 365884
rect 512258 365850 512288 365884
rect 512218 365794 512288 365850
rect 512218 365760 512224 365794
rect 512258 365760 512288 365794
rect 512218 365704 512288 365760
rect 512218 365670 512224 365704
rect 512258 365670 512288 365704
rect 512218 365614 512288 365670
rect 512218 365580 512224 365614
rect 512258 365580 512288 365614
rect 512218 365524 512288 365580
rect 512218 365490 512224 365524
rect 512258 365490 512288 365524
rect 512218 365434 512288 365490
rect 512218 365400 512224 365434
rect 512258 365400 512288 365434
rect 512218 365344 512288 365400
rect 512218 365310 512224 365344
rect 512258 365310 512288 365344
rect 512218 365254 512288 365310
rect 512218 365220 512224 365254
rect 512258 365220 512288 365254
rect 512218 365084 512288 365220
rect 512218 365050 512224 365084
rect 512258 365050 512288 365084
rect 512218 364994 512288 365050
rect 512218 364960 512224 364994
rect 512258 364960 512288 364994
rect 512218 364904 512288 364960
rect 512218 364870 512224 364904
rect 512258 364870 512288 364904
rect 512218 364814 512288 364870
rect 512218 364780 512224 364814
rect 512258 364780 512288 364814
rect 512218 364724 512288 364780
rect 512218 364690 512224 364724
rect 512258 364690 512288 364724
rect 512218 364634 512288 364690
rect 512218 364600 512224 364634
rect 512258 364600 512288 364634
rect 512218 364544 512288 364600
rect 512218 364510 512224 364544
rect 512258 364510 512288 364544
rect 512218 364454 512288 364510
rect 512218 364420 512224 364454
rect 512258 364420 512288 364454
rect 512218 364364 512288 364420
rect 512218 364330 512224 364364
rect 512258 364330 512288 364364
rect 512218 364274 512288 364330
rect 512218 364240 512224 364274
rect 512258 364240 512288 364274
rect 512218 364184 512288 364240
rect 512218 364150 512224 364184
rect 512258 364150 512288 364184
rect 512218 364094 512288 364150
rect 512218 364060 512224 364094
rect 512258 364060 512288 364094
rect 512218 364004 512288 364060
rect 512218 363970 512224 364004
rect 512258 363970 512288 364004
rect 512218 363914 512288 363970
rect 512218 363880 512224 363914
rect 512258 363880 512288 363914
rect 512218 363744 512288 363880
rect 512218 363710 512224 363744
rect 512258 363710 512288 363744
rect 512218 363654 512288 363710
rect 512218 363620 512224 363654
rect 512258 363620 512288 363654
rect 512218 363564 512288 363620
rect 512218 363530 512224 363564
rect 512258 363530 512288 363564
rect 512218 363474 512288 363530
rect 512218 363440 512224 363474
rect 512258 363440 512288 363474
rect 512218 363384 512288 363440
rect 512218 363350 512224 363384
rect 512258 363350 512288 363384
rect 512218 363294 512288 363350
rect 512218 363260 512224 363294
rect 512258 363260 512288 363294
rect 512218 363204 512288 363260
rect 512218 363170 512224 363204
rect 512258 363170 512288 363204
rect 512218 363114 512288 363170
rect 512218 363080 512224 363114
rect 512258 363080 512288 363114
rect 512218 363024 512288 363080
rect 512218 362990 512224 363024
rect 512258 362990 512288 363024
rect 512218 362934 512288 362990
rect 512218 362900 512224 362934
rect 512258 362900 512288 362934
rect 512218 362844 512288 362900
rect 512218 362810 512224 362844
rect 512258 362810 512288 362844
rect 512218 362754 512288 362810
rect 512218 362720 512224 362754
rect 512258 362720 512288 362754
rect 512218 362664 512288 362720
rect 512218 362630 512224 362664
rect 512258 362630 512288 362664
rect 512368 372690 512438 372740
rect 512368 372656 512384 372690
rect 512418 372656 512438 372690
rect 512368 372600 512438 372656
rect 512368 372566 512384 372600
rect 512418 372566 512438 372600
rect 512368 372510 512438 372566
rect 512368 372476 512384 372510
rect 512418 372476 512438 372510
rect 512368 372420 512438 372476
rect 512368 372386 512384 372420
rect 512418 372386 512438 372420
rect 512368 372330 512438 372386
rect 512368 372296 512384 372330
rect 512418 372296 512438 372330
rect 512368 372240 512438 372296
rect 512368 372206 512384 372240
rect 512418 372206 512438 372240
rect 512368 372150 512438 372206
rect 512368 372116 512384 372150
rect 512418 372116 512438 372150
rect 512368 372060 512438 372116
rect 512368 372026 512384 372060
rect 512418 372026 512438 372060
rect 512368 371620 512438 372026
rect 512368 371586 512384 371620
rect 512418 371586 512438 371620
rect 512368 371530 512438 371586
rect 512368 371496 512384 371530
rect 512418 371496 512438 371530
rect 512368 371440 512438 371496
rect 512368 371406 512384 371440
rect 512418 371406 512438 371440
rect 512368 371350 512438 371406
rect 512368 371316 512384 371350
rect 512418 371316 512438 371350
rect 512368 371260 512438 371316
rect 512368 371226 512384 371260
rect 512418 371226 512438 371260
rect 512368 371170 512438 371226
rect 512368 371136 512384 371170
rect 512418 371136 512438 371170
rect 512368 371080 512438 371136
rect 512368 371046 512384 371080
rect 512418 371046 512438 371080
rect 512368 370990 512438 371046
rect 512368 370956 512384 370990
rect 512418 370956 512438 370990
rect 512368 370900 512438 370956
rect 512368 370866 512384 370900
rect 512418 370866 512438 370900
rect 512368 370810 512438 370866
rect 512368 370776 512384 370810
rect 512418 370776 512438 370810
rect 512368 370720 512438 370776
rect 512368 370686 512384 370720
rect 512418 370686 512438 370720
rect 512368 370280 512438 370686
rect 512368 370246 512384 370280
rect 512418 370246 512438 370280
rect 512368 370190 512438 370246
rect 512368 370156 512384 370190
rect 512418 370156 512438 370190
rect 512368 370100 512438 370156
rect 512368 370066 512384 370100
rect 512418 370066 512438 370100
rect 512368 370010 512438 370066
rect 512368 369976 512384 370010
rect 512418 369976 512438 370010
rect 512368 369920 512438 369976
rect 512368 369886 512384 369920
rect 512418 369886 512438 369920
rect 512368 369830 512438 369886
rect 512368 369796 512384 369830
rect 512418 369796 512438 369830
rect 512368 369740 512438 369796
rect 512368 369706 512384 369740
rect 512418 369706 512438 369740
rect 512368 369650 512438 369706
rect 512368 369616 512384 369650
rect 512418 369616 512438 369650
rect 512368 369560 512438 369616
rect 512368 369526 512384 369560
rect 512418 369526 512438 369560
rect 512368 369470 512438 369526
rect 512368 369436 512384 369470
rect 512418 369436 512438 369470
rect 512368 369380 512438 369436
rect 512368 369346 512384 369380
rect 512418 369346 512438 369380
rect 512368 368940 512438 369346
rect 512368 368906 512384 368940
rect 512418 368906 512438 368940
rect 512368 368850 512438 368906
rect 512368 368816 512384 368850
rect 512418 368816 512438 368850
rect 512368 368760 512438 368816
rect 512368 368726 512384 368760
rect 512418 368726 512438 368760
rect 512368 368670 512438 368726
rect 512368 368636 512384 368670
rect 512418 368636 512438 368670
rect 512368 368580 512438 368636
rect 512368 368546 512384 368580
rect 512418 368546 512438 368580
rect 512368 368490 512438 368546
rect 512368 368456 512384 368490
rect 512418 368456 512438 368490
rect 512368 368400 512438 368456
rect 512368 368366 512384 368400
rect 512418 368366 512438 368400
rect 512368 368310 512438 368366
rect 512368 368276 512384 368310
rect 512418 368276 512438 368310
rect 512368 368220 512438 368276
rect 512368 368186 512384 368220
rect 512418 368186 512438 368220
rect 512368 368130 512438 368186
rect 512368 368096 512384 368130
rect 512418 368096 512438 368130
rect 512368 368040 512438 368096
rect 512368 368006 512384 368040
rect 512418 368006 512438 368040
rect 512368 367600 512438 368006
rect 512368 367566 512384 367600
rect 512418 367566 512438 367600
rect 512368 367510 512438 367566
rect 512368 367476 512384 367510
rect 512418 367476 512438 367510
rect 512368 367420 512438 367476
rect 512368 367386 512384 367420
rect 512418 367386 512438 367420
rect 512368 367330 512438 367386
rect 512368 367296 512384 367330
rect 512418 367296 512438 367330
rect 512368 367240 512438 367296
rect 512368 367206 512384 367240
rect 512418 367206 512438 367240
rect 512368 367150 512438 367206
rect 512368 367116 512384 367150
rect 512418 367116 512438 367150
rect 512368 367060 512438 367116
rect 512368 367026 512384 367060
rect 512418 367026 512438 367060
rect 512368 366970 512438 367026
rect 512368 366936 512384 366970
rect 512418 366936 512438 366970
rect 512368 366880 512438 366936
rect 512368 366846 512384 366880
rect 512418 366846 512438 366880
rect 512368 366790 512438 366846
rect 512368 366756 512384 366790
rect 512418 366756 512438 366790
rect 512368 366700 512438 366756
rect 512368 366666 512384 366700
rect 512418 366666 512438 366700
rect 512368 366260 512438 366666
rect 512368 366226 512384 366260
rect 512418 366226 512438 366260
rect 512368 366170 512438 366226
rect 512368 366136 512384 366170
rect 512418 366136 512438 366170
rect 512368 366080 512438 366136
rect 512368 366046 512384 366080
rect 512418 366046 512438 366080
rect 512368 365990 512438 366046
rect 512368 365956 512384 365990
rect 512418 365956 512438 365990
rect 512368 365900 512438 365956
rect 512368 365866 512384 365900
rect 512418 365866 512438 365900
rect 512368 365810 512438 365866
rect 512368 365776 512384 365810
rect 512418 365776 512438 365810
rect 512368 365720 512438 365776
rect 512368 365686 512384 365720
rect 512418 365686 512438 365720
rect 512368 365630 512438 365686
rect 512368 365596 512384 365630
rect 512418 365596 512438 365630
rect 512368 365540 512438 365596
rect 512368 365506 512384 365540
rect 512418 365506 512438 365540
rect 512368 365450 512438 365506
rect 512368 365416 512384 365450
rect 512418 365416 512438 365450
rect 512368 365360 512438 365416
rect 512368 365326 512384 365360
rect 512418 365326 512438 365360
rect 512368 364920 512438 365326
rect 512368 364886 512384 364920
rect 512418 364886 512438 364920
rect 512368 364830 512438 364886
rect 512368 364796 512384 364830
rect 512418 364796 512438 364830
rect 512368 364740 512438 364796
rect 512368 364706 512384 364740
rect 512418 364706 512438 364740
rect 512368 364650 512438 364706
rect 512368 364616 512384 364650
rect 512418 364616 512438 364650
rect 512368 364560 512438 364616
rect 512368 364526 512384 364560
rect 512418 364526 512438 364560
rect 512368 364470 512438 364526
rect 512368 364436 512384 364470
rect 512418 364436 512438 364470
rect 512368 364380 512438 364436
rect 512368 364346 512384 364380
rect 512418 364346 512438 364380
rect 512368 364290 512438 364346
rect 512368 364256 512384 364290
rect 512418 364256 512438 364290
rect 512368 364200 512438 364256
rect 512368 364166 512384 364200
rect 512418 364166 512438 364200
rect 512368 364110 512438 364166
rect 512368 364076 512384 364110
rect 512418 364076 512438 364110
rect 512368 364020 512438 364076
rect 512368 363986 512384 364020
rect 512418 363986 512438 364020
rect 512368 363580 512438 363986
rect 512368 363546 512384 363580
rect 512418 363546 512438 363580
rect 512368 363490 512438 363546
rect 512368 363456 512384 363490
rect 512418 363456 512438 363490
rect 512368 363400 512438 363456
rect 512368 363366 512384 363400
rect 512418 363366 512438 363400
rect 512368 363310 512438 363366
rect 512368 363276 512384 363310
rect 512418 363276 512438 363310
rect 512368 363220 512438 363276
rect 512368 363186 512384 363220
rect 512418 363186 512438 363220
rect 512368 363130 512438 363186
rect 512368 363096 512384 363130
rect 512418 363096 512438 363130
rect 512368 363040 512438 363096
rect 512368 363006 512384 363040
rect 512418 363006 512438 363040
rect 512368 362950 512438 363006
rect 512368 362916 512384 362950
rect 512418 362916 512438 362950
rect 512368 362860 512438 362916
rect 512368 362826 512384 362860
rect 512418 362826 512438 362860
rect 512368 362770 512438 362826
rect 512542 372774 513154 372806
rect 512542 372740 512588 372774
rect 512622 372740 512688 372774
rect 512722 372740 512788 372774
rect 512822 372740 512888 372774
rect 512922 372740 512988 372774
rect 513022 372740 513088 372774
rect 513122 372740 513154 372774
rect 512542 372706 513154 372740
rect 512542 372654 512556 372706
rect 512608 372674 513154 372706
rect 512542 372640 512588 372654
rect 512622 372640 512688 372674
rect 512722 372640 512788 372674
rect 512822 372640 512888 372674
rect 512922 372640 512988 372674
rect 513022 372640 513088 372674
rect 513122 372640 513154 372674
rect 512542 372574 513154 372640
rect 512542 372540 512588 372574
rect 512622 372540 512688 372574
rect 512722 372540 512788 372574
rect 512822 372540 512888 372574
rect 512922 372540 512988 372574
rect 513022 372540 513088 372574
rect 513122 372540 513154 372574
rect 512542 372474 513154 372540
rect 512542 372440 512588 372474
rect 512622 372440 512688 372474
rect 512722 372440 512788 372474
rect 512822 372440 512888 372474
rect 512922 372440 512988 372474
rect 513022 372440 513088 372474
rect 513122 372440 513154 372474
rect 512542 372374 513154 372440
rect 512542 372340 512588 372374
rect 512622 372340 512688 372374
rect 512722 372340 512788 372374
rect 512822 372340 512888 372374
rect 512922 372340 512988 372374
rect 513022 372340 513088 372374
rect 513122 372340 513154 372374
rect 512542 372274 513154 372340
rect 512542 372240 512588 372274
rect 512622 372240 512688 372274
rect 512722 372240 512788 372274
rect 512822 372240 512888 372274
rect 512922 372240 512988 372274
rect 513022 372240 513088 372274
rect 513122 372240 513154 372274
rect 512542 371434 513154 372240
rect 512542 371400 512588 371434
rect 512622 371400 512688 371434
rect 512722 371400 512788 371434
rect 512822 371400 512888 371434
rect 512922 371400 512988 371434
rect 513022 371400 513088 371434
rect 513122 371400 513154 371434
rect 512542 371334 513154 371400
rect 512542 371300 512588 371334
rect 512622 371300 512688 371334
rect 512722 371300 512788 371334
rect 512822 371300 512888 371334
rect 512922 371300 512988 371334
rect 513022 371300 513088 371334
rect 513122 371300 513154 371334
rect 512542 371234 513154 371300
rect 512542 371200 512588 371234
rect 512622 371200 512688 371234
rect 512722 371200 512788 371234
rect 512822 371200 512888 371234
rect 512922 371200 512988 371234
rect 513022 371200 513088 371234
rect 513122 371200 513154 371234
rect 512542 371134 513154 371200
rect 512542 371100 512588 371134
rect 512622 371100 512688 371134
rect 512722 371100 512788 371134
rect 512822 371100 512888 371134
rect 512922 371100 512988 371134
rect 513022 371100 513088 371134
rect 513122 371100 513154 371134
rect 512542 371034 513154 371100
rect 512542 371000 512588 371034
rect 512622 371000 512688 371034
rect 512722 371000 512788 371034
rect 512822 371000 512888 371034
rect 512922 371000 512988 371034
rect 513022 371000 513088 371034
rect 513122 371000 513154 371034
rect 512542 370934 513154 371000
rect 512542 370900 512588 370934
rect 512622 370900 512688 370934
rect 512722 370900 512788 370934
rect 512822 370900 512888 370934
rect 512922 370900 512988 370934
rect 513022 370900 513088 370934
rect 513122 370900 513154 370934
rect 512542 370094 513154 370900
rect 512542 370060 512588 370094
rect 512622 370060 512688 370094
rect 512722 370060 512788 370094
rect 512822 370060 512888 370094
rect 512922 370060 512988 370094
rect 513022 370060 513088 370094
rect 513122 370060 513154 370094
rect 512542 369994 513154 370060
rect 512542 369960 512588 369994
rect 512622 369960 512688 369994
rect 512722 369960 512788 369994
rect 512822 369960 512888 369994
rect 512922 369960 512988 369994
rect 513022 369960 513088 369994
rect 513122 369960 513154 369994
rect 512542 369894 513154 369960
rect 512542 369860 512588 369894
rect 512622 369860 512688 369894
rect 512722 369860 512788 369894
rect 512822 369860 512888 369894
rect 512922 369860 512988 369894
rect 513022 369860 513088 369894
rect 513122 369860 513154 369894
rect 512542 369794 513154 369860
rect 512542 369760 512588 369794
rect 512622 369760 512688 369794
rect 512722 369760 512788 369794
rect 512822 369760 512888 369794
rect 512922 369760 512988 369794
rect 513022 369760 513088 369794
rect 513122 369760 513154 369794
rect 512542 369694 513154 369760
rect 512542 369660 512588 369694
rect 512622 369660 512688 369694
rect 512722 369660 512788 369694
rect 512822 369660 512888 369694
rect 512922 369660 512988 369694
rect 513022 369660 513088 369694
rect 513122 369660 513154 369694
rect 512542 369594 513154 369660
rect 512542 369560 512588 369594
rect 512622 369560 512688 369594
rect 512722 369560 512788 369594
rect 512822 369560 512888 369594
rect 512922 369560 512988 369594
rect 513022 369560 513088 369594
rect 513122 369560 513154 369594
rect 512542 368754 513154 369560
rect 512542 368720 512588 368754
rect 512622 368720 512688 368754
rect 512722 368720 512788 368754
rect 512822 368720 512888 368754
rect 512922 368720 512988 368754
rect 513022 368720 513088 368754
rect 513122 368720 513154 368754
rect 512542 368654 513154 368720
rect 512542 368620 512588 368654
rect 512622 368620 512688 368654
rect 512722 368620 512788 368654
rect 512822 368620 512888 368654
rect 512922 368620 512988 368654
rect 513022 368620 513088 368654
rect 513122 368620 513154 368654
rect 512542 368554 513154 368620
rect 512542 368520 512588 368554
rect 512622 368520 512688 368554
rect 512722 368520 512788 368554
rect 512822 368520 512888 368554
rect 512922 368520 512988 368554
rect 513022 368520 513088 368554
rect 513122 368520 513154 368554
rect 512542 368454 513154 368520
rect 512542 368420 512588 368454
rect 512622 368420 512688 368454
rect 512722 368420 512788 368454
rect 512822 368420 512888 368454
rect 512922 368420 512988 368454
rect 513022 368420 513088 368454
rect 513122 368420 513154 368454
rect 512542 368354 513154 368420
rect 512542 368320 512588 368354
rect 512622 368320 512688 368354
rect 512722 368320 512788 368354
rect 512822 368320 512888 368354
rect 512922 368320 512988 368354
rect 513022 368320 513088 368354
rect 513122 368320 513154 368354
rect 512542 368254 513154 368320
rect 512542 368220 512588 368254
rect 512622 368220 512688 368254
rect 512722 368220 512788 368254
rect 512822 368220 512888 368254
rect 512922 368220 512988 368254
rect 513022 368220 513088 368254
rect 513122 368220 513154 368254
rect 512542 367414 513154 368220
rect 512542 367380 512588 367414
rect 512622 367380 512688 367414
rect 512722 367380 512788 367414
rect 512822 367380 512888 367414
rect 512922 367380 512988 367414
rect 513022 367380 513088 367414
rect 513122 367380 513154 367414
rect 512542 367314 513154 367380
rect 512542 367280 512588 367314
rect 512622 367280 512688 367314
rect 512722 367280 512788 367314
rect 512822 367280 512888 367314
rect 512922 367280 512988 367314
rect 513022 367280 513088 367314
rect 513122 367280 513154 367314
rect 512542 367214 513154 367280
rect 512542 367180 512588 367214
rect 512622 367180 512688 367214
rect 512722 367180 512788 367214
rect 512822 367180 512888 367214
rect 512922 367180 512988 367214
rect 513022 367180 513088 367214
rect 513122 367180 513154 367214
rect 512542 367114 513154 367180
rect 512542 367080 512588 367114
rect 512622 367080 512688 367114
rect 512722 367080 512788 367114
rect 512822 367080 512888 367114
rect 512922 367080 512988 367114
rect 513022 367080 513088 367114
rect 513122 367080 513154 367114
rect 512542 367014 513154 367080
rect 512542 366980 512588 367014
rect 512622 366980 512688 367014
rect 512722 366980 512788 367014
rect 512822 366980 512888 367014
rect 512922 366980 512988 367014
rect 513022 366980 513088 367014
rect 513122 366980 513154 367014
rect 512542 366914 513154 366980
rect 512542 366880 512588 366914
rect 512622 366880 512688 366914
rect 512722 366880 512788 366914
rect 512822 366880 512888 366914
rect 512922 366880 512988 366914
rect 513022 366880 513088 366914
rect 513122 366880 513154 366914
rect 512542 366542 513154 366880
rect 512542 366490 513100 366542
rect 513152 366490 513154 366542
rect 512542 366074 513154 366490
rect 512542 366040 512588 366074
rect 512622 366040 512688 366074
rect 512722 366040 512788 366074
rect 512822 366040 512888 366074
rect 512922 366040 512988 366074
rect 513022 366040 513088 366074
rect 513122 366040 513154 366074
rect 512542 365974 513154 366040
rect 512542 365940 512588 365974
rect 512622 365940 512688 365974
rect 512722 365940 512788 365974
rect 512822 365940 512888 365974
rect 512922 365940 512988 365974
rect 513022 365940 513088 365974
rect 513122 365940 513154 365974
rect 512542 365874 513154 365940
rect 512542 365840 512588 365874
rect 512622 365840 512688 365874
rect 512722 365840 512788 365874
rect 512822 365840 512888 365874
rect 512922 365840 512988 365874
rect 513022 365840 513088 365874
rect 513122 365840 513154 365874
rect 512542 365774 513154 365840
rect 512542 365740 512588 365774
rect 512622 365740 512688 365774
rect 512722 365740 512788 365774
rect 512822 365740 512888 365774
rect 512922 365740 512988 365774
rect 513022 365740 513088 365774
rect 513122 365740 513154 365774
rect 512542 365674 513154 365740
rect 512542 365640 512588 365674
rect 512622 365640 512688 365674
rect 512722 365640 512788 365674
rect 512822 365640 512888 365674
rect 512922 365640 512988 365674
rect 513022 365640 513088 365674
rect 513122 365640 513154 365674
rect 512542 365574 513154 365640
rect 512542 365540 512588 365574
rect 512622 365540 512688 365574
rect 512722 365540 512788 365574
rect 512822 365540 512888 365574
rect 512922 365540 512988 365574
rect 513022 365540 513088 365574
rect 513122 365540 513154 365574
rect 512542 364734 513154 365540
rect 512542 364700 512588 364734
rect 512622 364700 512688 364734
rect 512722 364700 512788 364734
rect 512822 364700 512888 364734
rect 512922 364700 512988 364734
rect 513022 364700 513088 364734
rect 513122 364700 513154 364734
rect 512542 364634 513154 364700
rect 512542 364600 512588 364634
rect 512622 364600 512688 364634
rect 512722 364600 512788 364634
rect 512822 364600 512888 364634
rect 512922 364600 512988 364634
rect 513022 364600 513088 364634
rect 513122 364600 513154 364634
rect 512542 364534 513154 364600
rect 512542 364500 512588 364534
rect 512622 364500 512688 364534
rect 512722 364500 512788 364534
rect 512822 364500 512888 364534
rect 512922 364500 512988 364534
rect 513022 364500 513088 364534
rect 513122 364500 513154 364534
rect 512542 364434 513154 364500
rect 512542 364400 512588 364434
rect 512622 364400 512688 364434
rect 512722 364400 512788 364434
rect 512822 364400 512888 364434
rect 512922 364400 512988 364434
rect 513022 364400 513088 364434
rect 513122 364400 513154 364434
rect 512542 364334 513154 364400
rect 512542 364300 512588 364334
rect 512622 364300 512688 364334
rect 512722 364300 512788 364334
rect 512822 364300 512888 364334
rect 512922 364300 512988 364334
rect 513022 364300 513088 364334
rect 513122 364300 513154 364334
rect 512542 364234 513154 364300
rect 512542 364200 512588 364234
rect 512622 364200 512688 364234
rect 512722 364200 512788 364234
rect 512822 364200 512888 364234
rect 512922 364200 512988 364234
rect 513022 364200 513088 364234
rect 513122 364200 513154 364234
rect 512542 363394 513154 364200
rect 512542 363360 512588 363394
rect 512622 363360 512688 363394
rect 512722 363360 512788 363394
rect 512822 363360 512888 363394
rect 512922 363360 512988 363394
rect 513022 363360 513088 363394
rect 513122 363360 513154 363394
rect 512542 363294 513154 363360
rect 512542 363260 512588 363294
rect 512622 363260 512688 363294
rect 512722 363260 512788 363294
rect 512822 363260 512888 363294
rect 512922 363260 512988 363294
rect 513022 363260 513088 363294
rect 513122 363260 513154 363294
rect 512542 363194 513154 363260
rect 512542 363160 512588 363194
rect 512622 363160 512688 363194
rect 512722 363160 512788 363194
rect 512822 363160 512888 363194
rect 512922 363160 512988 363194
rect 513022 363160 513088 363194
rect 513122 363160 513154 363194
rect 512542 363094 513154 363160
rect 512542 363060 512588 363094
rect 512622 363060 512688 363094
rect 512722 363060 512788 363094
rect 512822 363060 512888 363094
rect 512922 363060 512988 363094
rect 513022 363060 513088 363094
rect 513122 363060 513154 363094
rect 512542 362994 513154 363060
rect 512542 362960 512588 362994
rect 512622 362960 512688 362994
rect 512722 362960 512788 362994
rect 512822 362960 512888 362994
rect 512922 362960 512988 362994
rect 513022 362960 513088 362994
rect 513122 362960 513154 362994
rect 512542 362894 513154 362960
rect 512542 362860 512588 362894
rect 512622 362860 512688 362894
rect 512722 362860 512788 362894
rect 512822 362860 512888 362894
rect 512922 362860 512988 362894
rect 513022 362860 513088 362894
rect 513122 362860 513154 362894
rect 512542 362814 513154 362860
rect 513728 372798 513848 372953
rect 513728 372787 513780 372798
rect 513728 372753 513771 372787
rect 513728 372746 513780 372753
rect 513832 372746 513848 372798
rect 513728 372587 513848 372746
rect 513728 372553 513771 372587
rect 513805 372553 513848 372587
rect 513728 372387 513848 372553
rect 513728 372353 513771 372387
rect 513805 372353 513848 372387
rect 513728 372187 513848 372353
rect 513728 372153 513771 372187
rect 513805 372153 513848 372187
rect 513728 371987 513848 372153
rect 513728 371953 513771 371987
rect 513805 371953 513848 371987
rect 513728 371787 513848 371953
rect 513728 371753 513771 371787
rect 513805 371753 513848 371787
rect 513728 371587 513848 371753
rect 513728 371553 513771 371587
rect 513805 371553 513848 371587
rect 513728 371387 513848 371553
rect 513728 371353 513771 371387
rect 513805 371353 513848 371387
rect 513728 371187 513848 371353
rect 513728 371153 513771 371187
rect 513805 371153 513848 371187
rect 513728 370987 513848 371153
rect 513728 370953 513771 370987
rect 513805 370953 513848 370987
rect 513728 370787 513848 370953
rect 513728 370753 513771 370787
rect 513805 370753 513848 370787
rect 513728 370587 513848 370753
rect 513728 370553 513771 370587
rect 513805 370553 513848 370587
rect 513728 370387 513848 370553
rect 513728 370353 513771 370387
rect 513805 370353 513848 370387
rect 513728 370187 513848 370353
rect 513728 370153 513771 370187
rect 513805 370153 513848 370187
rect 513728 369987 513848 370153
rect 513728 369953 513771 369987
rect 513805 369953 513848 369987
rect 513728 369787 513848 369953
rect 513728 369753 513771 369787
rect 513805 369753 513848 369787
rect 513728 369587 513848 369753
rect 513728 369553 513771 369587
rect 513805 369553 513848 369587
rect 513728 369387 513848 369553
rect 513728 369353 513771 369387
rect 513805 369353 513848 369387
rect 513728 369187 513848 369353
rect 513728 369153 513771 369187
rect 513805 369153 513848 369187
rect 513728 368987 513848 369153
rect 513728 368953 513771 368987
rect 513805 368953 513848 368987
rect 513728 368787 513848 368953
rect 513728 368753 513771 368787
rect 513805 368753 513848 368787
rect 513728 368587 513848 368753
rect 513728 368553 513771 368587
rect 513805 368553 513848 368587
rect 513728 368387 513848 368553
rect 513728 368353 513771 368387
rect 513805 368353 513848 368387
rect 513728 368187 513848 368353
rect 513728 368153 513771 368187
rect 513805 368153 513848 368187
rect 513728 367987 513848 368153
rect 513728 367953 513771 367987
rect 513805 367953 513848 367987
rect 513728 367787 513848 367953
rect 513728 367753 513771 367787
rect 513805 367753 513848 367787
rect 513728 367587 513848 367753
rect 513728 367553 513771 367587
rect 513805 367553 513848 367587
rect 513728 367387 513848 367553
rect 513728 367353 513771 367387
rect 513805 367353 513848 367387
rect 513728 367187 513848 367353
rect 513728 367153 513771 367187
rect 513805 367153 513848 367187
rect 513728 366987 513848 367153
rect 513728 366953 513771 366987
rect 513805 366953 513848 366987
rect 513728 366787 513848 366953
rect 513728 366753 513771 366787
rect 513805 366753 513848 366787
rect 513728 366587 513848 366753
rect 513728 366553 513771 366587
rect 513805 366553 513848 366587
rect 513728 366387 513848 366553
rect 513728 366353 513771 366387
rect 513805 366353 513848 366387
rect 513728 366187 513848 366353
rect 513728 366153 513771 366187
rect 513805 366153 513848 366187
rect 513728 365987 513848 366153
rect 513728 365953 513771 365987
rect 513805 365953 513848 365987
rect 513728 365787 513848 365953
rect 513728 365753 513771 365787
rect 513805 365753 513848 365787
rect 513728 365587 513848 365753
rect 513728 365553 513771 365587
rect 513805 365553 513848 365587
rect 513728 365387 513848 365553
rect 513728 365353 513771 365387
rect 513805 365353 513848 365387
rect 513728 365187 513848 365353
rect 513728 365153 513771 365187
rect 513805 365153 513848 365187
rect 513728 364987 513848 365153
rect 513728 364953 513771 364987
rect 513805 364953 513848 364987
rect 513728 364787 513848 364953
rect 513728 364753 513771 364787
rect 513805 364753 513848 364787
rect 513728 364587 513848 364753
rect 513728 364553 513771 364587
rect 513805 364553 513848 364587
rect 513728 364387 513848 364553
rect 513728 364353 513771 364387
rect 513805 364353 513848 364387
rect 513728 364187 513848 364353
rect 513728 364153 513771 364187
rect 513805 364153 513848 364187
rect 513728 363987 513848 364153
rect 513728 363953 513771 363987
rect 513805 363953 513848 363987
rect 513728 363787 513848 363953
rect 513728 363753 513771 363787
rect 513805 363753 513848 363787
rect 513728 363587 513848 363753
rect 513728 363553 513771 363587
rect 513805 363553 513848 363587
rect 513728 363387 513848 363553
rect 513728 363353 513771 363387
rect 513805 363353 513848 363387
rect 513728 363187 513848 363353
rect 513728 363153 513771 363187
rect 513805 363153 513848 363187
rect 513728 362987 513848 363153
rect 513728 362953 513771 362987
rect 513805 362953 513848 362987
rect 512368 362736 512384 362770
rect 512418 362736 512438 362770
rect 512368 362680 512438 362736
rect 512368 362646 512384 362680
rect 512418 362646 512438 362680
rect 512368 362640 512438 362646
rect 513728 362787 513848 362953
rect 513728 362753 513771 362787
rect 513805 362753 513848 362787
rect 512218 362574 512288 362630
rect 512218 362540 512224 362574
rect 512258 362540 512288 362574
rect 512218 362476 512288 362540
rect 513728 362587 513848 362753
rect 513728 362553 513771 362587
rect 513805 362553 513848 362587
rect 511848 359888 511850 361476
rect 511966 359888 511968 361476
rect 511848 359866 511968 359888
rect 509968 357440 509970 359028
rect 510086 357440 510088 359028
rect 509968 357418 510088 357440
rect 513728 359028 513848 362553
rect 515608 411584 515728 411606
rect 515608 409996 515610 411584
rect 515726 409996 515728 411584
rect 515608 392371 515728 409996
rect 516160 401042 516212 401048
rect 516160 400984 516212 400990
rect 516172 392543 516200 400984
rect 515608 392337 515651 392371
rect 515685 392337 515728 392371
rect 515608 392171 515728 392337
rect 515608 392137 515651 392171
rect 515685 392137 515728 392171
rect 515608 391971 515728 392137
rect 515907 392535 516469 392543
rect 515907 392141 515919 392535
rect 516457 392141 516469 392535
rect 515907 392133 516469 392141
rect 516867 392535 517429 392543
rect 516867 392141 516879 392535
rect 517417 392141 517429 392535
rect 516867 392133 517429 392141
rect 517488 392371 517608 412444
rect 521248 414032 521368 414054
rect 521248 412444 521250 414032
rect 521366 412444 521368 414032
rect 517488 392337 517531 392371
rect 517565 392337 517608 392371
rect 517488 392171 517608 392337
rect 517488 392137 517531 392171
rect 517565 392137 517608 392171
rect 517396 392032 517424 392133
rect 515608 391937 515651 391971
rect 515685 391937 515728 391971
rect 517384 392026 517436 392032
rect 517384 391968 517436 391974
rect 517488 391971 517608 392137
rect 515608 391771 515728 391937
rect 515608 391737 515651 391771
rect 515685 391737 515728 391771
rect 515608 391571 515728 391737
rect 515608 391537 515651 391571
rect 515685 391537 515728 391571
rect 515608 391371 515728 391537
rect 515608 391337 515651 391371
rect 515685 391337 515728 391371
rect 515608 391171 515728 391337
rect 515608 391137 515651 391171
rect 515685 391137 515728 391171
rect 515608 390971 515728 391137
rect 515608 390937 515651 390971
rect 515685 390937 515728 390971
rect 515608 390771 515728 390937
rect 515608 390737 515651 390771
rect 515685 390737 515728 390771
rect 515608 390571 515728 390737
rect 515608 390537 515651 390571
rect 515685 390537 515728 390571
rect 517488 391937 517531 391971
rect 517565 391937 517608 391971
rect 517488 391771 517608 391937
rect 517488 391737 517531 391771
rect 517565 391737 517608 391771
rect 517488 391571 517608 391737
rect 517488 391537 517531 391571
rect 517565 391537 517608 391571
rect 517488 391371 517608 391537
rect 517488 391337 517531 391371
rect 517565 391337 517608 391371
rect 517488 391171 517608 391337
rect 517488 391137 517531 391171
rect 517565 391137 517608 391171
rect 517488 390971 517608 391137
rect 517488 390937 517531 390971
rect 517565 390937 517608 390971
rect 517488 390771 517608 390937
rect 517488 390737 517531 390771
rect 517565 390737 517608 390771
rect 517488 390571 517608 390737
rect 515608 390371 515728 390537
rect 516469 390535 517433 390546
rect 515608 390337 515651 390371
rect 515685 390337 515728 390371
rect 515608 389353 515728 390337
rect 515907 390528 517433 390535
rect 515907 390134 515919 390528
rect 516457 390134 516879 390528
rect 517417 390134 517433 390528
rect 515907 390125 517433 390134
rect 516469 390114 517433 390125
rect 517488 390537 517531 390571
rect 517565 390537 517608 390571
rect 517488 390371 517608 390537
rect 517488 390337 517531 390371
rect 517565 390337 517608 390371
rect 516908 389542 516960 389548
rect 516148 389524 516908 389530
rect 516148 389490 516171 389524
rect 516205 389490 516243 389524
rect 516277 389490 516315 389524
rect 516349 389490 516387 389524
rect 516421 389490 516459 389524
rect 516493 389490 516531 389524
rect 516565 389490 516603 389524
rect 516637 389490 516675 389524
rect 516709 389490 516747 389524
rect 516781 389490 516819 389524
rect 516853 389490 516891 389524
rect 516148 389484 516960 389490
rect 515608 389319 515651 389353
rect 515685 389319 515728 389353
rect 515608 388953 515728 389319
rect 517488 389353 517608 390337
rect 517488 389319 517531 389353
rect 517565 389319 517608 389353
rect 516148 389070 516948 389072
rect 517488 389070 517608 389319
rect 516148 389066 517608 389070
rect 516148 389032 516171 389066
rect 516205 389032 516243 389066
rect 516277 389032 516315 389066
rect 516349 389032 516387 389066
rect 516421 389032 516459 389066
rect 516493 389032 516531 389066
rect 516565 389032 516603 389066
rect 516637 389032 516675 389066
rect 516709 389032 516747 389066
rect 516781 389032 516819 389066
rect 516853 389032 516891 389066
rect 516925 389042 517608 389066
rect 516925 389032 516948 389042
rect 516148 389026 516948 389032
rect 515608 388919 515651 388953
rect 515685 388919 515728 388953
rect 515608 388553 515728 388919
rect 517488 388953 517608 389042
rect 517488 388919 517531 388953
rect 517565 388919 517608 388953
rect 516148 388608 516948 388614
rect 516148 388574 516171 388608
rect 516205 388574 516243 388608
rect 516277 388574 516315 388608
rect 516349 388574 516387 388608
rect 516421 388574 516459 388608
rect 516493 388574 516531 388608
rect 516565 388574 516603 388608
rect 516637 388574 516675 388608
rect 516709 388574 516747 388608
rect 516781 388574 516819 388608
rect 516853 388574 516891 388608
rect 516925 388574 516948 388608
rect 516148 388568 516948 388574
rect 515608 388519 515651 388553
rect 515685 388519 515728 388553
rect 515608 388153 515728 388519
rect 517488 388553 517608 388919
rect 517488 388519 517531 388553
rect 517565 388519 517608 388553
rect 515608 388119 515651 388153
rect 515685 388119 515728 388153
rect 515608 387753 515728 388119
rect 516148 388150 516948 388156
rect 516148 388116 516171 388150
rect 516205 388116 516243 388150
rect 516277 388116 516315 388150
rect 516349 388116 516387 388150
rect 516421 388116 516459 388150
rect 516493 388116 516531 388150
rect 516565 388116 516603 388150
rect 516637 388116 516675 388150
rect 516709 388116 516747 388150
rect 516781 388116 516819 388150
rect 516853 388116 516891 388150
rect 516925 388116 516948 388150
rect 516148 388110 516948 388116
rect 517488 388153 517608 388519
rect 517488 388119 517531 388153
rect 517565 388119 517608 388153
rect 515608 387719 515651 387753
rect 515685 387719 515728 387753
rect 515608 387353 515728 387719
rect 517488 387753 517608 388119
rect 517488 387719 517531 387753
rect 517565 387719 517608 387753
rect 516148 387692 516948 387698
rect 516148 387658 516171 387692
rect 516205 387658 516243 387692
rect 516277 387658 516315 387692
rect 516349 387658 516387 387692
rect 516421 387658 516459 387692
rect 516493 387658 516531 387692
rect 516565 387658 516603 387692
rect 516637 387658 516675 387692
rect 516709 387658 516747 387692
rect 516781 387658 516819 387692
rect 516853 387658 516891 387692
rect 516925 387658 516948 387692
rect 516148 387652 516948 387658
rect 517192 387432 517220 387487
rect 517180 387426 517232 387432
rect 517180 387368 517232 387374
rect 515608 387319 515651 387353
rect 515685 387319 515728 387353
rect 515608 386953 515728 387319
rect 517488 387353 517608 387719
rect 517488 387319 517531 387353
rect 517565 387319 517608 387353
rect 516148 387234 516948 387240
rect 516148 387200 516171 387234
rect 516205 387200 516243 387234
rect 516277 387200 516315 387234
rect 516349 387200 516387 387234
rect 516421 387200 516459 387234
rect 516493 387200 516531 387234
rect 516565 387200 516603 387234
rect 516637 387200 516675 387234
rect 516709 387200 516747 387234
rect 516781 387200 516819 387234
rect 516853 387200 516891 387234
rect 516925 387200 516948 387234
rect 516148 387194 516948 387200
rect 515608 386919 515651 386953
rect 515685 386919 515728 386953
rect 515608 386553 515728 386919
rect 517488 386953 517608 387319
rect 517488 386919 517531 386953
rect 517565 386919 517608 386953
rect 516148 386776 516948 386782
rect 516148 386742 516171 386776
rect 516205 386742 516243 386776
rect 516277 386742 516315 386776
rect 516349 386742 516387 386776
rect 516421 386742 516459 386776
rect 516493 386742 516531 386776
rect 516565 386742 516603 386776
rect 516637 386742 516675 386776
rect 516709 386742 516747 386776
rect 516781 386742 516819 386776
rect 516853 386742 516891 386776
rect 516925 386742 516948 386776
rect 516148 386736 516948 386742
rect 515608 386519 515651 386553
rect 515685 386519 515728 386553
rect 515608 386153 515728 386519
rect 517488 386553 517608 386919
rect 517488 386519 517531 386553
rect 517565 386519 517608 386553
rect 516148 386318 516948 386324
rect 516148 386284 516171 386318
rect 516205 386284 516243 386318
rect 516277 386284 516315 386318
rect 516349 386284 516387 386318
rect 516421 386284 516459 386318
rect 516493 386284 516531 386318
rect 516565 386284 516603 386318
rect 516637 386284 516675 386318
rect 516709 386284 516747 386318
rect 516781 386284 516819 386318
rect 516853 386284 516891 386318
rect 516925 386284 516948 386318
rect 516148 386278 516948 386284
rect 515608 386119 515651 386153
rect 515685 386119 515728 386153
rect 515608 385753 515728 386119
rect 517488 386153 517608 386519
rect 517488 386119 517531 386153
rect 517565 386119 517608 386153
rect 516148 385860 516948 385866
rect 516148 385826 516171 385860
rect 516205 385826 516243 385860
rect 516277 385826 516315 385860
rect 516349 385826 516387 385860
rect 516421 385826 516459 385860
rect 516493 385826 516531 385860
rect 516565 385826 516603 385860
rect 516637 385826 516675 385860
rect 516709 385826 516747 385860
rect 516781 385826 516819 385860
rect 516853 385826 516891 385860
rect 516925 385826 516948 385860
rect 516148 385820 516948 385826
rect 515608 385719 515651 385753
rect 515685 385719 515728 385753
rect 515608 384843 515728 385719
rect 516308 385500 516336 385820
rect 517488 385753 517608 386119
rect 517488 385719 517531 385753
rect 517565 385719 517608 385753
rect 516296 385494 516348 385500
rect 516296 385436 516348 385442
rect 516148 385402 516948 385408
rect 516148 385368 516171 385402
rect 516205 385368 516243 385402
rect 516277 385368 516315 385402
rect 516349 385368 516387 385402
rect 516421 385368 516459 385402
rect 516493 385368 516531 385402
rect 516565 385368 516603 385402
rect 516637 385368 516675 385402
rect 516709 385368 516747 385402
rect 516781 385368 516819 385402
rect 516853 385368 516891 385402
rect 516925 385368 516948 385402
rect 516148 385362 516948 385368
rect 515608 384809 515651 384843
rect 515685 384809 515728 384843
rect 515608 384443 515728 384809
rect 515608 384409 515651 384443
rect 515685 384409 515728 384443
rect 515608 384043 515728 384409
rect 515608 384009 515651 384043
rect 515685 384009 515728 384043
rect 515608 383643 515728 384009
rect 515608 383609 515651 383643
rect 515685 383609 515728 383643
rect 515608 383243 515728 383609
rect 515608 383209 515651 383243
rect 515685 383209 515728 383243
rect 515608 382843 515728 383209
rect 515608 382809 515651 382843
rect 515685 382809 515728 382843
rect 515608 382443 515728 382809
rect 515608 382409 515651 382443
rect 515685 382409 515728 382443
rect 515608 382043 515728 382409
rect 515608 382009 515651 382043
rect 515685 382009 515728 382043
rect 515608 381643 515728 382009
rect 515608 381609 515651 381643
rect 515685 381609 515728 381643
rect 515608 381538 515728 381609
rect 515608 381486 515616 381538
rect 515668 381486 515728 381538
rect 515608 381243 515728 381486
rect 515608 381209 515651 381243
rect 515685 381209 515728 381243
rect 515608 380843 515728 381209
rect 515608 380809 515651 380843
rect 515685 380809 515728 380843
rect 515608 380443 515728 380809
rect 515608 380409 515651 380443
rect 515685 380409 515728 380443
rect 515608 380043 515728 380409
rect 515608 380009 515651 380043
rect 515685 380009 515728 380043
rect 515608 379643 515728 380009
rect 515608 379609 515651 379643
rect 515685 379609 515728 379643
rect 515608 379243 515728 379609
rect 515608 379209 515651 379243
rect 515685 379209 515728 379243
rect 515608 378843 515728 379209
rect 515608 378809 515651 378843
rect 515685 378809 515728 378843
rect 515608 378443 515728 378809
rect 515608 378409 515651 378443
rect 515685 378409 515728 378443
rect 515608 378043 515728 378409
rect 515608 378009 515651 378043
rect 515685 378009 515728 378043
rect 515608 377377 515728 378009
rect 517488 384843 517608 385719
rect 517488 384809 517531 384843
rect 517565 384809 517608 384843
rect 517488 384443 517608 384809
rect 517488 384409 517531 384443
rect 517565 384409 517608 384443
rect 517488 384043 517608 384409
rect 517488 384009 517531 384043
rect 517565 384009 517608 384043
rect 519368 411584 519488 411606
rect 519368 409996 519370 411584
rect 519486 409996 519488 411584
rect 519368 390901 519488 409996
rect 520648 398282 520700 398288
rect 520648 398224 520700 398230
rect 519696 392026 519748 392032
rect 519696 391968 519748 391974
rect 519708 391073 519736 391968
rect 520660 391073 520688 398224
rect 519368 390867 519411 390901
rect 519445 390867 519488 390901
rect 519368 390701 519488 390867
rect 519368 390667 519411 390701
rect 519445 390667 519488 390701
rect 519368 390501 519488 390667
rect 519667 391065 520229 391073
rect 519667 390671 519679 391065
rect 520217 390671 520229 391065
rect 519667 390663 520229 390671
rect 520627 391065 521189 391073
rect 520627 390671 520639 391065
rect 521177 390671 521189 391065
rect 520627 390663 521189 390671
rect 521248 390901 521368 412444
rect 525008 414032 525128 414054
rect 525008 412444 525010 414032
rect 525126 412444 525128 414032
rect 521248 390867 521291 390901
rect 521325 390867 521368 390901
rect 521248 390701 521368 390867
rect 521248 390667 521291 390701
rect 521325 390667 521368 390701
rect 519368 390467 519411 390501
rect 519445 390467 519488 390501
rect 519368 390301 519488 390467
rect 519368 390267 519411 390301
rect 519445 390267 519488 390301
rect 519368 390101 519488 390267
rect 519368 390067 519411 390101
rect 519445 390067 519488 390101
rect 519368 389901 519488 390067
rect 519368 389867 519411 389901
rect 519445 389867 519488 389901
rect 519368 389701 519488 389867
rect 519368 389667 519411 389701
rect 519445 389667 519488 389701
rect 519368 389501 519488 389667
rect 519368 389467 519411 389501
rect 519445 389467 519488 389501
rect 519368 389301 519488 389467
rect 519368 389267 519411 389301
rect 519445 389267 519488 389301
rect 519368 389101 519488 389267
rect 519368 389067 519411 389101
rect 519445 389067 519488 389101
rect 521248 390501 521368 390667
rect 521248 390467 521291 390501
rect 521325 390467 521368 390501
rect 521248 390301 521368 390467
rect 521248 390267 521291 390301
rect 521325 390267 521368 390301
rect 521248 390101 521368 390267
rect 521248 390067 521291 390101
rect 521325 390067 521368 390101
rect 521248 389901 521368 390067
rect 521248 389867 521291 389901
rect 521325 389867 521368 389901
rect 521248 389701 521368 389867
rect 521248 389667 521291 389701
rect 521325 389667 521368 389701
rect 521248 389501 521368 389667
rect 521248 389467 521291 389501
rect 521325 389467 521368 389501
rect 521248 389301 521368 389467
rect 521248 389267 521291 389301
rect 521325 389267 521368 389301
rect 521248 389101 521368 389267
rect 519368 388901 519488 389067
rect 520229 389065 521193 389076
rect 519368 388867 519411 388901
rect 519445 388867 519488 388901
rect 519368 387569 519488 388867
rect 519667 389058 521193 389065
rect 519667 388664 519679 389058
rect 520217 388664 520639 389058
rect 521177 388664 521193 389058
rect 519667 388655 521193 388664
rect 520229 388644 521193 388655
rect 521248 389067 521291 389101
rect 521325 389067 521368 389101
rect 521248 388901 521368 389067
rect 521248 388867 521291 388901
rect 521325 388867 521368 388901
rect 519368 387535 519411 387569
rect 519445 387535 519488 387569
rect 519368 387369 519488 387535
rect 519368 387335 519411 387369
rect 519445 387335 519488 387369
rect 519368 387169 519488 387335
rect 519667 387733 520229 387741
rect 519667 387339 519679 387733
rect 520217 387339 520229 387733
rect 519667 387331 520229 387339
rect 520627 387733 521189 387741
rect 520627 387339 520639 387733
rect 521177 387339 521189 387733
rect 520627 387331 521189 387339
rect 521248 387569 521368 388867
rect 521248 387535 521291 387569
rect 521325 387535 521368 387569
rect 521248 387369 521368 387535
rect 521248 387335 521291 387369
rect 521325 387335 521368 387369
rect 519368 387135 519411 387169
rect 519445 387135 519488 387169
rect 519368 386969 519488 387135
rect 519368 386935 519411 386969
rect 519445 386935 519488 386969
rect 519368 386769 519488 386935
rect 519368 386735 519411 386769
rect 519445 386735 519488 386769
rect 519368 386569 519488 386735
rect 519368 386535 519411 386569
rect 519445 386535 519488 386569
rect 519368 386369 519488 386535
rect 519368 386335 519411 386369
rect 519445 386335 519488 386369
rect 519368 386169 519488 386335
rect 519368 386135 519411 386169
rect 519445 386135 519488 386169
rect 519368 385969 519488 386135
rect 519368 385935 519411 385969
rect 519445 385935 519488 385969
rect 519368 385769 519488 385935
rect 520184 385868 520212 387331
rect 521248 387169 521368 387335
rect 521248 387135 521291 387169
rect 521325 387135 521368 387169
rect 521248 386969 521368 387135
rect 521248 386935 521291 386969
rect 521325 386935 521368 386969
rect 521248 386769 521368 386935
rect 521248 386735 521291 386769
rect 521325 386735 521368 386769
rect 521248 386569 521368 386735
rect 521248 386535 521291 386569
rect 521325 386535 521368 386569
rect 521248 386369 521368 386535
rect 521248 386335 521291 386369
rect 521325 386335 521368 386369
rect 521248 386169 521368 386335
rect 521248 386135 521291 386169
rect 521325 386135 521368 386169
rect 521248 385969 521368 386135
rect 521248 385935 521291 385969
rect 521325 385935 521368 385969
rect 520172 385862 520224 385868
rect 520172 385804 520224 385810
rect 519368 385735 519411 385769
rect 519445 385735 519488 385769
rect 521248 385769 521368 385935
rect 519368 385569 519488 385735
rect 520229 385733 521193 385744
rect 519368 385535 519411 385569
rect 519445 385535 519488 385569
rect 519368 384825 519488 385535
rect 519667 385726 521193 385733
rect 519667 385332 519679 385726
rect 520217 385332 520639 385726
rect 521177 385332 521193 385726
rect 519667 385323 521193 385332
rect 520229 385312 521193 385323
rect 521248 385735 521291 385769
rect 521325 385735 521368 385769
rect 521248 385569 521368 385735
rect 521248 385535 521291 385569
rect 521325 385535 521368 385569
rect 520648 385218 520700 385224
rect 520648 385160 520700 385166
rect 520660 384997 520688 385160
rect 519368 384791 519411 384825
rect 519445 384791 519488 384825
rect 519368 384625 519488 384791
rect 519368 384591 519411 384625
rect 519445 384591 519488 384625
rect 519368 384425 519488 384591
rect 519667 384989 520229 384997
rect 519667 384595 519679 384989
rect 520217 384595 520229 384989
rect 519667 384587 520229 384595
rect 520627 384989 521189 384997
rect 520627 384595 520639 384989
rect 521177 384595 521189 384989
rect 520627 384587 521189 384595
rect 521248 384825 521368 385535
rect 521248 384791 521291 384825
rect 521325 384791 521368 384825
rect 521248 384625 521368 384791
rect 521248 384591 521291 384625
rect 521325 384591 521368 384625
rect 519368 384391 519411 384425
rect 519445 384391 519488 384425
rect 519368 384225 519488 384391
rect 519368 384191 519411 384225
rect 519445 384191 519488 384225
rect 517488 383643 517608 384009
rect 518608 384022 518660 384028
rect 518608 383964 518660 383970
rect 519368 384025 519488 384191
rect 519708 384028 519736 384587
rect 521248 384425 521368 384591
rect 521248 384391 521291 384425
rect 521325 384391 521368 384425
rect 521248 384225 521368 384391
rect 521248 384191 521291 384225
rect 521325 384191 521368 384225
rect 519368 383991 519411 384025
rect 519445 383991 519488 384025
rect 517488 383609 517531 383643
rect 517565 383609 517608 383643
rect 517488 383243 517608 383609
rect 517488 383209 517531 383243
rect 517565 383209 517608 383243
rect 517488 382843 517608 383209
rect 517488 382809 517531 382843
rect 517565 382809 517608 382843
rect 517488 382443 517608 382809
rect 517488 382409 517531 382443
rect 517565 382409 517608 382443
rect 517488 382043 517608 382409
rect 517488 382009 517531 382043
rect 517565 382009 517608 382043
rect 517488 381643 517608 382009
rect 517488 381609 517531 381643
rect 517565 381609 517608 381643
rect 517488 381243 517608 381609
rect 517488 381209 517531 381243
rect 517565 381209 517608 381243
rect 517488 380843 517608 381209
rect 517488 380809 517531 380843
rect 517565 380809 517608 380843
rect 517488 380443 517608 380809
rect 517488 380409 517531 380443
rect 517565 380409 517608 380443
rect 517488 380043 517608 380409
rect 517488 380009 517531 380043
rect 517565 380009 517608 380043
rect 517488 379643 517608 380009
rect 517488 379609 517531 379643
rect 517565 379609 517608 379643
rect 517488 379243 517608 379609
rect 517488 379209 517531 379243
rect 517565 379209 517608 379243
rect 517488 378843 517608 379209
rect 517488 378809 517531 378843
rect 517565 378809 517608 378843
rect 517488 378443 517608 378809
rect 517488 378409 517531 378443
rect 517565 378409 517608 378443
rect 517488 378043 517608 378409
rect 517488 378009 517531 378043
rect 517565 378009 517608 378043
rect 517384 377582 517436 377588
rect 515608 377343 515651 377377
rect 515685 377343 515728 377377
rect 515608 377177 515728 377343
rect 515907 377541 516469 377549
rect 515907 377202 515919 377541
rect 515608 377143 515651 377177
rect 515685 377143 515728 377177
rect 515608 376977 515728 377143
rect 515608 376943 515651 376977
rect 515685 376943 515728 376977
rect 515608 376777 515728 376943
rect 515608 376743 515651 376777
rect 515685 376743 515728 376777
rect 515608 376577 515728 376743
rect 515608 376543 515651 376577
rect 515685 376543 515728 376577
rect 515608 376377 515728 376543
rect 515608 376343 515651 376377
rect 515685 376343 515728 376377
rect 515608 376177 515728 376343
rect 515608 376143 515651 376177
rect 515685 376143 515728 376177
rect 515608 375977 515728 376143
rect 515608 375943 515651 375977
rect 515685 375943 515728 375977
rect 515608 375777 515728 375943
rect 515608 375743 515651 375777
rect 515685 375743 515728 375777
rect 515608 375577 515728 375743
rect 515608 375543 515651 375577
rect 515685 375543 515728 375577
rect 515608 375377 515728 375543
rect 515608 375343 515651 375377
rect 515685 375343 515728 375377
rect 515608 374633 515728 375343
rect 515832 377174 515919 377202
rect 515832 375012 515860 377174
rect 515907 377147 515919 377174
rect 516457 377147 516469 377541
rect 515907 377139 516469 377147
rect 516867 377541 517384 377549
rect 516867 377147 516879 377541
rect 517417 377524 517436 377530
rect 517417 377147 517429 377524
rect 516867 377139 517429 377147
rect 517488 377377 517608 378009
rect 518620 377588 518648 383964
rect 519368 383825 519488 383991
rect 519696 384022 519748 384028
rect 519696 383964 519748 383970
rect 521248 384025 521368 384191
rect 521248 383991 521291 384025
rect 521325 383991 521368 384025
rect 519368 383791 519411 383825
rect 519445 383791 519488 383825
rect 519368 383625 519488 383791
rect 519368 383591 519411 383625
rect 519445 383591 519488 383625
rect 519368 383425 519488 383591
rect 519368 383391 519411 383425
rect 519445 383391 519488 383425
rect 519368 383225 519488 383391
rect 519368 383191 519411 383225
rect 519445 383191 519488 383225
rect 519368 383025 519488 383191
rect 519368 382991 519411 383025
rect 519445 382991 519488 383025
rect 521248 383825 521368 383991
rect 521248 383791 521291 383825
rect 521325 383791 521368 383825
rect 521248 383625 521368 383791
rect 521248 383591 521291 383625
rect 521325 383591 521368 383625
rect 521248 383425 521368 383591
rect 521248 383391 521291 383425
rect 521325 383391 521368 383425
rect 521248 383225 521368 383391
rect 521248 383191 521291 383225
rect 521325 383191 521368 383225
rect 521248 383025 521368 383191
rect 519368 382825 519488 382991
rect 520229 382989 521193 383000
rect 519368 382791 519411 382825
rect 519445 382791 519488 382825
rect 519368 381591 519488 382791
rect 519667 382982 521193 382989
rect 519667 382588 519679 382982
rect 520217 382588 520639 382982
rect 521177 382588 521193 382982
rect 519667 382579 521193 382588
rect 520229 382568 521193 382579
rect 521248 382991 521291 383025
rect 521325 382991 521368 383025
rect 521248 382825 521368 382991
rect 521248 382791 521291 382825
rect 521325 382791 521368 382825
rect 519368 381557 519411 381591
rect 519445 381557 519488 381591
rect 519368 381391 519488 381557
rect 519368 381357 519411 381391
rect 519445 381357 519488 381391
rect 519368 381191 519488 381357
rect 519667 381755 520229 381763
rect 519667 381361 519679 381755
rect 520217 381361 520229 381755
rect 519667 381353 520229 381361
rect 520627 381755 521189 381763
rect 520627 381361 520639 381755
rect 521177 381361 521189 381755
rect 520627 381353 521189 381361
rect 521248 381591 521368 382791
rect 521248 381557 521291 381591
rect 521325 381557 521368 381591
rect 521248 381391 521368 381557
rect 521248 381357 521291 381391
rect 521325 381357 521368 381391
rect 519368 381157 519411 381191
rect 519445 381157 519488 381191
rect 519368 380991 519488 381157
rect 519368 380957 519411 380991
rect 519445 380957 519488 380991
rect 519368 380791 519488 380957
rect 519368 380757 519411 380791
rect 519445 380757 519488 380791
rect 519368 380591 519488 380757
rect 519368 380557 519411 380591
rect 519445 380557 519488 380591
rect 519368 380391 519488 380557
rect 519368 380357 519411 380391
rect 519445 380357 519488 380391
rect 519368 380191 519488 380357
rect 519368 380157 519411 380191
rect 519445 380157 519488 380191
rect 519368 379991 519488 380157
rect 519368 379957 519411 379991
rect 519445 379957 519488 379991
rect 519368 379791 519488 379957
rect 519560 379974 519612 379980
rect 519560 379916 519612 379922
rect 519368 379757 519411 379791
rect 519445 379757 519488 379791
rect 519368 379591 519488 379757
rect 519368 379557 519411 379591
rect 519445 379557 519488 379591
rect 518608 377582 518660 377588
rect 518608 377524 518660 377530
rect 517488 377343 517531 377377
rect 517565 377343 517608 377377
rect 517488 377177 517608 377343
rect 517488 377143 517531 377177
rect 517565 377143 517608 377177
rect 517488 376977 517608 377143
rect 517488 376943 517531 376977
rect 517565 376943 517608 376977
rect 517488 376777 517608 376943
rect 517488 376743 517531 376777
rect 517565 376743 517608 376777
rect 517488 376577 517608 376743
rect 519368 377377 519488 379557
rect 519368 377343 519411 377377
rect 519445 377343 519488 377377
rect 519368 377177 519488 377343
rect 519368 377143 519411 377177
rect 519445 377143 519488 377177
rect 519368 376977 519488 377143
rect 519368 376943 519411 376977
rect 519445 376943 519488 376977
rect 519368 376777 519488 376943
rect 519368 376743 519411 376777
rect 519445 376743 519488 376777
rect 517860 376662 517912 376668
rect 517860 376604 517912 376610
rect 517488 376543 517531 376577
rect 517565 376543 517608 376577
rect 517488 376377 517608 376543
rect 517488 376343 517531 376377
rect 517565 376343 517608 376377
rect 517488 376177 517608 376343
rect 517488 376143 517531 376177
rect 517565 376143 517608 376177
rect 517488 375977 517608 376143
rect 517488 375943 517531 375977
rect 517565 375943 517608 375977
rect 517488 375777 517608 375943
rect 517488 375743 517531 375777
rect 517565 375743 517608 375777
rect 517488 375577 517608 375743
rect 516469 375541 517433 375552
rect 515907 375534 517433 375541
rect 515907 375140 515919 375534
rect 516457 375140 516879 375534
rect 517417 375140 517433 375534
rect 515907 375131 517433 375140
rect 516469 375120 517433 375131
rect 517488 375543 517531 375577
rect 517565 375543 517608 375577
rect 517488 375377 517608 375543
rect 517488 375343 517531 375377
rect 517565 375343 517608 375377
rect 515820 375006 515872 375012
rect 515820 374948 515872 374954
rect 516908 375006 516960 375012
rect 516908 374948 516960 374954
rect 516432 374822 516484 374828
rect 515608 374599 515651 374633
rect 515685 374599 515728 374633
rect 515608 374433 515728 374599
rect 515608 374399 515651 374433
rect 515685 374399 515728 374433
rect 515608 374233 515728 374399
rect 515907 374797 516432 374805
rect 516920 374805 516948 374948
rect 515907 374403 515919 374797
rect 516457 374764 516484 374770
rect 516867 374797 517429 374805
rect 516457 374403 516469 374764
rect 515907 374395 516469 374403
rect 516867 374403 516879 374797
rect 517417 374403 517429 374797
rect 516867 374395 517429 374403
rect 517488 374633 517608 375343
rect 517488 374599 517531 374633
rect 517565 374599 517608 374633
rect 517488 374433 517608 374599
rect 517488 374399 517531 374433
rect 517565 374399 517608 374433
rect 515608 374199 515651 374233
rect 515685 374199 515728 374233
rect 515608 374033 515728 374199
rect 515608 373999 515651 374033
rect 515685 373999 515728 374033
rect 515608 373833 515728 373999
rect 515608 373799 515651 373833
rect 515685 373799 515728 373833
rect 515608 373633 515728 373799
rect 515608 373599 515651 373633
rect 515685 373599 515728 373633
rect 515608 373433 515728 373599
rect 517488 374233 517608 374399
rect 517488 374199 517531 374233
rect 517565 374199 517608 374233
rect 517488 374033 517608 374199
rect 517488 373999 517531 374033
rect 517565 373999 517608 374033
rect 517488 373833 517608 373999
rect 517488 373799 517531 373833
rect 517565 373799 517608 373833
rect 517488 373633 517608 373799
rect 517488 373599 517531 373633
rect 517565 373599 517608 373633
rect 515888 373534 515940 373540
rect 515608 373399 515651 373433
rect 515685 373399 515728 373433
rect 515608 373233 515728 373399
rect 515608 373199 515651 373233
rect 515685 373199 515728 373233
rect 515608 373033 515728 373199
rect 515608 372999 515651 373033
rect 515685 372999 515728 373033
rect 515608 372833 515728 372999
rect 515608 372799 515651 372833
rect 515685 372799 515728 372833
rect 515608 372633 515728 372799
rect 515608 372599 515651 372633
rect 515685 372599 515728 372633
rect 515608 371889 515728 372599
rect 515608 371855 515651 371889
rect 515685 371855 515728 371889
rect 515608 371689 515728 371855
rect 515608 371655 515651 371689
rect 515685 371655 515728 371689
rect 515608 371489 515728 371655
rect 515608 371455 515651 371489
rect 515685 371455 515728 371489
rect 515608 371289 515728 371455
rect 515608 371255 515651 371289
rect 515685 371255 515728 371289
rect 515608 371089 515728 371255
rect 515608 371055 515651 371089
rect 515685 371055 515728 371089
rect 515608 370889 515728 371055
rect 515608 370855 515651 370889
rect 515685 370855 515728 370889
rect 515608 370689 515728 370855
rect 515608 370655 515651 370689
rect 515685 370655 515728 370689
rect 515608 370489 515728 370655
rect 515608 370455 515651 370489
rect 515685 370455 515728 370489
rect 515608 370289 515728 370455
rect 515608 370255 515651 370289
rect 515685 370255 515728 370289
rect 515608 370089 515728 370255
rect 515608 370055 515651 370089
rect 515685 370055 515728 370089
rect 515608 369889 515728 370055
rect 515608 369855 515651 369889
rect 515685 369855 515728 369889
rect 515608 369145 515728 369855
rect 515832 373494 515888 373522
rect 515832 369290 515860 373494
rect 515888 373476 515940 373482
rect 517488 373433 517608 373599
rect 517488 373399 517531 373433
rect 517565 373399 517608 373433
rect 517488 373233 517608 373399
rect 517488 373199 517531 373233
rect 517565 373199 517608 373233
rect 517488 373033 517608 373199
rect 517488 372999 517531 373033
rect 517565 372999 517608 373033
rect 517488 372833 517608 372999
rect 516469 372797 517433 372808
rect 515907 372790 517433 372797
rect 515907 372396 515919 372790
rect 516457 372396 516879 372790
rect 517417 372396 517433 372790
rect 515907 372387 517433 372396
rect 516469 372376 517433 372387
rect 517488 372799 517531 372833
rect 517565 372799 517608 372833
rect 517488 372633 517608 372799
rect 517488 372599 517531 372633
rect 517565 372599 517608 372633
rect 516364 372246 516416 372252
rect 516364 372188 516416 372194
rect 516376 372061 516404 372188
rect 517384 372062 517436 372068
rect 515907 372053 516469 372061
rect 515907 371659 515919 372053
rect 516457 371659 516469 372053
rect 515907 371651 516469 371659
rect 516867 372053 517384 372061
rect 516867 371659 516879 372053
rect 517417 372004 517436 372010
rect 517417 371659 517429 372004
rect 516867 371651 517429 371659
rect 517488 371889 517608 372599
rect 517872 372068 517900 376604
rect 519368 376577 519488 376743
rect 519368 376543 519411 376577
rect 519445 376543 519488 376577
rect 519368 376377 519488 376543
rect 519368 376343 519411 376377
rect 519445 376343 519488 376377
rect 519368 376177 519488 376343
rect 519368 376143 519411 376177
rect 519445 376143 519488 376177
rect 519368 375977 519488 376143
rect 519368 375943 519411 375977
rect 519445 375943 519488 375977
rect 519368 375777 519488 375943
rect 519368 375743 519411 375777
rect 519445 375743 519488 375777
rect 519368 375577 519488 375743
rect 519368 375543 519411 375577
rect 519445 375543 519488 375577
rect 519368 375377 519488 375543
rect 519368 375343 519411 375377
rect 519445 375343 519488 375377
rect 519368 374633 519488 375343
rect 519572 374828 519600 379916
rect 520184 379888 520212 381353
rect 520660 379980 520688 381353
rect 521248 381191 521368 381357
rect 521248 381157 521291 381191
rect 521325 381157 521368 381191
rect 521248 380991 521368 381157
rect 521248 380957 521291 380991
rect 521325 380957 521368 380991
rect 521248 380791 521368 380957
rect 521248 380757 521291 380791
rect 521325 380757 521368 380791
rect 521248 380591 521368 380757
rect 521248 380557 521291 380591
rect 521325 380557 521368 380591
rect 521248 380391 521368 380557
rect 521248 380357 521291 380391
rect 521325 380357 521368 380391
rect 521248 380191 521368 380357
rect 521248 380157 521291 380191
rect 521325 380157 521368 380191
rect 521248 379991 521368 380157
rect 520648 379974 520700 379980
rect 520648 379916 520700 379922
rect 521248 379957 521291 379991
rect 521325 379957 521368 379991
rect 520172 379882 520224 379888
rect 520172 379824 520224 379830
rect 521248 379791 521368 379957
rect 520229 379755 521193 379766
rect 519667 379748 521193 379755
rect 519667 379354 519679 379748
rect 520217 379354 520639 379748
rect 521177 379354 521193 379748
rect 519667 379345 521193 379354
rect 520229 379334 521193 379345
rect 521248 379757 521291 379791
rect 521325 379757 521368 379791
rect 521248 379591 521368 379757
rect 521248 379557 521291 379591
rect 521325 379557 521368 379591
rect 520648 379238 520700 379244
rect 520648 379180 520700 379186
rect 520660 377549 520688 379180
rect 519667 377541 520229 377549
rect 519667 377147 519679 377541
rect 520217 377147 520229 377541
rect 519667 377139 520229 377147
rect 520627 377541 521189 377549
rect 520627 377147 520639 377541
rect 521177 377147 521189 377541
rect 520627 377139 521189 377147
rect 521248 377377 521368 379557
rect 521248 377343 521291 377377
rect 521325 377343 521368 377377
rect 521248 377177 521368 377343
rect 521248 377143 521291 377177
rect 521325 377143 521368 377177
rect 519708 376668 519736 377139
rect 521248 376977 521368 377143
rect 521248 376943 521291 376977
rect 521325 376943 521368 376977
rect 521248 376777 521368 376943
rect 521248 376743 521291 376777
rect 521325 376743 521368 376777
rect 519696 376662 519748 376668
rect 519696 376604 519748 376610
rect 521248 376577 521368 376743
rect 521248 376543 521291 376577
rect 521325 376543 521368 376577
rect 521248 376377 521368 376543
rect 521248 376343 521291 376377
rect 521325 376343 521368 376377
rect 521248 376177 521368 376343
rect 521248 376143 521291 376177
rect 521325 376143 521368 376177
rect 521248 375977 521368 376143
rect 521248 375943 521291 375977
rect 521325 375943 521368 375977
rect 521248 375777 521368 375943
rect 521248 375743 521291 375777
rect 521325 375743 521368 375777
rect 521248 375577 521368 375743
rect 520229 375541 521193 375552
rect 519667 375534 521193 375541
rect 519667 375140 519679 375534
rect 520217 375140 520639 375534
rect 521177 375140 521193 375534
rect 519667 375131 521193 375140
rect 520229 375120 521193 375131
rect 521248 375543 521291 375577
rect 521325 375543 521368 375577
rect 521248 375377 521368 375543
rect 521248 375343 521291 375377
rect 521325 375343 521368 375377
rect 519560 374822 519612 374828
rect 519560 374764 519612 374770
rect 519667 374797 520229 374805
rect 519368 374599 519411 374633
rect 519445 374599 519488 374633
rect 519368 374433 519488 374599
rect 519667 374442 519679 374797
rect 519368 374399 519411 374433
rect 519445 374399 519488 374433
rect 519368 374233 519488 374399
rect 519368 374199 519411 374233
rect 519445 374199 519488 374233
rect 519368 374033 519488 374199
rect 519368 373999 519411 374033
rect 519445 373999 519488 374033
rect 519368 373833 519488 373999
rect 519368 373799 519411 373833
rect 519445 373799 519488 373833
rect 519368 373633 519488 373799
rect 519368 373599 519411 373633
rect 519445 373599 519488 373633
rect 519368 373433 519488 373599
rect 519368 373399 519411 373433
rect 519445 373399 519488 373433
rect 519368 373233 519488 373399
rect 519368 373199 519411 373233
rect 519445 373199 519488 373233
rect 519368 373033 519488 373199
rect 519368 372999 519411 373033
rect 519445 372999 519488 373033
rect 519368 372833 519488 372999
rect 519368 372799 519411 372833
rect 519445 372799 519488 372833
rect 519368 372633 519488 372799
rect 519368 372599 519411 372633
rect 519445 372599 519488 372633
rect 517860 372062 517912 372068
rect 517860 372004 517912 372010
rect 517488 371855 517531 371889
rect 517565 371855 517608 371889
rect 517488 371689 517608 371855
rect 517488 371655 517531 371689
rect 517565 371655 517608 371689
rect 517488 371489 517608 371655
rect 517488 371455 517531 371489
rect 517565 371455 517608 371489
rect 517488 371289 517608 371455
rect 517488 371255 517531 371289
rect 517565 371255 517608 371289
rect 517488 371089 517608 371255
rect 517488 371055 517531 371089
rect 517565 371055 517608 371089
rect 517488 370889 517608 371055
rect 517488 370855 517531 370889
rect 517565 370855 517608 370889
rect 517488 370689 517608 370855
rect 517488 370655 517531 370689
rect 517565 370655 517608 370689
rect 517488 370489 517608 370655
rect 517488 370455 517531 370489
rect 517565 370455 517608 370489
rect 517488 370289 517608 370455
rect 517488 370255 517531 370289
rect 517565 370255 517608 370289
rect 517488 370089 517608 370255
rect 516469 370053 517433 370064
rect 515907 370046 517433 370053
rect 515907 369652 515919 370046
rect 516457 369652 516879 370046
rect 517417 369652 517433 370046
rect 515907 369643 517433 369652
rect 516469 369632 517433 369643
rect 517488 370055 517531 370089
rect 517565 370055 517608 370089
rect 517488 369889 517608 370055
rect 517488 369855 517531 369889
rect 517565 369855 517608 369889
rect 515907 369309 516469 369317
rect 515907 369290 515919 369309
rect 515832 369262 515919 369290
rect 515608 369111 515651 369145
rect 515685 369111 515728 369145
rect 515608 368945 515728 369111
rect 515608 368911 515651 368945
rect 515685 368911 515728 368945
rect 515608 368745 515728 368911
rect 515820 368934 515872 368940
rect 515907 368915 515919 369262
rect 516457 368915 516469 369309
rect 515907 368907 516469 368915
rect 516867 369309 517429 369317
rect 516867 368915 516879 369309
rect 517417 368915 517429 369309
rect 516867 368907 516908 368915
rect 515820 368876 515872 368882
rect 516960 368907 517429 368915
rect 517488 369145 517608 369855
rect 517488 369111 517531 369145
rect 517565 369111 517608 369145
rect 517488 368945 517608 369111
rect 517488 368911 517531 368945
rect 517565 368911 517608 368945
rect 516908 368876 516960 368882
rect 515608 368711 515651 368745
rect 515685 368711 515728 368745
rect 515608 368545 515728 368711
rect 515608 368511 515651 368545
rect 515685 368511 515728 368545
rect 515608 368345 515728 368511
rect 515608 368311 515651 368345
rect 515685 368311 515728 368345
rect 515608 368145 515728 368311
rect 515608 368111 515651 368145
rect 515685 368111 515728 368145
rect 515608 367945 515728 368111
rect 515608 367911 515651 367945
rect 515685 367911 515728 367945
rect 515608 367745 515728 367911
rect 515608 367711 515651 367745
rect 515685 367711 515728 367745
rect 515608 367545 515728 367711
rect 515608 367511 515651 367545
rect 515685 367511 515728 367545
rect 515608 367345 515728 367511
rect 515608 367311 515651 367345
rect 515685 367311 515728 367345
rect 515608 367145 515728 367311
rect 515608 367111 515651 367145
rect 515685 367111 515728 367145
rect 515608 366401 515728 367111
rect 515832 366456 515860 368876
rect 517488 368745 517608 368911
rect 517488 368711 517531 368745
rect 517565 368711 517608 368745
rect 517488 368545 517608 368711
rect 517488 368511 517531 368545
rect 517565 368511 517608 368545
rect 517488 368345 517608 368511
rect 517488 368311 517531 368345
rect 517565 368311 517608 368345
rect 517488 368145 517608 368311
rect 517488 368111 517531 368145
rect 517565 368111 517608 368145
rect 517488 367945 517608 368111
rect 517488 367911 517531 367945
rect 517565 367911 517608 367945
rect 517488 367745 517608 367911
rect 517488 367711 517531 367745
rect 517565 367711 517608 367745
rect 517488 367545 517608 367711
rect 517488 367511 517531 367545
rect 517565 367511 517608 367545
rect 517488 367345 517608 367511
rect 516469 367309 517433 367320
rect 515907 367302 517433 367309
rect 515907 366908 515919 367302
rect 516457 366908 516879 367302
rect 517417 366908 517433 367302
rect 515907 366899 517433 366908
rect 516469 366888 517433 366899
rect 517488 367311 517531 367345
rect 517565 367311 517608 367345
rect 517488 367145 517608 367311
rect 517488 367111 517531 367145
rect 517565 367111 517608 367145
rect 515907 366565 516469 366573
rect 515608 366367 515651 366401
rect 515685 366367 515728 366401
rect 515820 366450 515872 366456
rect 515820 366392 515872 366398
rect 515608 366201 515728 366367
rect 515608 366167 515651 366201
rect 515685 366167 515728 366201
rect 515608 366001 515728 366167
rect 515907 366171 515919 366565
rect 516457 366364 516469 366565
rect 516867 366565 517429 366573
rect 516457 366358 516484 366364
rect 516457 366300 516484 366306
rect 516457 366171 516469 366300
rect 515907 366163 516469 366171
rect 516867 366171 516879 366565
rect 517417 366171 517429 366565
rect 516867 366163 517429 366171
rect 517488 366401 517608 367111
rect 517488 366367 517531 366401
rect 517565 366367 517608 366401
rect 517488 366201 517608 366367
rect 517488 366167 517531 366201
rect 517565 366167 517608 366201
rect 515608 365967 515651 366001
rect 515685 365967 515728 366001
rect 515608 365801 515728 365967
rect 515608 365767 515651 365801
rect 515685 365767 515728 365801
rect 515608 365601 515728 365767
rect 515608 365567 515651 365601
rect 515685 365567 515728 365601
rect 515608 365401 515728 365567
rect 515608 365367 515651 365401
rect 515685 365367 515728 365401
rect 515608 365201 515728 365367
rect 515608 365167 515651 365201
rect 515685 365167 515728 365201
rect 515608 365001 515728 365167
rect 515608 364967 515651 365001
rect 515685 364967 515728 365001
rect 515608 364801 515728 364967
rect 515608 364767 515651 364801
rect 515685 364767 515728 364801
rect 515608 364601 515728 364767
rect 515608 364567 515651 364601
rect 515685 364567 515728 364601
rect 517488 366001 517608 366167
rect 517488 365967 517531 366001
rect 517565 365967 517608 366001
rect 517488 365801 517608 365967
rect 517488 365767 517531 365801
rect 517565 365767 517608 365801
rect 517488 365601 517608 365767
rect 517488 365567 517531 365601
rect 517565 365567 517608 365601
rect 517488 365401 517608 365567
rect 517488 365367 517531 365401
rect 517565 365367 517608 365401
rect 517488 365201 517608 365367
rect 517488 365167 517531 365201
rect 517565 365167 517608 365201
rect 517488 365001 517608 365167
rect 517488 364967 517531 365001
rect 517565 364967 517608 365001
rect 517488 364801 517608 364967
rect 517488 364767 517531 364801
rect 517565 364767 517608 364801
rect 517488 364601 517608 364767
rect 515608 364401 515728 364567
rect 516469 364565 517433 364576
rect 515608 364367 515651 364401
rect 515685 364367 515728 364401
rect 515608 361476 515728 364367
rect 515907 364558 517433 364565
rect 515907 364164 515919 364558
rect 516457 364164 516879 364558
rect 517417 364164 517433 364558
rect 515907 364155 517433 364164
rect 516469 364144 517433 364155
rect 517488 364567 517531 364601
rect 517565 364567 517608 364601
rect 517488 364401 517608 364567
rect 517488 364367 517531 364401
rect 517565 364367 517608 364401
rect 515608 359888 515610 361476
rect 515726 359888 515728 361476
rect 515608 359866 515728 359888
rect 513728 357440 513730 359028
rect 513846 357440 513848 359028
rect 513728 357418 513848 357440
rect 517488 359028 517608 364367
rect 519368 366401 519488 372599
rect 519572 374414 519679 374442
rect 519572 372252 519600 374414
rect 519667 374403 519679 374414
rect 520217 374403 520229 374797
rect 519667 374395 520229 374403
rect 520627 374797 521189 374805
rect 520627 374403 520639 374797
rect 521177 374403 521189 374797
rect 520627 374395 521189 374403
rect 521248 374633 521368 375343
rect 521248 374599 521291 374633
rect 521325 374599 521368 374633
rect 521248 374433 521368 374599
rect 521248 374399 521291 374433
rect 521325 374399 521368 374433
rect 520660 373540 520688 374395
rect 521248 374233 521368 374399
rect 521248 374199 521291 374233
rect 521325 374199 521368 374233
rect 521248 374033 521368 374199
rect 521248 373999 521291 374033
rect 521325 373999 521368 374033
rect 521248 373833 521368 373999
rect 521248 373799 521291 373833
rect 521325 373799 521368 373833
rect 521248 373633 521368 373799
rect 521248 373599 521291 373633
rect 521325 373599 521368 373633
rect 520648 373534 520700 373540
rect 520648 373476 520700 373482
rect 521248 373433 521368 373599
rect 521248 373399 521291 373433
rect 521325 373399 521368 373433
rect 521248 373233 521368 373399
rect 521248 373199 521291 373233
rect 521325 373199 521368 373233
rect 521248 373033 521368 373199
rect 521248 372999 521291 373033
rect 521325 372999 521368 373033
rect 521248 372833 521368 372999
rect 520229 372797 521193 372808
rect 519667 372790 521193 372797
rect 519667 372396 519679 372790
rect 520217 372396 520639 372790
rect 521177 372396 521193 372790
rect 519667 372387 521193 372396
rect 520229 372376 521193 372387
rect 521248 372799 521291 372833
rect 521325 372799 521368 372833
rect 521248 372633 521368 372799
rect 521248 372599 521291 372633
rect 521325 372599 521368 372633
rect 519560 372246 519612 372252
rect 519560 372188 519612 372194
rect 519667 366565 520229 366573
rect 519368 366367 519411 366401
rect 519445 366367 519488 366401
rect 519560 366450 519612 366456
rect 519667 366438 519679 366565
rect 519612 366410 519679 366438
rect 519560 366392 519612 366398
rect 519368 366201 519488 366367
rect 519368 366167 519411 366201
rect 519445 366167 519488 366201
rect 519368 366001 519488 366167
rect 519667 366171 519679 366410
rect 520217 366171 520229 366565
rect 519667 366163 520229 366171
rect 520627 366565 521189 366573
rect 520627 366171 520639 366565
rect 521177 366171 521189 366565
rect 520627 366163 521189 366171
rect 521248 366401 521368 372599
rect 521248 366367 521291 366401
rect 521325 366367 521368 366401
rect 521248 366201 521368 366367
rect 521248 366167 521291 366201
rect 521325 366167 521368 366201
rect 519368 365967 519411 366001
rect 519445 365967 519488 366001
rect 519368 365801 519488 365967
rect 519368 365767 519411 365801
rect 519445 365767 519488 365801
rect 519368 365601 519488 365767
rect 519368 365567 519411 365601
rect 519445 365567 519488 365601
rect 519368 365401 519488 365567
rect 519368 365367 519411 365401
rect 519445 365367 519488 365401
rect 519368 365201 519488 365367
rect 519368 365167 519411 365201
rect 519445 365167 519488 365201
rect 519368 365001 519488 365167
rect 519368 364967 519411 365001
rect 519445 364967 519488 365001
rect 519368 364801 519488 364967
rect 519368 364767 519411 364801
rect 519445 364767 519488 364801
rect 519368 364601 519488 364767
rect 519368 364567 519411 364601
rect 519445 364567 519488 364601
rect 521248 366001 521368 366167
rect 521248 365967 521291 366001
rect 521325 365967 521368 366001
rect 521248 365801 521368 365967
rect 521248 365767 521291 365801
rect 521325 365767 521368 365801
rect 521248 365601 521368 365767
rect 521248 365567 521291 365601
rect 521325 365567 521368 365601
rect 521248 365401 521368 365567
rect 521248 365367 521291 365401
rect 521325 365367 521368 365401
rect 521248 365201 521368 365367
rect 521248 365167 521291 365201
rect 521325 365167 521368 365201
rect 521248 365001 521368 365167
rect 521248 364967 521291 365001
rect 521325 364967 521368 365001
rect 521248 364801 521368 364967
rect 521248 364767 521291 364801
rect 521325 364767 521368 364801
rect 521248 364601 521368 364767
rect 519368 364401 519488 364567
rect 520229 364565 521193 364576
rect 519368 364367 519411 364401
rect 519445 364367 519488 364401
rect 519368 361476 519488 364367
rect 519667 364558 521193 364565
rect 519667 364164 519679 364558
rect 520217 364164 520639 364558
rect 521177 364164 521193 364558
rect 519667 364155 521193 364164
rect 520229 364144 521193 364155
rect 521248 364567 521291 364601
rect 521325 364567 521368 364601
rect 521248 364401 521368 364567
rect 521248 364367 521291 364401
rect 521325 364367 521368 364401
rect 519368 359888 519370 361476
rect 519486 359888 519488 361476
rect 519368 359866 519488 359888
rect 517488 357440 517490 359028
rect 517606 357440 517608 359028
rect 517488 357418 517608 357440
rect 521248 359028 521368 364367
rect 523128 411584 523248 411606
rect 523128 409996 523130 411584
rect 523246 409996 523248 411584
rect 523128 389941 523248 409996
rect 523423 390077 524713 390083
rect 523423 390043 523439 390077
rect 523473 390043 523511 390077
rect 523545 390043 523583 390077
rect 523617 390043 523655 390077
rect 523689 390043 523727 390077
rect 523761 390043 523799 390077
rect 523833 390043 523871 390077
rect 523905 390043 523943 390077
rect 523977 390043 524015 390077
rect 524049 390043 524087 390077
rect 524121 390043 524159 390077
rect 524193 390043 524231 390077
rect 524265 390043 524303 390077
rect 524337 390043 524375 390077
rect 524409 390043 524447 390077
rect 524481 390043 524519 390077
rect 524553 390043 524591 390077
rect 524625 390043 524663 390077
rect 524697 390043 524713 390077
rect 523423 390037 524713 390043
rect 523128 389907 523171 389941
rect 523205 389907 523248 389941
rect 523128 389622 523248 389907
rect 525008 389941 525128 412444
rect 528768 414032 528888 414054
rect 528768 412444 528770 414032
rect 528886 412444 528888 414032
rect 525008 389907 525051 389941
rect 525085 389907 525128 389941
rect 523423 389622 524713 389625
rect 523128 389619 524713 389622
rect 523128 389594 523439 389619
rect 523128 389541 523248 389594
rect 523423 389585 523439 389594
rect 523473 389585 523511 389619
rect 523545 389585 523583 389619
rect 523617 389585 523655 389619
rect 523689 389585 523727 389619
rect 523761 389585 523799 389619
rect 523833 389585 523871 389619
rect 523905 389585 523943 389619
rect 523977 389585 524015 389619
rect 524049 389585 524087 389619
rect 524121 389585 524159 389619
rect 524193 389585 524231 389619
rect 524265 389585 524303 389619
rect 524337 389585 524375 389619
rect 524409 389585 524447 389619
rect 524481 389585 524519 389619
rect 524553 389585 524591 389619
rect 524625 389585 524663 389619
rect 524697 389585 524713 389619
rect 523423 389579 524713 389585
rect 523128 389507 523171 389541
rect 523205 389507 523248 389541
rect 523128 389141 523248 389507
rect 524864 389545 524916 389548
rect 524864 389542 524947 389545
rect 524916 389533 524947 389542
rect 524941 389499 524947 389533
rect 524916 389490 524947 389499
rect 524864 389487 524947 389490
rect 525008 389541 525128 389907
rect 525008 389507 525051 389541
rect 525085 389507 525128 389541
rect 524864 389484 524916 389487
rect 523128 389107 523171 389141
rect 523205 389107 523248 389141
rect 523423 389161 524713 389167
rect 523423 389127 523439 389161
rect 523473 389127 523511 389161
rect 523545 389127 523583 389161
rect 523617 389127 523655 389161
rect 523689 389127 523727 389161
rect 523761 389127 523799 389161
rect 523833 389127 523871 389161
rect 523905 389127 523943 389161
rect 523977 389127 524015 389161
rect 524049 389127 524087 389161
rect 524121 389127 524159 389161
rect 524193 389127 524231 389161
rect 524265 389127 524303 389161
rect 524337 389127 524375 389161
rect 524409 389127 524447 389161
rect 524481 389127 524519 389161
rect 524553 389127 524591 389161
rect 524625 389127 524663 389161
rect 524697 389127 524713 389161
rect 523423 389121 524713 389127
rect 525008 389141 525128 389507
rect 523128 388741 523248 389107
rect 523128 388707 523171 388741
rect 523205 388707 523248 388741
rect 525008 389107 525051 389141
rect 525085 389107 525128 389141
rect 525008 388741 525128 389107
rect 523128 388341 523248 388707
rect 523423 388703 524713 388709
rect 523423 388669 523439 388703
rect 523473 388669 523511 388703
rect 523545 388669 523583 388703
rect 523617 388669 523655 388703
rect 523689 388669 523727 388703
rect 523761 388669 523799 388703
rect 523833 388669 523871 388703
rect 523905 388669 523943 388703
rect 523977 388669 524015 388703
rect 524049 388669 524087 388703
rect 524121 388669 524159 388703
rect 524193 388669 524231 388703
rect 524265 388669 524303 388703
rect 524337 388669 524375 388703
rect 524409 388669 524447 388703
rect 524481 388669 524519 388703
rect 524553 388669 524591 388703
rect 524625 388669 524663 388703
rect 524697 388669 524713 388703
rect 523423 388663 524713 388669
rect 525008 388707 525051 388741
rect 525085 388707 525128 388741
rect 523128 388307 523171 388341
rect 523205 388307 523248 388341
rect 523128 387941 523248 388307
rect 525008 388341 525128 388707
rect 525008 388307 525051 388341
rect 525085 388307 525128 388341
rect 523423 388245 524713 388251
rect 523423 388211 523439 388245
rect 523473 388211 523511 388245
rect 523545 388211 523583 388245
rect 523617 388211 523655 388245
rect 523689 388211 523727 388245
rect 523761 388211 523799 388245
rect 523833 388211 523871 388245
rect 523905 388211 523943 388245
rect 523977 388211 524015 388245
rect 524049 388211 524087 388245
rect 524121 388211 524159 388245
rect 524193 388211 524231 388245
rect 524265 388211 524303 388245
rect 524337 388211 524375 388245
rect 524409 388211 524447 388245
rect 524481 388211 524519 388245
rect 524553 388211 524591 388245
rect 524625 388211 524663 388245
rect 524697 388211 524713 388245
rect 523423 388205 524713 388211
rect 523128 387907 523171 387941
rect 523205 387907 523248 387941
rect 523128 387541 523248 387907
rect 525008 387941 525128 388307
rect 525008 387907 525051 387941
rect 525085 387907 525128 387941
rect 523423 387787 524713 387793
rect 523423 387753 523439 387787
rect 523473 387753 523511 387787
rect 523545 387753 523583 387787
rect 523617 387753 523655 387787
rect 523689 387753 523727 387787
rect 523761 387753 523799 387787
rect 523833 387753 523871 387787
rect 523905 387753 523943 387787
rect 523977 387753 524015 387787
rect 524049 387753 524087 387787
rect 524121 387753 524159 387787
rect 524193 387753 524231 387787
rect 524265 387753 524303 387787
rect 524337 387753 524375 387787
rect 524409 387753 524447 387787
rect 524481 387753 524519 387787
rect 524553 387753 524591 387787
rect 524625 387753 524663 387787
rect 524697 387753 524713 387787
rect 523423 387747 524713 387753
rect 523128 387507 523171 387541
rect 523205 387507 523248 387541
rect 523128 387141 523248 387507
rect 525008 387541 525128 387907
rect 525008 387507 525051 387541
rect 525085 387507 525128 387541
rect 523423 387329 524713 387335
rect 523423 387295 523439 387329
rect 523473 387295 523511 387329
rect 523545 387295 523583 387329
rect 523617 387295 523655 387329
rect 523689 387295 523727 387329
rect 523761 387295 523799 387329
rect 523833 387295 523871 387329
rect 523905 387295 523943 387329
rect 523977 387295 524015 387329
rect 524049 387295 524087 387329
rect 524121 387295 524159 387329
rect 524193 387295 524231 387329
rect 524265 387295 524303 387329
rect 524337 387295 524375 387329
rect 524409 387295 524447 387329
rect 524481 387295 524519 387329
rect 524553 387295 524591 387329
rect 524625 387295 524663 387329
rect 524697 387295 524713 387329
rect 523423 387289 524713 387295
rect 523128 387107 523171 387141
rect 523205 387107 523248 387141
rect 523128 386741 523248 387107
rect 525008 387141 525128 387507
rect 525008 387107 525051 387141
rect 525085 387107 525128 387141
rect 523423 386871 524713 386877
rect 523423 386837 523439 386871
rect 523473 386837 523511 386871
rect 523545 386837 523583 386871
rect 523617 386837 523655 386871
rect 523689 386837 523727 386871
rect 523761 386837 523799 386871
rect 523833 386837 523871 386871
rect 523905 386837 523943 386871
rect 523977 386837 524015 386871
rect 524049 386837 524087 386871
rect 524121 386837 524159 386871
rect 524193 386837 524231 386871
rect 524265 386837 524303 386871
rect 524337 386837 524375 386871
rect 524409 386837 524447 386871
rect 524481 386837 524519 386871
rect 524553 386837 524591 386871
rect 524625 386837 524663 386871
rect 524697 386837 524713 386871
rect 523423 386831 524713 386837
rect 523128 386707 523171 386741
rect 523205 386707 523248 386741
rect 523128 386341 523248 386707
rect 525008 386741 525128 387107
rect 525008 386707 525051 386741
rect 525085 386707 525128 386741
rect 523423 386413 524713 386419
rect 523423 386379 523439 386413
rect 523473 386379 523511 386413
rect 523545 386379 523583 386413
rect 523617 386379 523655 386413
rect 523689 386379 523727 386413
rect 523761 386379 523799 386413
rect 523833 386379 523871 386413
rect 523905 386379 523943 386413
rect 523977 386379 524015 386413
rect 524049 386379 524087 386413
rect 524121 386379 524159 386413
rect 524193 386379 524231 386413
rect 524265 386379 524303 386413
rect 524337 386379 524375 386413
rect 524409 386379 524447 386413
rect 524481 386379 524519 386413
rect 524553 386379 524591 386413
rect 524625 386379 524663 386413
rect 524697 386379 524713 386413
rect 523423 386373 524713 386379
rect 523128 386307 523171 386341
rect 523205 386307 523248 386341
rect 523128 385941 523248 386307
rect 525008 386341 525128 386707
rect 525008 386307 525051 386341
rect 525085 386307 525128 386341
rect 523128 385907 523171 385941
rect 523205 385907 523248 385941
rect 523423 385955 524713 385961
rect 523423 385921 523439 385955
rect 523473 385921 523511 385955
rect 523545 385921 523583 385955
rect 523617 385921 523655 385955
rect 523689 385921 523727 385955
rect 523761 385921 523799 385955
rect 523833 385921 523871 385955
rect 523905 385921 523943 385955
rect 523977 385921 524015 385955
rect 524049 385921 524087 385955
rect 524121 385921 524159 385955
rect 524193 385921 524231 385955
rect 524265 385921 524303 385955
rect 524337 385921 524375 385955
rect 524409 385921 524447 385955
rect 524481 385921 524519 385955
rect 524553 385921 524591 385955
rect 524625 385921 524663 385955
rect 524697 385921 524713 385955
rect 523423 385915 524713 385921
rect 525008 385941 525128 386307
rect 523128 385541 523248 385907
rect 523128 385507 523171 385541
rect 523205 385507 523248 385541
rect 523128 385141 523248 385507
rect 525008 385907 525051 385941
rect 525085 385907 525128 385941
rect 525008 385541 525128 385907
rect 525008 385507 525051 385541
rect 525085 385507 525128 385541
rect 523423 385497 524713 385503
rect 523423 385463 523439 385497
rect 523473 385463 523511 385497
rect 523545 385463 523583 385497
rect 523617 385463 523655 385497
rect 523689 385463 523727 385497
rect 523761 385463 523799 385497
rect 523833 385463 523871 385497
rect 523905 385463 523943 385497
rect 523977 385463 524015 385497
rect 524049 385463 524087 385497
rect 524121 385463 524159 385497
rect 524193 385463 524231 385497
rect 524265 385463 524303 385497
rect 524337 385463 524375 385497
rect 524409 385463 524447 385497
rect 524481 385463 524519 385497
rect 524553 385463 524591 385497
rect 524625 385463 524663 385497
rect 524697 385463 524713 385497
rect 523423 385457 524713 385463
rect 523128 385107 523171 385141
rect 523205 385107 523248 385141
rect 523128 384741 523248 385107
rect 525008 385141 525128 385507
rect 525008 385107 525051 385141
rect 525085 385107 525128 385141
rect 523423 385039 524713 385045
rect 523423 385005 523439 385039
rect 523473 385005 523511 385039
rect 523545 385005 523583 385039
rect 523617 385005 523655 385039
rect 523689 385005 523727 385039
rect 523761 385005 523799 385039
rect 523833 385005 523871 385039
rect 523905 385005 523943 385039
rect 523977 385005 524015 385039
rect 524049 385005 524087 385039
rect 524121 385005 524159 385039
rect 524193 385005 524231 385039
rect 524265 385005 524303 385039
rect 524337 385005 524375 385039
rect 524409 385005 524447 385039
rect 524481 385005 524519 385039
rect 524553 385005 524591 385039
rect 524625 385005 524663 385039
rect 524697 385005 524713 385039
rect 523423 384999 524713 385005
rect 523128 384707 523171 384741
rect 523205 384707 523248 384741
rect 523128 384341 523248 384707
rect 525008 384741 525128 385107
rect 525008 384707 525051 384741
rect 525085 384707 525128 384741
rect 523423 384581 524713 384587
rect 523423 384547 523439 384581
rect 523473 384547 523511 384581
rect 523545 384547 523583 384581
rect 523617 384547 523655 384581
rect 523689 384547 523727 384581
rect 523761 384547 523799 384581
rect 523833 384547 523871 384581
rect 523905 384547 523943 384581
rect 523977 384547 524015 384581
rect 524049 384547 524087 384581
rect 524121 384547 524159 384581
rect 524193 384547 524231 384581
rect 524265 384547 524303 384581
rect 524337 384547 524375 384581
rect 524409 384547 524447 384581
rect 524481 384547 524519 384581
rect 524553 384547 524591 384581
rect 524625 384547 524663 384581
rect 524697 384547 524713 384581
rect 523423 384541 524713 384547
rect 523128 384307 523171 384341
rect 523205 384307 523248 384341
rect 523128 383941 523248 384307
rect 525008 384341 525128 384707
rect 525008 384307 525051 384341
rect 525085 384307 525128 384341
rect 523423 384123 524713 384129
rect 523423 384089 523439 384123
rect 523473 384089 523511 384123
rect 523545 384089 523583 384123
rect 523617 384089 523655 384123
rect 523689 384089 523727 384123
rect 523761 384089 523799 384123
rect 523833 384089 523871 384123
rect 523905 384089 523943 384123
rect 523977 384089 524015 384123
rect 524049 384089 524087 384123
rect 524121 384089 524159 384123
rect 524193 384089 524231 384123
rect 524265 384089 524303 384123
rect 524337 384089 524375 384123
rect 524409 384089 524447 384123
rect 524481 384089 524519 384123
rect 524553 384089 524591 384123
rect 524625 384089 524663 384123
rect 524697 384089 524713 384123
rect 523423 384083 524713 384089
rect 523128 383907 523171 383941
rect 523205 383907 523248 383941
rect 523128 383541 523248 383907
rect 525008 383941 525128 384307
rect 525008 383907 525051 383941
rect 525085 383907 525128 383941
rect 523423 383665 524713 383671
rect 523423 383631 523439 383665
rect 523473 383631 523511 383665
rect 523545 383631 523583 383665
rect 523617 383631 523655 383665
rect 523689 383631 523727 383665
rect 523761 383631 523799 383665
rect 523833 383631 523871 383665
rect 523905 383631 523943 383665
rect 523977 383631 524015 383665
rect 524049 383631 524087 383665
rect 524121 383631 524159 383665
rect 524193 383631 524231 383665
rect 524265 383631 524303 383665
rect 524337 383631 524375 383665
rect 524409 383631 524447 383665
rect 524481 383631 524519 383665
rect 524553 383631 524591 383665
rect 524625 383631 524663 383665
rect 524697 383631 524713 383665
rect 523423 383625 524713 383631
rect 523128 383507 523171 383541
rect 523205 383507 523248 383541
rect 523128 383141 523248 383507
rect 525008 383541 525128 383907
rect 525008 383507 525051 383541
rect 525085 383507 525128 383541
rect 523423 383207 524713 383213
rect 523423 383173 523439 383207
rect 523473 383173 523511 383207
rect 523545 383173 523583 383207
rect 523617 383173 523655 383207
rect 523689 383173 523727 383207
rect 523761 383173 523799 383207
rect 523833 383173 523871 383207
rect 523905 383173 523943 383207
rect 523977 383173 524015 383207
rect 524049 383173 524087 383207
rect 524121 383173 524159 383207
rect 524193 383173 524231 383207
rect 524265 383173 524303 383207
rect 524337 383173 524375 383207
rect 524409 383173 524447 383207
rect 524481 383173 524519 383207
rect 524553 383173 524591 383207
rect 524625 383173 524663 383207
rect 524697 383173 524713 383207
rect 523423 383167 524713 383173
rect 523128 383107 523171 383141
rect 523205 383107 523248 383141
rect 523128 382741 523248 383107
rect 525008 383141 525128 383507
rect 525008 383107 525051 383141
rect 525085 383107 525128 383141
rect 523128 382707 523171 382741
rect 523205 382707 523248 382741
rect 523423 382749 524713 382755
rect 523423 382715 523439 382749
rect 523473 382715 523511 382749
rect 523545 382715 523583 382749
rect 523617 382715 523655 382749
rect 523689 382715 523727 382749
rect 523761 382715 523799 382749
rect 523833 382715 523871 382749
rect 523905 382715 523943 382749
rect 523977 382715 524015 382749
rect 524049 382715 524087 382749
rect 524121 382715 524159 382749
rect 524193 382715 524231 382749
rect 524265 382715 524303 382749
rect 524337 382715 524375 382749
rect 524409 382715 524447 382749
rect 524481 382715 524519 382749
rect 524553 382715 524591 382749
rect 524625 382715 524663 382749
rect 524697 382715 524713 382749
rect 523423 382709 524713 382715
rect 525008 382741 525128 383107
rect 523128 382341 523248 382707
rect 523128 382307 523171 382341
rect 523205 382307 523248 382341
rect 523128 381941 523248 382307
rect 525008 382707 525051 382741
rect 525085 382707 525128 382741
rect 525008 382341 525128 382707
rect 525008 382307 525051 382341
rect 525085 382307 525128 382341
rect 523423 382291 524713 382297
rect 523423 382257 523439 382291
rect 523473 382257 523511 382291
rect 523545 382257 523583 382291
rect 523617 382257 523655 382291
rect 523689 382257 523727 382291
rect 523761 382257 523799 382291
rect 523833 382257 523871 382291
rect 523905 382257 523943 382291
rect 523977 382257 524015 382291
rect 524049 382257 524087 382291
rect 524121 382257 524159 382291
rect 524193 382257 524231 382291
rect 524265 382257 524303 382291
rect 524337 382257 524375 382291
rect 524409 382257 524447 382291
rect 524481 382257 524519 382291
rect 524553 382257 524591 382291
rect 524625 382257 524663 382291
rect 524697 382257 524713 382291
rect 523423 382251 524713 382257
rect 523128 381907 523171 381941
rect 523205 381907 523248 381941
rect 523128 381541 523248 381907
rect 525008 381941 525128 382307
rect 525008 381907 525051 381941
rect 525085 381907 525128 381941
rect 523423 381833 524713 381839
rect 523423 381799 523439 381833
rect 523473 381799 523511 381833
rect 523545 381799 523583 381833
rect 523617 381799 523655 381833
rect 523689 381799 523727 381833
rect 523761 381799 523799 381833
rect 523833 381799 523871 381833
rect 523905 381799 523943 381833
rect 523977 381799 524015 381833
rect 524049 381799 524087 381833
rect 524121 381799 524159 381833
rect 524193 381799 524231 381833
rect 524265 381799 524303 381833
rect 524337 381799 524375 381833
rect 524409 381799 524447 381833
rect 524481 381799 524519 381833
rect 524553 381799 524591 381833
rect 524625 381799 524663 381833
rect 524697 381799 524713 381833
rect 523423 381793 524713 381799
rect 523128 381507 523171 381541
rect 523205 381507 523248 381541
rect 523128 381141 523248 381507
rect 525008 381541 525128 381907
rect 525008 381507 525051 381541
rect 525085 381507 525128 381541
rect 523423 381375 524713 381381
rect 523423 381341 523439 381375
rect 523473 381341 523511 381375
rect 523545 381341 523583 381375
rect 523617 381341 523655 381375
rect 523689 381341 523727 381375
rect 523761 381341 523799 381375
rect 523833 381341 523871 381375
rect 523905 381341 523943 381375
rect 523977 381341 524015 381375
rect 524049 381341 524087 381375
rect 524121 381341 524159 381375
rect 524193 381341 524231 381375
rect 524265 381341 524303 381375
rect 524337 381341 524375 381375
rect 524409 381341 524447 381375
rect 524481 381341 524519 381375
rect 524553 381341 524591 381375
rect 524625 381341 524663 381375
rect 524697 381341 524713 381375
rect 523423 381335 524713 381341
rect 523128 381107 523171 381141
rect 523205 381107 523248 381141
rect 523128 380741 523248 381107
rect 525008 381141 525128 381507
rect 525008 381107 525051 381141
rect 525085 381107 525128 381141
rect 523423 380917 524713 380923
rect 523423 380883 523439 380917
rect 523473 380883 523511 380917
rect 523545 380883 523583 380917
rect 523617 380883 523655 380917
rect 523689 380883 523727 380917
rect 523761 380883 523799 380917
rect 523833 380883 523871 380917
rect 523905 380883 523943 380917
rect 523977 380883 524015 380917
rect 524049 380883 524087 380917
rect 524121 380883 524159 380917
rect 524193 380883 524231 380917
rect 524265 380883 524303 380917
rect 524337 380883 524375 380917
rect 524409 380883 524447 380917
rect 524481 380883 524519 380917
rect 524553 380883 524591 380917
rect 524625 380883 524663 380917
rect 524697 380883 524713 380917
rect 523423 380877 524713 380883
rect 523128 380707 523171 380741
rect 523205 380707 523248 380741
rect 523128 380341 523248 380707
rect 525008 380741 525128 381107
rect 525008 380707 525051 380741
rect 525085 380707 525128 380741
rect 524808 380624 524836 380679
rect 524796 380618 524848 380624
rect 524796 380560 524848 380566
rect 523423 380459 524713 380465
rect 523423 380425 523439 380459
rect 523473 380425 523511 380459
rect 523545 380425 523583 380459
rect 523617 380425 523655 380459
rect 523689 380425 523727 380459
rect 523761 380425 523799 380459
rect 523833 380425 523871 380459
rect 523905 380425 523943 380459
rect 523977 380425 524015 380459
rect 524049 380425 524087 380459
rect 524121 380425 524159 380459
rect 524193 380425 524231 380459
rect 524265 380425 524303 380459
rect 524337 380425 524375 380459
rect 524409 380425 524447 380459
rect 524481 380425 524519 380459
rect 524553 380425 524591 380459
rect 524625 380425 524663 380459
rect 524697 380425 524713 380459
rect 523423 380419 524713 380425
rect 523128 380307 523171 380341
rect 523205 380307 523248 380341
rect 523128 379941 523248 380307
rect 525008 380341 525128 380707
rect 525008 380307 525051 380341
rect 525085 380307 525128 380341
rect 523423 380001 524713 380007
rect 523423 379967 523439 380001
rect 523473 379967 523511 380001
rect 523545 379967 523583 380001
rect 523617 379967 523655 380001
rect 523689 379967 523727 380001
rect 523761 379967 523799 380001
rect 523833 379967 523871 380001
rect 523905 379967 523943 380001
rect 523977 379967 524015 380001
rect 524049 379967 524087 380001
rect 524121 379967 524159 380001
rect 524193 379967 524231 380001
rect 524265 379967 524303 380001
rect 524337 379967 524375 380001
rect 524409 379967 524447 380001
rect 524481 379967 524519 380001
rect 524553 379967 524591 380001
rect 524625 379967 524663 380001
rect 524697 379967 524713 380001
rect 523423 379961 524713 379967
rect 523128 379907 523171 379941
rect 523205 379907 523248 379941
rect 523128 379541 523248 379907
rect 525008 379941 525128 380307
rect 525008 379907 525051 379941
rect 525085 379907 525128 379941
rect 523128 379507 523171 379541
rect 523205 379507 523248 379541
rect 523128 379141 523248 379507
rect 523423 379543 524713 379549
rect 523423 379509 523439 379543
rect 523473 379509 523511 379543
rect 523545 379509 523583 379543
rect 523617 379509 523655 379543
rect 523689 379509 523727 379543
rect 523761 379509 523799 379543
rect 523833 379509 523871 379543
rect 523905 379509 523943 379543
rect 523977 379509 524015 379543
rect 524049 379509 524087 379543
rect 524121 379509 524159 379543
rect 524193 379509 524231 379543
rect 524265 379509 524303 379543
rect 524337 379509 524375 379543
rect 524409 379509 524447 379543
rect 524481 379509 524519 379543
rect 524553 379509 524591 379543
rect 524625 379509 524663 379543
rect 524697 379509 524713 379543
rect 523423 379503 524713 379509
rect 525008 379541 525128 379907
rect 525008 379507 525051 379541
rect 525085 379507 525128 379541
rect 523128 379107 523171 379141
rect 523205 379107 523248 379141
rect 523128 378741 523248 379107
rect 525008 379141 525128 379507
rect 525008 379107 525051 379141
rect 525085 379107 525128 379141
rect 523423 379085 524713 379091
rect 523423 379051 523439 379085
rect 523473 379051 523511 379085
rect 523545 379051 523583 379085
rect 523617 379051 523655 379085
rect 523689 379051 523727 379085
rect 523761 379051 523799 379085
rect 523833 379051 523871 379085
rect 523905 379051 523943 379085
rect 523977 379051 524015 379085
rect 524049 379051 524087 379085
rect 524121 379051 524159 379085
rect 524193 379051 524231 379085
rect 524265 379051 524303 379085
rect 524337 379051 524375 379085
rect 524409 379051 524447 379085
rect 524481 379051 524519 379085
rect 524553 379051 524591 379085
rect 524625 379051 524663 379085
rect 524697 379051 524713 379085
rect 523423 379045 524713 379051
rect 523128 378707 523171 378741
rect 523205 378707 523248 378741
rect 523128 378341 523248 378707
rect 525008 378741 525128 379107
rect 525008 378707 525051 378741
rect 525085 378707 525128 378741
rect 523423 378627 524713 378633
rect 523423 378593 523439 378627
rect 523473 378593 523511 378627
rect 523545 378593 523583 378627
rect 523617 378593 523655 378627
rect 523689 378593 523727 378627
rect 523761 378593 523799 378627
rect 523833 378593 523871 378627
rect 523905 378593 523943 378627
rect 523977 378593 524015 378627
rect 524049 378593 524087 378627
rect 524121 378593 524159 378627
rect 524193 378593 524231 378627
rect 524265 378593 524303 378627
rect 524337 378593 524375 378627
rect 524409 378593 524447 378627
rect 524481 378593 524519 378627
rect 524553 378593 524591 378627
rect 524625 378593 524663 378627
rect 524697 378593 524713 378627
rect 523423 378587 524713 378593
rect 523128 378307 523171 378341
rect 523205 378307 523248 378341
rect 523128 377941 523248 378307
rect 525008 378341 525128 378707
rect 525008 378307 525051 378341
rect 525085 378307 525128 378341
rect 523423 378169 524713 378175
rect 523423 378135 523439 378169
rect 523473 378135 523511 378169
rect 523545 378135 523583 378169
rect 523617 378135 523655 378169
rect 523689 378135 523727 378169
rect 523761 378135 523799 378169
rect 523833 378135 523871 378169
rect 523905 378135 523943 378169
rect 523977 378135 524015 378169
rect 524049 378135 524087 378169
rect 524121 378135 524159 378169
rect 524193 378135 524231 378169
rect 524265 378135 524303 378169
rect 524337 378135 524375 378169
rect 524409 378135 524447 378169
rect 524481 378135 524519 378169
rect 524553 378135 524591 378169
rect 524625 378135 524663 378169
rect 524697 378135 524713 378169
rect 523423 378129 524713 378135
rect 523128 377907 523171 377941
rect 523205 377907 523248 377941
rect 523128 377541 523248 377907
rect 525008 377941 525128 378307
rect 525008 377907 525051 377941
rect 525085 377907 525128 377941
rect 523423 377711 524713 377717
rect 523423 377677 523439 377711
rect 523473 377677 523511 377711
rect 523545 377677 523583 377711
rect 523617 377677 523655 377711
rect 523689 377677 523727 377711
rect 523761 377677 523799 377711
rect 523833 377677 523871 377711
rect 523905 377677 523943 377711
rect 523977 377677 524015 377711
rect 524049 377677 524087 377711
rect 524121 377677 524159 377711
rect 524193 377677 524231 377711
rect 524265 377677 524303 377711
rect 524337 377677 524375 377711
rect 524409 377677 524447 377711
rect 524481 377677 524519 377711
rect 524553 377677 524591 377711
rect 524625 377677 524663 377711
rect 524697 377677 524713 377711
rect 523423 377671 524713 377677
rect 523128 377507 523171 377541
rect 523205 377507 523248 377541
rect 523128 377141 523248 377507
rect 525008 377541 525128 377907
rect 525008 377507 525051 377541
rect 525085 377507 525128 377541
rect 523423 377253 524713 377259
rect 523423 377219 523439 377253
rect 523473 377219 523511 377253
rect 523545 377219 523583 377253
rect 523617 377219 523655 377253
rect 523689 377219 523727 377253
rect 523761 377219 523799 377253
rect 523833 377219 523871 377253
rect 523905 377219 523943 377253
rect 523977 377219 524015 377253
rect 524049 377219 524087 377253
rect 524121 377219 524159 377253
rect 524193 377219 524231 377253
rect 524265 377219 524303 377253
rect 524337 377219 524375 377253
rect 524409 377219 524447 377253
rect 524481 377219 524519 377253
rect 524553 377219 524591 377253
rect 524625 377219 524663 377253
rect 524697 377219 524713 377253
rect 523423 377213 524713 377219
rect 523128 377107 523171 377141
rect 523205 377107 523248 377141
rect 523128 376741 523248 377107
rect 525008 377141 525128 377507
rect 525008 377107 525051 377141
rect 525085 377107 525128 377141
rect 523423 376795 524713 376801
rect 523423 376761 523439 376795
rect 523473 376761 523511 376795
rect 523545 376761 523583 376795
rect 523617 376761 523655 376795
rect 523689 376761 523727 376795
rect 523761 376761 523799 376795
rect 523833 376761 523871 376795
rect 523905 376761 523943 376795
rect 523977 376761 524015 376795
rect 524049 376761 524087 376795
rect 524121 376761 524159 376795
rect 524193 376761 524231 376795
rect 524265 376761 524303 376795
rect 524337 376761 524375 376795
rect 524409 376761 524447 376795
rect 524481 376761 524519 376795
rect 524553 376761 524591 376795
rect 524625 376761 524663 376795
rect 524697 376761 524713 376795
rect 523423 376755 524713 376761
rect 523128 376707 523171 376741
rect 523205 376707 523248 376741
rect 523128 376341 523248 376707
rect 525008 376741 525128 377107
rect 525008 376707 525051 376741
rect 525085 376707 525128 376741
rect 523128 376307 523171 376341
rect 523205 376307 523248 376341
rect 523128 375941 523248 376307
rect 523423 376337 524713 376343
rect 523423 376303 523439 376337
rect 523473 376303 523511 376337
rect 523545 376303 523583 376337
rect 523617 376303 523655 376337
rect 523689 376303 523727 376337
rect 523761 376303 523799 376337
rect 523833 376303 523871 376337
rect 523905 376303 523943 376337
rect 523977 376303 524015 376337
rect 524049 376303 524087 376337
rect 524121 376303 524159 376337
rect 524193 376303 524231 376337
rect 524265 376303 524303 376337
rect 524337 376303 524375 376337
rect 524409 376303 524447 376337
rect 524481 376303 524519 376337
rect 524553 376303 524591 376337
rect 524625 376303 524663 376337
rect 524697 376303 524713 376337
rect 523423 376297 524713 376303
rect 525008 376341 525128 376707
rect 525008 376307 525051 376341
rect 525085 376307 525128 376341
rect 523128 375907 523171 375941
rect 523205 375907 523248 375941
rect 523128 375541 523248 375907
rect 525008 375941 525128 376307
rect 525008 375907 525051 375941
rect 525085 375907 525128 375941
rect 523423 375879 524713 375885
rect 523423 375845 523439 375879
rect 523473 375845 523511 375879
rect 523545 375845 523583 375879
rect 523617 375845 523655 375879
rect 523689 375845 523727 375879
rect 523761 375845 523799 375879
rect 523833 375845 523871 375879
rect 523905 375845 523943 375879
rect 523977 375845 524015 375879
rect 524049 375845 524087 375879
rect 524121 375845 524159 375879
rect 524193 375845 524231 375879
rect 524265 375845 524303 375879
rect 524337 375845 524375 375879
rect 524409 375845 524447 375879
rect 524481 375845 524519 375879
rect 524553 375845 524591 375879
rect 524625 375845 524663 375879
rect 524697 375845 524713 375879
rect 523423 375839 524713 375845
rect 523128 375507 523171 375541
rect 523205 375507 523248 375541
rect 523128 375141 523248 375507
rect 525008 375541 525128 375907
rect 525008 375507 525051 375541
rect 525085 375507 525128 375541
rect 523423 375421 524713 375427
rect 523423 375387 523439 375421
rect 523473 375387 523511 375421
rect 523545 375387 523583 375421
rect 523617 375387 523655 375421
rect 523689 375387 523727 375421
rect 523761 375387 523799 375421
rect 523833 375387 523871 375421
rect 523905 375387 523943 375421
rect 523977 375387 524015 375421
rect 524049 375387 524087 375421
rect 524121 375387 524159 375421
rect 524193 375387 524231 375421
rect 524265 375387 524303 375421
rect 524337 375387 524375 375421
rect 524409 375387 524447 375421
rect 524481 375387 524519 375421
rect 524553 375387 524591 375421
rect 524625 375387 524663 375421
rect 524697 375387 524713 375421
rect 523423 375381 524713 375387
rect 523128 375107 523171 375141
rect 523205 375107 523248 375141
rect 523128 374741 523248 375107
rect 525008 375141 525128 375507
rect 525008 375107 525051 375141
rect 525085 375107 525128 375141
rect 523423 374963 524713 374969
rect 523423 374929 523439 374963
rect 523473 374929 523511 374963
rect 523545 374929 523583 374963
rect 523617 374929 523655 374963
rect 523689 374929 523727 374963
rect 523761 374929 523799 374963
rect 523833 374929 523871 374963
rect 523905 374929 523943 374963
rect 523977 374929 524015 374963
rect 524049 374929 524087 374963
rect 524121 374929 524159 374963
rect 524193 374929 524231 374963
rect 524265 374929 524303 374963
rect 524337 374929 524375 374963
rect 524409 374929 524447 374963
rect 524481 374929 524519 374963
rect 524553 374929 524591 374963
rect 524625 374929 524663 374963
rect 524697 374929 524713 374963
rect 523423 374923 524713 374929
rect 523128 374707 523171 374741
rect 523205 374707 523248 374741
rect 523128 374341 523248 374707
rect 525008 374741 525128 375107
rect 525008 374707 525051 374741
rect 525085 374707 525128 374741
rect 523423 374505 524713 374511
rect 523423 374471 523439 374505
rect 523473 374471 523511 374505
rect 523545 374471 523583 374505
rect 523617 374471 523655 374505
rect 523689 374471 523727 374505
rect 523761 374471 523799 374505
rect 523833 374471 523871 374505
rect 523905 374471 523943 374505
rect 523977 374471 524015 374505
rect 524049 374471 524087 374505
rect 524121 374471 524159 374505
rect 524193 374471 524231 374505
rect 524265 374471 524303 374505
rect 524337 374471 524375 374505
rect 524409 374471 524447 374505
rect 524481 374471 524519 374505
rect 524553 374471 524591 374505
rect 524625 374471 524663 374505
rect 524697 374471 524713 374505
rect 523423 374465 524713 374471
rect 523128 374307 523171 374341
rect 523205 374307 523248 374341
rect 523128 373941 523248 374307
rect 525008 374341 525128 374707
rect 525008 374307 525051 374341
rect 525085 374307 525128 374341
rect 523423 374047 524713 374053
rect 523423 374013 523439 374047
rect 523473 374013 523511 374047
rect 523545 374013 523583 374047
rect 523617 374013 523655 374047
rect 523689 374013 523727 374047
rect 523761 374013 523799 374047
rect 523833 374013 523871 374047
rect 523905 374013 523943 374047
rect 523977 374013 524015 374047
rect 524049 374013 524087 374047
rect 524121 374013 524159 374047
rect 524193 374013 524231 374047
rect 524265 374013 524303 374047
rect 524337 374013 524375 374047
rect 524409 374013 524447 374047
rect 524481 374013 524519 374047
rect 524553 374013 524591 374047
rect 524625 374013 524663 374047
rect 524697 374013 524713 374047
rect 523423 374007 524713 374013
rect 523128 373907 523171 373941
rect 523205 373907 523248 373941
rect 523128 373541 523248 373907
rect 525008 373941 525128 374307
rect 525008 373907 525051 373941
rect 525085 373907 525128 373941
rect 523423 373589 524713 373595
rect 523423 373555 523439 373589
rect 523473 373555 523511 373589
rect 523545 373555 523583 373589
rect 523617 373555 523655 373589
rect 523689 373555 523727 373589
rect 523761 373555 523799 373589
rect 523833 373555 523871 373589
rect 523905 373555 523943 373589
rect 523977 373555 524015 373589
rect 524049 373555 524087 373589
rect 524121 373555 524159 373589
rect 524193 373555 524231 373589
rect 524265 373555 524303 373589
rect 524337 373555 524375 373589
rect 524409 373555 524447 373589
rect 524481 373555 524519 373589
rect 524553 373555 524591 373589
rect 524625 373555 524663 373589
rect 524697 373555 524713 373589
rect 523423 373549 524713 373555
rect 523128 373507 523171 373541
rect 523205 373507 523248 373541
rect 523128 373141 523248 373507
rect 523128 373107 523171 373141
rect 523205 373107 523248 373141
rect 525008 373541 525128 373907
rect 525008 373507 525051 373541
rect 525085 373507 525128 373541
rect 525008 373141 525128 373507
rect 523128 372741 523248 373107
rect 523423 373131 524713 373137
rect 523423 373097 523439 373131
rect 523473 373097 523511 373131
rect 523545 373097 523583 373131
rect 523617 373097 523655 373131
rect 523689 373097 523727 373131
rect 523761 373097 523799 373131
rect 523833 373097 523871 373131
rect 523905 373097 523943 373131
rect 523977 373097 524015 373131
rect 524049 373097 524087 373131
rect 524121 373097 524159 373131
rect 524193 373097 524231 373131
rect 524265 373097 524303 373131
rect 524337 373097 524375 373131
rect 524409 373097 524447 373131
rect 524481 373097 524519 373131
rect 524553 373097 524591 373131
rect 524625 373097 524663 373131
rect 524697 373097 524713 373131
rect 523423 373091 524713 373097
rect 525008 373107 525051 373141
rect 525085 373107 525128 373141
rect 523128 372707 523171 372741
rect 523205 372707 523248 372741
rect 523128 372341 523248 372707
rect 525008 372741 525128 373107
rect 525008 372707 525051 372741
rect 525085 372707 525128 372741
rect 523423 372673 524713 372679
rect 523423 372639 523439 372673
rect 523473 372639 523511 372673
rect 523545 372639 523583 372673
rect 523617 372639 523655 372673
rect 523689 372639 523727 372673
rect 523761 372639 523799 372673
rect 523833 372639 523871 372673
rect 523905 372639 523943 372673
rect 523977 372639 524015 372673
rect 524049 372639 524087 372673
rect 524121 372639 524159 372673
rect 524193 372639 524231 372673
rect 524265 372639 524303 372673
rect 524337 372639 524375 372673
rect 524409 372639 524447 372673
rect 524481 372639 524519 372673
rect 524553 372639 524591 372673
rect 524625 372639 524663 372673
rect 524697 372639 524713 372673
rect 523423 372633 524713 372639
rect 523128 372307 523171 372341
rect 523205 372307 523248 372341
rect 523128 371941 523248 372307
rect 525008 372341 525128 372707
rect 525008 372307 525051 372341
rect 525085 372307 525128 372341
rect 523423 372215 524713 372221
rect 523423 372181 523439 372215
rect 523473 372181 523511 372215
rect 523545 372181 523583 372215
rect 523617 372181 523655 372215
rect 523689 372181 523727 372215
rect 523761 372181 523799 372215
rect 523833 372181 523871 372215
rect 523905 372181 523943 372215
rect 523977 372181 524015 372215
rect 524049 372181 524087 372215
rect 524121 372181 524159 372215
rect 524193 372181 524231 372215
rect 524265 372181 524303 372215
rect 524337 372181 524375 372215
rect 524409 372181 524447 372215
rect 524481 372181 524519 372215
rect 524553 372181 524591 372215
rect 524625 372181 524663 372215
rect 524697 372181 524713 372215
rect 523423 372175 524713 372181
rect 523128 371907 523171 371941
rect 523205 371907 523248 371941
rect 523128 371541 523248 371907
rect 525008 371941 525128 372307
rect 525008 371907 525051 371941
rect 525085 371907 525128 371941
rect 523423 371757 524713 371763
rect 523423 371723 523439 371757
rect 523473 371723 523511 371757
rect 523545 371723 523583 371757
rect 523617 371723 523655 371757
rect 523689 371723 523727 371757
rect 523761 371723 523799 371757
rect 523833 371723 523871 371757
rect 523905 371723 523943 371757
rect 523977 371723 524015 371757
rect 524049 371723 524087 371757
rect 524121 371723 524159 371757
rect 524193 371723 524231 371757
rect 524265 371723 524303 371757
rect 524337 371723 524375 371757
rect 524409 371723 524447 371757
rect 524481 371723 524519 371757
rect 524553 371723 524591 371757
rect 524625 371723 524663 371757
rect 524697 371723 524713 371757
rect 523423 371717 524713 371723
rect 523128 371507 523171 371541
rect 523205 371507 523248 371541
rect 523128 371141 523248 371507
rect 525008 371541 525128 371907
rect 525008 371507 525051 371541
rect 525085 371507 525128 371541
rect 523423 371299 524713 371305
rect 523423 371265 523439 371299
rect 523473 371265 523511 371299
rect 523545 371265 523583 371299
rect 523617 371265 523655 371299
rect 523689 371265 523727 371299
rect 523761 371265 523799 371299
rect 523833 371265 523871 371299
rect 523905 371265 523943 371299
rect 523977 371265 524015 371299
rect 524049 371265 524087 371299
rect 524121 371265 524159 371299
rect 524193 371265 524231 371299
rect 524265 371265 524303 371299
rect 524337 371265 524375 371299
rect 524409 371265 524447 371299
rect 524481 371265 524519 371299
rect 524553 371265 524591 371299
rect 524625 371265 524663 371299
rect 524697 371265 524713 371299
rect 523423 371259 524713 371265
rect 523128 371107 523171 371141
rect 523205 371107 523248 371141
rect 523128 370741 523248 371107
rect 525008 371141 525128 371507
rect 525008 371107 525051 371141
rect 525085 371107 525128 371141
rect 524660 370958 524712 370964
rect 524660 370900 524712 370906
rect 524672 370847 524700 370900
rect 523423 370841 524713 370847
rect 523423 370807 523439 370841
rect 523473 370807 523511 370841
rect 523545 370807 523583 370841
rect 523617 370807 523655 370841
rect 523689 370807 523727 370841
rect 523761 370807 523799 370841
rect 523833 370807 523871 370841
rect 523905 370807 523943 370841
rect 523977 370807 524015 370841
rect 524049 370807 524087 370841
rect 524121 370807 524159 370841
rect 524193 370807 524231 370841
rect 524265 370807 524303 370841
rect 524337 370807 524375 370841
rect 524409 370807 524447 370841
rect 524481 370807 524519 370841
rect 524553 370807 524591 370841
rect 524625 370807 524663 370841
rect 524697 370807 524713 370841
rect 523423 370801 524713 370807
rect 523128 370707 523171 370741
rect 523205 370707 523248 370741
rect 523128 370341 523248 370707
rect 525008 370741 525128 371107
rect 525008 370707 525051 370741
rect 525085 370707 525128 370741
rect 523423 370383 524713 370389
rect 523423 370349 523439 370383
rect 523473 370349 523511 370383
rect 523545 370349 523583 370383
rect 523617 370349 523655 370383
rect 523689 370349 523727 370383
rect 523761 370349 523799 370383
rect 523833 370349 523871 370383
rect 523905 370349 523943 370383
rect 523977 370349 524015 370383
rect 524049 370349 524087 370383
rect 524121 370349 524159 370383
rect 524193 370349 524231 370383
rect 524265 370349 524303 370383
rect 524337 370349 524375 370383
rect 524409 370349 524447 370383
rect 524481 370349 524519 370383
rect 524553 370349 524591 370383
rect 524625 370349 524663 370383
rect 524697 370349 524713 370383
rect 523423 370343 524713 370349
rect 523128 370307 523171 370341
rect 523205 370307 523248 370341
rect 523128 369941 523248 370307
rect 523128 369907 523171 369941
rect 523205 369907 523248 369941
rect 525008 370341 525128 370707
rect 525008 370307 525051 370341
rect 525085 370307 525128 370341
rect 525008 369941 525128 370307
rect 523128 369541 523248 369907
rect 523423 369925 524713 369931
rect 523423 369891 523439 369925
rect 523473 369891 523511 369925
rect 523545 369891 523583 369925
rect 523617 369891 523655 369925
rect 523689 369891 523727 369925
rect 523761 369891 523799 369925
rect 523833 369891 523871 369925
rect 523905 369891 523943 369925
rect 523977 369891 524015 369925
rect 524049 369891 524087 369925
rect 524121 369891 524159 369925
rect 524193 369891 524231 369925
rect 524265 369891 524303 369925
rect 524337 369891 524375 369925
rect 524409 369891 524447 369925
rect 524481 369891 524519 369925
rect 524553 369891 524591 369925
rect 524625 369891 524663 369925
rect 524697 369891 524713 369925
rect 523423 369885 524713 369891
rect 525008 369907 525051 369941
rect 525085 369907 525128 369941
rect 523128 369507 523171 369541
rect 523205 369507 523248 369541
rect 523128 369141 523248 369507
rect 525008 369541 525128 369907
rect 525008 369507 525051 369541
rect 525085 369507 525128 369541
rect 523423 369467 524713 369473
rect 523423 369433 523439 369467
rect 523473 369433 523511 369467
rect 523545 369433 523583 369467
rect 523617 369433 523655 369467
rect 523689 369433 523727 369467
rect 523761 369433 523799 369467
rect 523833 369433 523871 369467
rect 523905 369433 523943 369467
rect 523977 369433 524015 369467
rect 524049 369433 524087 369467
rect 524121 369433 524159 369467
rect 524193 369433 524231 369467
rect 524265 369433 524303 369467
rect 524337 369433 524375 369467
rect 524409 369433 524447 369467
rect 524481 369433 524519 369467
rect 524553 369433 524591 369467
rect 524625 369433 524663 369467
rect 524697 369433 524713 369467
rect 523423 369427 524713 369433
rect 523128 369107 523171 369141
rect 523205 369107 523248 369141
rect 523128 368741 523248 369107
rect 525008 369141 525128 369507
rect 525008 369107 525051 369141
rect 525085 369107 525128 369141
rect 523423 369009 524713 369015
rect 523423 368975 523439 369009
rect 523473 368975 523511 369009
rect 523545 368975 523583 369009
rect 523617 368975 523655 369009
rect 523689 368975 523727 369009
rect 523761 368975 523799 369009
rect 523833 368975 523871 369009
rect 523905 368975 523943 369009
rect 523977 368975 524015 369009
rect 524049 368975 524087 369009
rect 524121 368975 524159 369009
rect 524193 368975 524231 369009
rect 524265 368975 524303 369009
rect 524337 368975 524375 369009
rect 524409 368975 524447 369009
rect 524481 368975 524519 369009
rect 524553 368975 524591 369009
rect 524625 368975 524663 369009
rect 524697 368975 524713 369009
rect 523423 368969 524713 368975
rect 523128 368707 523171 368741
rect 523205 368707 523248 368741
rect 523128 368341 523248 368707
rect 525008 368741 525128 369107
rect 525008 368707 525051 368741
rect 525085 368707 525128 368741
rect 523423 368551 524713 368557
rect 523423 368517 523439 368551
rect 523473 368517 523511 368551
rect 523545 368517 523583 368551
rect 523617 368517 523655 368551
rect 523689 368517 523727 368551
rect 523761 368517 523799 368551
rect 523833 368517 523871 368551
rect 523905 368517 523943 368551
rect 523977 368517 524015 368551
rect 524049 368517 524087 368551
rect 524121 368517 524159 368551
rect 524193 368517 524231 368551
rect 524265 368517 524303 368551
rect 524337 368517 524375 368551
rect 524409 368517 524447 368551
rect 524481 368517 524519 368551
rect 524553 368517 524591 368551
rect 524625 368517 524663 368551
rect 524697 368517 524713 368551
rect 523423 368511 524713 368517
rect 523128 368307 523171 368341
rect 523205 368307 523248 368341
rect 523128 367941 523248 368307
rect 525008 368341 525128 368707
rect 525008 368307 525051 368341
rect 525085 368307 525128 368341
rect 523423 368093 524713 368099
rect 523423 368059 523439 368093
rect 523473 368059 523511 368093
rect 523545 368059 523583 368093
rect 523617 368059 523655 368093
rect 523689 368059 523727 368093
rect 523761 368059 523799 368093
rect 523833 368059 523871 368093
rect 523905 368059 523943 368093
rect 523977 368059 524015 368093
rect 524049 368059 524087 368093
rect 524121 368059 524159 368093
rect 524193 368059 524231 368093
rect 524265 368059 524303 368093
rect 524337 368059 524375 368093
rect 524409 368059 524447 368093
rect 524481 368059 524519 368093
rect 524553 368059 524591 368093
rect 524625 368059 524663 368093
rect 524697 368059 524713 368093
rect 523423 368053 524713 368059
rect 523128 367907 523171 367941
rect 523205 367907 523248 367941
rect 523128 367541 523248 367907
rect 525008 367941 525128 368307
rect 525008 367907 525051 367941
rect 525085 367907 525128 367941
rect 523423 367635 524713 367641
rect 523423 367601 523439 367635
rect 523473 367601 523511 367635
rect 523545 367601 523583 367635
rect 523617 367601 523655 367635
rect 523689 367601 523727 367635
rect 523761 367601 523799 367635
rect 523833 367601 523871 367635
rect 523905 367601 523943 367635
rect 523977 367601 524015 367635
rect 524049 367601 524087 367635
rect 524121 367601 524159 367635
rect 524193 367601 524231 367635
rect 524265 367601 524303 367635
rect 524337 367601 524375 367635
rect 524409 367601 524447 367635
rect 524481 367601 524519 367635
rect 524553 367601 524591 367635
rect 524625 367601 524663 367635
rect 524697 367601 524713 367635
rect 523423 367595 524713 367601
rect 523128 367507 523171 367541
rect 523205 367507 523248 367541
rect 523128 367141 523248 367507
rect 525008 367541 525128 367907
rect 525008 367507 525051 367541
rect 525085 367507 525128 367541
rect 523128 367107 523171 367141
rect 523205 367107 523248 367141
rect 523423 367177 524713 367183
rect 523423 367143 523439 367177
rect 523473 367143 523511 367177
rect 523545 367143 523583 367177
rect 523617 367143 523655 367177
rect 523689 367143 523727 367177
rect 523761 367143 523799 367177
rect 523833 367143 523871 367177
rect 523905 367143 523943 367177
rect 523977 367143 524015 367177
rect 524049 367143 524087 367177
rect 524121 367143 524159 367177
rect 524193 367143 524231 367177
rect 524265 367143 524303 367177
rect 524337 367143 524375 367177
rect 524409 367143 524447 367177
rect 524481 367143 524519 367177
rect 524553 367143 524591 367177
rect 524625 367143 524663 367177
rect 524697 367143 524713 367177
rect 523423 367137 524713 367143
rect 525008 367141 525128 367507
rect 523128 366741 523248 367107
rect 523128 366707 523171 366741
rect 523205 366707 523248 366741
rect 525008 367107 525051 367141
rect 525085 367107 525128 367141
rect 525008 366741 525128 367107
rect 523128 366341 523248 366707
rect 523423 366719 524713 366725
rect 523423 366685 523439 366719
rect 523473 366685 523511 366719
rect 523545 366685 523583 366719
rect 523617 366685 523655 366719
rect 523689 366685 523727 366719
rect 523761 366685 523799 366719
rect 523833 366685 523871 366719
rect 523905 366685 523943 366719
rect 523977 366685 524015 366719
rect 524049 366685 524087 366719
rect 524121 366685 524159 366719
rect 524193 366685 524231 366719
rect 524265 366685 524303 366719
rect 524337 366685 524375 366719
rect 524409 366685 524447 366719
rect 524481 366685 524519 366719
rect 524553 366685 524591 366719
rect 524625 366685 524663 366719
rect 524697 366685 524713 366719
rect 523423 366679 524713 366685
rect 525008 366707 525051 366741
rect 525085 366707 525128 366741
rect 523128 366307 523171 366341
rect 523205 366307 523248 366341
rect 523128 365941 523248 366307
rect 525008 366341 525128 366707
rect 525008 366307 525051 366341
rect 525085 366307 525128 366341
rect 523423 366261 524713 366267
rect 523423 366227 523439 366261
rect 523473 366227 523511 366261
rect 523545 366227 523583 366261
rect 523617 366227 523655 366261
rect 523689 366227 523727 366261
rect 523761 366227 523799 366261
rect 523833 366227 523871 366261
rect 523905 366227 523943 366261
rect 523977 366227 524015 366261
rect 524049 366227 524087 366261
rect 524121 366227 524159 366261
rect 524193 366227 524231 366261
rect 524265 366227 524303 366261
rect 524337 366227 524375 366261
rect 524409 366227 524447 366261
rect 524481 366227 524519 366261
rect 524553 366227 524591 366261
rect 524625 366227 524663 366261
rect 524697 366227 524713 366261
rect 523423 366221 524713 366227
rect 523128 365907 523171 365941
rect 523205 365907 523248 365941
rect 523128 365541 523248 365907
rect 525008 365941 525128 366307
rect 525008 365907 525051 365941
rect 525085 365907 525128 365941
rect 523423 365803 524713 365809
rect 523423 365769 523439 365803
rect 523473 365769 523511 365803
rect 523545 365769 523583 365803
rect 523617 365769 523655 365803
rect 523689 365769 523727 365803
rect 523761 365769 523799 365803
rect 523833 365769 523871 365803
rect 523905 365769 523943 365803
rect 523977 365769 524015 365803
rect 524049 365769 524087 365803
rect 524121 365769 524159 365803
rect 524193 365769 524231 365803
rect 524265 365769 524303 365803
rect 524337 365769 524375 365803
rect 524409 365769 524447 365803
rect 524481 365769 524519 365803
rect 524553 365769 524591 365803
rect 524625 365769 524663 365803
rect 524697 365769 524713 365803
rect 523423 365763 524713 365769
rect 523128 365507 523171 365541
rect 523205 365507 523248 365541
rect 523128 365141 523248 365507
rect 525008 365541 525128 365907
rect 525008 365507 525051 365541
rect 525085 365507 525128 365541
rect 523423 365345 524713 365351
rect 523423 365311 523439 365345
rect 523473 365311 523511 365345
rect 523545 365311 523583 365345
rect 523617 365311 523655 365345
rect 523689 365311 523727 365345
rect 523761 365311 523799 365345
rect 523833 365311 523871 365345
rect 523905 365311 523943 365345
rect 523977 365311 524015 365345
rect 524049 365311 524087 365345
rect 524121 365311 524159 365345
rect 524193 365311 524231 365345
rect 524265 365311 524303 365345
rect 524337 365311 524375 365345
rect 524409 365311 524447 365345
rect 524481 365311 524519 365345
rect 524553 365311 524591 365345
rect 524625 365311 524663 365345
rect 524697 365311 524713 365345
rect 523423 365305 524713 365311
rect 523128 365107 523171 365141
rect 523205 365107 523248 365141
rect 523128 364741 523248 365107
rect 525008 365141 525128 365507
rect 525008 365107 525051 365141
rect 525085 365107 525128 365141
rect 523423 364887 524713 364893
rect 523423 364853 523439 364887
rect 523473 364853 523511 364887
rect 523545 364853 523583 364887
rect 523617 364853 523655 364887
rect 523689 364853 523727 364887
rect 523761 364853 523799 364887
rect 523833 364853 523871 364887
rect 523905 364853 523943 364887
rect 523977 364853 524015 364887
rect 524049 364853 524087 364887
rect 524121 364853 524159 364887
rect 524193 364853 524231 364887
rect 524265 364853 524303 364887
rect 524337 364853 524375 364887
rect 524409 364853 524447 364887
rect 524481 364853 524519 364887
rect 524553 364853 524591 364887
rect 524625 364853 524663 364887
rect 524697 364853 524713 364887
rect 523423 364847 524713 364853
rect 523128 364707 523171 364741
rect 523205 364707 523248 364741
rect 523128 364341 523248 364707
rect 525008 364741 525128 365107
rect 525008 364707 525051 364741
rect 525085 364707 525128 364741
rect 523423 364429 524713 364435
rect 523423 364395 523439 364429
rect 523473 364395 523511 364429
rect 523545 364395 523583 364429
rect 523617 364395 523655 364429
rect 523689 364395 523727 364429
rect 523761 364395 523799 364429
rect 523833 364395 523871 364429
rect 523905 364395 523943 364429
rect 523977 364395 524015 364429
rect 524049 364395 524087 364429
rect 524121 364395 524159 364429
rect 524193 364395 524231 364429
rect 524265 364395 524303 364429
rect 524337 364395 524375 364429
rect 524409 364395 524447 364429
rect 524481 364395 524519 364429
rect 524553 364395 524591 364429
rect 524625 364395 524663 364429
rect 524697 364395 524713 364429
rect 523423 364389 524713 364395
rect 523128 364307 523171 364341
rect 523205 364307 523248 364341
rect 523128 363941 523248 364307
rect 525008 364341 525128 364707
rect 525008 364307 525051 364341
rect 525085 364307 525128 364341
rect 523128 363907 523171 363941
rect 523205 363907 523248 363941
rect 523423 363971 524713 363977
rect 523423 363937 523439 363971
rect 523473 363937 523511 363971
rect 523545 363937 523583 363971
rect 523617 363937 523655 363971
rect 523689 363937 523727 363971
rect 523761 363937 523799 363971
rect 523833 363937 523871 363971
rect 523905 363937 523943 363971
rect 523977 363937 524015 363971
rect 524049 363937 524087 363971
rect 524121 363937 524159 363971
rect 524193 363937 524231 363971
rect 524265 363937 524303 363971
rect 524337 363937 524375 363971
rect 524409 363937 524447 363971
rect 524481 363937 524519 363971
rect 524553 363937 524591 363971
rect 524625 363937 524663 363971
rect 524697 363937 524713 363971
rect 523423 363931 524713 363937
rect 525008 363941 525128 364307
rect 523128 363541 523248 363907
rect 523128 363507 523171 363541
rect 523205 363507 523248 363541
rect 525008 363907 525051 363941
rect 525085 363907 525128 363941
rect 525008 363541 525128 363907
rect 523128 363141 523248 363507
rect 523423 363513 524713 363519
rect 523423 363479 523439 363513
rect 523473 363479 523511 363513
rect 523545 363479 523583 363513
rect 523617 363479 523655 363513
rect 523689 363479 523727 363513
rect 523761 363479 523799 363513
rect 523833 363479 523871 363513
rect 523905 363479 523943 363513
rect 523977 363479 524015 363513
rect 524049 363479 524087 363513
rect 524121 363479 524159 363513
rect 524193 363479 524231 363513
rect 524265 363479 524303 363513
rect 524337 363479 524375 363513
rect 524409 363479 524447 363513
rect 524481 363479 524519 363513
rect 524553 363479 524591 363513
rect 524625 363479 524663 363513
rect 524697 363479 524713 363513
rect 523423 363473 524713 363479
rect 525008 363507 525051 363541
rect 525085 363507 525128 363541
rect 523128 363107 523171 363141
rect 523205 363107 523248 363141
rect 523128 362741 523248 363107
rect 525008 363141 525128 363507
rect 525008 363107 525051 363141
rect 525085 363107 525128 363141
rect 523423 363055 524713 363061
rect 523423 363021 523439 363055
rect 523473 363021 523511 363055
rect 523545 363021 523583 363055
rect 523617 363021 523655 363055
rect 523689 363021 523727 363055
rect 523761 363021 523799 363055
rect 523833 363021 523871 363055
rect 523905 363021 523943 363055
rect 523977 363021 524015 363055
rect 524049 363021 524087 363055
rect 524121 363021 524159 363055
rect 524193 363021 524231 363055
rect 524265 363021 524303 363055
rect 524337 363021 524375 363055
rect 524409 363021 524447 363055
rect 524481 363021 524519 363055
rect 524553 363021 524591 363055
rect 524625 363021 524663 363055
rect 524697 363021 524713 363055
rect 523423 363015 524713 363021
rect 523128 362707 523171 362741
rect 523205 362707 523248 362741
rect 523128 361476 523248 362707
rect 525008 362741 525128 363107
rect 525008 362707 525051 362741
rect 525085 362707 525128 362741
rect 523423 362597 524713 362603
rect 523423 362563 523439 362597
rect 523473 362563 523511 362597
rect 523545 362563 523583 362597
rect 523617 362563 523655 362597
rect 523689 362563 523727 362597
rect 523761 362563 523799 362597
rect 523833 362563 523871 362597
rect 523905 362563 523943 362597
rect 523977 362563 524015 362597
rect 524049 362563 524087 362597
rect 524121 362563 524159 362597
rect 524193 362563 524231 362597
rect 524265 362563 524303 362597
rect 524337 362563 524375 362597
rect 524409 362563 524447 362597
rect 524481 362563 524519 362597
rect 524553 362563 524591 362597
rect 524625 362563 524663 362597
rect 524697 362563 524713 362597
rect 523423 362557 524713 362563
rect 523128 359888 523130 361476
rect 523246 359888 523248 361476
rect 523128 359866 523248 359888
rect 521248 357440 521250 359028
rect 521366 357440 521368 359028
rect 521248 357418 521368 357440
rect 525008 359028 525128 362707
rect 526888 411584 527008 411606
rect 526888 409996 526890 411584
rect 527006 409996 527008 411584
rect 526888 370909 527008 409996
rect 526888 370875 526931 370909
rect 526965 370875 527008 370909
rect 526888 370709 527008 370875
rect 527187 371073 527749 371081
rect 527187 370762 527199 371073
rect 526888 370675 526931 370709
rect 526965 370675 527008 370709
rect 526888 370509 527008 370675
rect 526888 370475 526931 370509
rect 526965 370475 527008 370509
rect 526888 370309 527008 370475
rect 526888 370275 526931 370309
rect 526965 370275 527008 370309
rect 526888 370109 527008 370275
rect 526888 370075 526931 370109
rect 526965 370075 527008 370109
rect 526888 369909 527008 370075
rect 526888 369875 526931 369909
rect 526965 369875 527008 369909
rect 526888 369709 527008 369875
rect 526888 369675 526931 369709
rect 526965 369675 527008 369709
rect 526888 369509 527008 369675
rect 526888 369475 526931 369509
rect 526965 369475 527008 369509
rect 526888 369309 527008 369475
rect 526888 369275 526931 369309
rect 526965 369275 527008 369309
rect 526888 369109 527008 369275
rect 526888 369075 526931 369109
rect 526965 369075 527008 369109
rect 526888 368909 527008 369075
rect 526888 368875 526931 368909
rect 526965 368875 527008 368909
rect 526888 368165 527008 368875
rect 526888 368131 526931 368165
rect 526965 368131 527008 368165
rect 526888 367965 527008 368131
rect 526888 367931 526931 367965
rect 526965 367931 527008 367965
rect 526888 367765 527008 367931
rect 526888 367731 526931 367765
rect 526965 367731 527008 367765
rect 526888 367565 527008 367731
rect 526888 367531 526931 367565
rect 526965 367531 527008 367565
rect 526888 367365 527008 367531
rect 526888 367331 526931 367365
rect 526965 367331 527008 367365
rect 526888 367165 527008 367331
rect 526888 367131 526931 367165
rect 526965 367131 527008 367165
rect 526888 366965 527008 367131
rect 526888 366931 526931 366965
rect 526965 366931 527008 366965
rect 526888 366765 527008 366931
rect 526888 366731 526931 366765
rect 526965 366731 527008 366765
rect 526888 366565 527008 366731
rect 526888 366531 526931 366565
rect 526965 366531 527008 366565
rect 526888 366365 527008 366531
rect 526888 366331 526931 366365
rect 526965 366331 527008 366365
rect 526888 366165 527008 366331
rect 526888 366131 526931 366165
rect 526965 366131 527008 366165
rect 526888 365421 527008 366131
rect 527052 370734 527199 370762
rect 527052 365904 527080 370734
rect 527187 370679 527199 370734
rect 527737 370679 527749 371073
rect 527187 370671 527749 370679
rect 528147 371073 528709 371081
rect 528147 370679 528159 371073
rect 528697 370679 528709 371073
rect 528147 370671 528196 370679
rect 528248 370671 528709 370679
rect 528768 370909 528888 412444
rect 532528 414032 532648 414054
rect 532528 412444 532530 414032
rect 532646 412444 532648 414032
rect 528768 370875 528811 370909
rect 528845 370875 528888 370909
rect 528768 370709 528888 370875
rect 528768 370675 528811 370709
rect 528845 370675 528888 370709
rect 528196 370624 528248 370630
rect 527176 370590 527228 370596
rect 527120 370550 527176 370578
rect 527040 365898 527092 365904
rect 527120 365886 527148 370550
rect 527176 370532 527228 370538
rect 528768 370509 528888 370675
rect 528768 370475 528811 370509
rect 528845 370475 528888 370509
rect 528768 370309 528888 370475
rect 528768 370275 528811 370309
rect 528845 370275 528888 370309
rect 528768 370109 528888 370275
rect 528768 370075 528811 370109
rect 528845 370075 528888 370109
rect 528768 369909 528888 370075
rect 528768 369875 528811 369909
rect 528845 369875 528888 369909
rect 528768 369709 528888 369875
rect 528768 369675 528811 369709
rect 528845 369675 528888 369709
rect 528768 369509 528888 369675
rect 528768 369475 528811 369509
rect 528845 369475 528888 369509
rect 528768 369309 528888 369475
rect 528768 369275 528811 369309
rect 528845 369275 528888 369309
rect 528768 369109 528888 369275
rect 527749 369073 528713 369084
rect 527187 369066 528713 369073
rect 527187 368672 527199 369066
rect 527737 368672 528159 369066
rect 528697 368672 528713 369066
rect 527187 368663 528713 368672
rect 527749 368652 528713 368663
rect 528768 369075 528811 369109
rect 528845 369075 528888 369109
rect 528768 368909 528888 369075
rect 528768 368875 528811 368909
rect 528845 368875 528888 368909
rect 527187 368329 527749 368337
rect 527187 367935 527199 368329
rect 527737 368296 527749 368329
rect 528147 368329 528709 368337
rect 527737 368290 527772 368296
rect 527737 368232 527772 368238
rect 527737 367935 527749 368232
rect 527187 367927 527749 367935
rect 528147 367935 528159 368329
rect 528697 368020 528709 368329
rect 528768 368165 528888 368875
rect 528768 368131 528811 368165
rect 528845 368131 528888 368165
rect 528697 368014 528724 368020
rect 528697 367956 528724 367962
rect 528768 367965 528888 368131
rect 528697 367935 528709 367956
rect 528147 367927 528709 367935
rect 528768 367931 528811 367965
rect 528845 367931 528888 367965
rect 528768 367765 528888 367931
rect 528768 367731 528811 367765
rect 528845 367731 528888 367765
rect 528768 367565 528888 367731
rect 528768 367531 528811 367565
rect 528845 367531 528888 367565
rect 528768 367365 528888 367531
rect 528768 367331 528811 367365
rect 528845 367331 528888 367365
rect 528768 367165 528888 367331
rect 528768 367131 528811 367165
rect 528845 367131 528888 367165
rect 528768 366965 528888 367131
rect 528768 366931 528811 366965
rect 528845 366931 528888 366965
rect 528768 366765 528888 366931
rect 528768 366731 528811 366765
rect 528845 366731 528888 366765
rect 528768 366565 528888 366731
rect 528768 366531 528811 366565
rect 528845 366531 528888 366565
rect 528768 366365 528888 366531
rect 527749 366329 528713 366340
rect 527187 366322 528713 366329
rect 527187 365928 527199 366322
rect 527737 365928 528159 366322
rect 528697 365928 528713 366322
rect 527187 365919 528713 365928
rect 527749 365908 528713 365919
rect 528768 366331 528811 366365
rect 528845 366331 528888 366365
rect 528768 366165 528888 366331
rect 528768 366131 528811 366165
rect 528845 366131 528888 366165
rect 527120 365858 527216 365886
rect 527040 365840 527092 365846
rect 527188 365593 527216 365858
rect 526888 365387 526931 365421
rect 526965 365387 527008 365421
rect 526888 365221 527008 365387
rect 526888 365187 526931 365221
rect 526965 365187 527008 365221
rect 526888 365021 527008 365187
rect 527187 365585 527749 365593
rect 527187 365191 527199 365585
rect 527737 365191 527749 365585
rect 527187 365183 527749 365191
rect 528147 365585 528709 365593
rect 528147 365191 528159 365585
rect 528697 365444 528709 365585
rect 528697 365438 528724 365444
rect 528697 365380 528724 365386
rect 528768 365421 528888 366131
rect 528768 365387 528811 365421
rect 528845 365387 528888 365421
rect 528697 365191 528709 365380
rect 528147 365183 528709 365191
rect 528768 365221 528888 365387
rect 528768 365187 528811 365221
rect 528845 365187 528888 365221
rect 526888 364987 526931 365021
rect 526965 364987 527008 365021
rect 526888 364821 527008 364987
rect 526888 364787 526931 364821
rect 526965 364787 527008 364821
rect 526888 364621 527008 364787
rect 526888 364587 526931 364621
rect 526965 364587 527008 364621
rect 526888 364421 527008 364587
rect 526888 364387 526931 364421
rect 526965 364387 527008 364421
rect 526888 364221 527008 364387
rect 526888 364187 526931 364221
rect 526965 364187 527008 364221
rect 526888 364021 527008 364187
rect 526888 363987 526931 364021
rect 526965 363987 527008 364021
rect 526888 363821 527008 363987
rect 526888 363787 526931 363821
rect 526965 363787 527008 363821
rect 526888 363621 527008 363787
rect 526888 363587 526931 363621
rect 526965 363587 527008 363621
rect 528768 365021 528888 365187
rect 528768 364987 528811 365021
rect 528845 364987 528888 365021
rect 528768 364821 528888 364987
rect 528768 364787 528811 364821
rect 528845 364787 528888 364821
rect 528768 364621 528888 364787
rect 528768 364587 528811 364621
rect 528845 364587 528888 364621
rect 528768 364421 528888 364587
rect 528768 364387 528811 364421
rect 528845 364387 528888 364421
rect 528768 364221 528888 364387
rect 528768 364187 528811 364221
rect 528845 364187 528888 364221
rect 528768 364021 528888 364187
rect 528768 363987 528811 364021
rect 528845 363987 528888 364021
rect 528768 363821 528888 363987
rect 528768 363787 528811 363821
rect 528845 363787 528888 363821
rect 528768 363621 528888 363787
rect 526888 363421 527008 363587
rect 527749 363585 528713 363596
rect 526888 363387 526931 363421
rect 526965 363387 527008 363421
rect 526888 361476 527008 363387
rect 527187 363578 528713 363585
rect 527187 363184 527199 363578
rect 527737 363184 528159 363578
rect 528697 363184 528713 363578
rect 527187 363175 528713 363184
rect 527749 363164 528713 363175
rect 528768 363587 528811 363621
rect 528845 363587 528888 363621
rect 528768 363421 528888 363587
rect 528768 363387 528811 363421
rect 528845 363387 528888 363421
rect 526888 359888 526890 361476
rect 527006 359888 527008 361476
rect 526888 359866 527008 359888
rect 525008 357440 525010 359028
rect 525126 357440 525128 359028
rect 525008 357418 525128 357440
rect 528768 359028 528888 363387
rect 530648 411584 530768 411606
rect 530648 409996 530650 411584
rect 530766 409996 530768 411584
rect 530648 371007 530768 409996
rect 530648 370973 530691 371007
rect 530725 370973 530768 371007
rect 530648 370807 530768 370973
rect 530648 370773 530691 370807
rect 530725 370773 530768 370807
rect 530648 370607 530768 370773
rect 530947 371171 531509 371179
rect 530947 370777 530959 371171
rect 531497 370777 531509 371171
rect 530947 370769 531509 370777
rect 531907 371171 532469 371179
rect 531907 370777 531919 371171
rect 532457 370777 532469 371171
rect 531907 370769 532469 370777
rect 532528 371007 532648 412444
rect 536288 414032 536408 414054
rect 536288 412444 536290 414032
rect 536406 412444 536408 414032
rect 532528 370973 532571 371007
rect 532605 370973 532648 371007
rect 532528 370807 532648 370973
rect 532528 370773 532571 370807
rect 532605 370773 532648 370807
rect 530648 370573 530691 370607
rect 530725 370573 530768 370607
rect 530648 370407 530768 370573
rect 530648 370373 530691 370407
rect 530725 370373 530768 370407
rect 530648 370207 530768 370373
rect 530648 370173 530691 370207
rect 530725 370173 530768 370207
rect 530648 370007 530768 370173
rect 530848 370222 530900 370228
rect 530848 370164 530900 370170
rect 530648 369973 530691 370007
rect 530725 369973 530768 370007
rect 530648 369807 530768 369973
rect 530648 369773 530691 369807
rect 530725 369773 530768 369807
rect 530648 369607 530768 369773
rect 530648 369573 530691 369607
rect 530725 369573 530768 369607
rect 530648 369407 530768 369573
rect 530648 369373 530691 369407
rect 530725 369373 530768 369407
rect 530648 369207 530768 369373
rect 530648 369173 530691 369207
rect 530725 369173 530768 369207
rect 530648 369007 530768 369173
rect 530648 368973 530691 369007
rect 530725 368973 530768 369007
rect 530648 368263 530768 368973
rect 530860 368646 530888 370164
rect 532424 369308 532452 370769
rect 532528 370607 532648 370773
rect 532528 370573 532571 370607
rect 532605 370573 532648 370607
rect 532528 370407 532648 370573
rect 532528 370373 532571 370407
rect 532605 370373 532648 370407
rect 532528 370207 532648 370373
rect 532528 370173 532571 370207
rect 532605 370173 532648 370207
rect 532528 370007 532648 370173
rect 532528 369973 532571 370007
rect 532605 369973 532648 370007
rect 532528 369807 532648 369973
rect 532528 369773 532571 369807
rect 532605 369773 532648 369807
rect 532528 369607 532648 369773
rect 532528 369573 532571 369607
rect 532605 369573 532648 369607
rect 532528 369407 532648 369573
rect 532528 369373 532571 369407
rect 532605 369373 532648 369407
rect 532412 369302 532464 369308
rect 532412 369244 532464 369250
rect 532528 369207 532648 369373
rect 534408 411584 534528 411606
rect 534408 409996 534410 411584
rect 534526 409996 534528 411584
rect 534408 370223 534528 409996
rect 534408 370189 534451 370223
rect 534485 370189 534528 370223
rect 534408 370023 534528 370189
rect 534408 369989 534451 370023
rect 534485 369989 534528 370023
rect 534408 369823 534528 369989
rect 534707 370387 535269 370395
rect 534707 369993 534719 370387
rect 535257 369993 535269 370387
rect 534707 369985 535269 369993
rect 535667 370387 536229 370395
rect 535667 370222 535679 370387
rect 535667 370170 535676 370222
rect 535667 369993 535679 370170
rect 536217 369993 536229 370387
rect 535667 369985 536229 369993
rect 536288 370223 536408 412444
rect 566254 405476 566462 405488
rect 566246 405258 566256 405476
rect 566462 405258 566472 405476
rect 580076 405402 580180 405420
rect 580064 405292 580074 405402
rect 580182 405292 580192 405402
rect 560592 404708 565906 404738
rect 560592 404648 560860 404708
rect 560920 404648 561060 404708
rect 561120 404648 561260 404708
rect 561320 404648 561460 404708
rect 561520 404648 561660 404708
rect 561720 404648 561860 404708
rect 561920 404648 562060 404708
rect 562120 404648 562260 404708
rect 562320 404648 562460 404708
rect 562520 404648 562660 404708
rect 562720 404648 562860 404708
rect 562920 404648 563060 404708
rect 563120 404648 563260 404708
rect 563320 404648 563460 404708
rect 563520 404648 563660 404708
rect 563720 404648 563860 404708
rect 563920 404648 564060 404708
rect 564120 404648 564260 404708
rect 564320 404648 564460 404708
rect 564520 404648 564660 404708
rect 564720 404648 564860 404708
rect 564920 404648 565060 404708
rect 565120 404648 565260 404708
rect 565320 404648 565460 404708
rect 565520 404648 565660 404708
rect 565720 404648 565906 404708
rect 560592 404618 565906 404648
rect 560695 404286 560741 404298
rect 559722 403368 559976 403390
rect 559722 403192 559736 403368
rect 559926 403310 559976 403368
rect 560695 403310 560701 404286
rect 560735 403310 560741 404286
rect 559926 403286 560498 403310
rect 560695 403298 560741 403310
rect 560953 404286 560999 404298
rect 560953 403310 560959 404286
rect 560993 403310 560999 404286
rect 560953 403298 560999 403310
rect 561211 404286 561257 404298
rect 561211 403310 561217 404286
rect 561251 403310 561257 404286
rect 561211 403298 561257 403310
rect 561469 404286 561515 404298
rect 561469 403310 561475 404286
rect 561509 403310 561515 404286
rect 561469 403298 561515 403310
rect 561727 404286 561773 404298
rect 561727 403310 561733 404286
rect 561767 403310 561773 404286
rect 561727 403298 561773 403310
rect 561985 404286 562031 404298
rect 561985 403310 561991 404286
rect 562025 403310 562031 404286
rect 561985 403298 562031 403310
rect 562243 404286 562289 404298
rect 562243 403310 562249 404286
rect 562283 403310 562289 404286
rect 562243 403298 562289 403310
rect 562501 404286 562547 404298
rect 562501 403310 562507 404286
rect 562541 403310 562547 404286
rect 562501 403298 562547 403310
rect 562759 404286 562805 404298
rect 562759 403310 562765 404286
rect 562799 403310 562805 404286
rect 562759 403298 562805 403310
rect 563017 404286 563063 404298
rect 563017 403310 563023 404286
rect 563057 403310 563063 404286
rect 563017 403298 563063 403310
rect 563275 404286 563321 404298
rect 563275 403310 563281 404286
rect 563315 403310 563321 404286
rect 563275 403298 563321 403310
rect 563533 404286 563579 404298
rect 563533 403310 563539 404286
rect 563573 403310 563579 404286
rect 563533 403298 563579 403310
rect 563791 404286 563837 404298
rect 563791 403310 563797 404286
rect 563831 403310 563837 404286
rect 563791 403298 563837 403310
rect 564049 404286 564095 404298
rect 564049 403310 564055 404286
rect 564089 403310 564095 404286
rect 564049 403298 564095 403310
rect 564307 404286 564353 404298
rect 564307 403310 564313 404286
rect 564347 403310 564353 404286
rect 564307 403298 564353 403310
rect 564565 404286 564611 404298
rect 564565 403310 564571 404286
rect 564605 403310 564611 404286
rect 564565 403298 564611 403310
rect 564823 404286 564869 404298
rect 564823 403310 564829 404286
rect 564863 403310 564869 404286
rect 564823 403298 564869 403310
rect 565081 404286 565127 404298
rect 565081 403310 565087 404286
rect 565121 403310 565127 404286
rect 565081 403298 565127 403310
rect 565339 404286 565385 404298
rect 565339 403310 565345 404286
rect 565379 403310 565385 404286
rect 565339 403298 565385 403310
rect 565597 404286 565643 404298
rect 565597 403310 565603 404286
rect 565637 403310 565643 404286
rect 565597 403298 565643 403310
rect 565855 404286 565901 404298
rect 565855 403310 565861 404286
rect 565895 403310 565901 404286
rect 566254 403370 566462 405258
rect 574448 404748 579834 404778
rect 574448 404688 574506 404748
rect 574566 404688 574706 404748
rect 574766 404688 574906 404748
rect 574966 404688 575106 404748
rect 575166 404688 575306 404748
rect 575366 404688 575506 404748
rect 575566 404688 575706 404748
rect 575766 404688 575906 404748
rect 575966 404688 576106 404748
rect 576166 404688 576306 404748
rect 576366 404688 576506 404748
rect 576566 404688 576706 404748
rect 576766 404688 576906 404748
rect 576966 404688 577106 404748
rect 577166 404688 577306 404748
rect 577366 404688 577506 404748
rect 577566 404688 577706 404748
rect 577766 404688 577906 404748
rect 577966 404688 578106 404748
rect 578166 404688 578306 404748
rect 578366 404688 578506 404748
rect 578566 404688 578706 404748
rect 578766 404688 578906 404748
rect 578966 404688 579106 404748
rect 579166 404688 579306 404748
rect 579366 404688 579506 404748
rect 579566 404688 579834 404748
rect 574448 404658 579834 404688
rect 565855 403298 565901 403310
rect 566070 403340 566462 403370
rect 574489 404326 574535 404338
rect 559926 403192 560322 403286
rect 559722 403178 560322 403192
rect 560482 403178 560498 403286
rect 559722 403162 560498 403178
rect 566070 403190 566084 403340
rect 566216 403190 566462 403340
rect 566070 403162 566462 403190
rect 573509 403312 574144 403353
rect 574489 403350 574495 404326
rect 574529 403350 574535 404326
rect 574489 403338 574535 403350
rect 574747 404326 574793 404338
rect 574747 403350 574753 404326
rect 574787 403350 574793 404326
rect 574747 403338 574793 403350
rect 575005 404326 575051 404338
rect 575005 403350 575011 404326
rect 575045 403350 575051 404326
rect 575005 403338 575051 403350
rect 575263 404326 575309 404338
rect 575263 403350 575269 404326
rect 575303 403350 575309 404326
rect 575263 403338 575309 403350
rect 575521 404326 575567 404338
rect 575521 403350 575527 404326
rect 575561 403350 575567 404326
rect 575521 403338 575567 403350
rect 575779 404326 575825 404338
rect 575779 403350 575785 404326
rect 575819 403350 575825 404326
rect 575779 403338 575825 403350
rect 576037 404326 576083 404338
rect 576037 403350 576043 404326
rect 576077 403350 576083 404326
rect 576037 403338 576083 403350
rect 576295 404326 576341 404338
rect 576295 403350 576301 404326
rect 576335 403350 576341 404326
rect 576295 403338 576341 403350
rect 576553 404326 576599 404338
rect 576553 403350 576559 404326
rect 576593 403350 576599 404326
rect 576553 403338 576599 403350
rect 576811 404326 576857 404338
rect 576811 403350 576817 404326
rect 576851 403350 576857 404326
rect 576811 403338 576857 403350
rect 577069 404326 577115 404338
rect 577069 403350 577075 404326
rect 577109 403350 577115 404326
rect 577069 403338 577115 403350
rect 577327 404326 577373 404338
rect 577327 403350 577333 404326
rect 577367 403350 577373 404326
rect 577327 403338 577373 403350
rect 577585 404326 577631 404338
rect 577585 403350 577591 404326
rect 577625 403350 577631 404326
rect 577585 403338 577631 403350
rect 577843 404326 577889 404338
rect 577843 403350 577849 404326
rect 577883 403350 577889 404326
rect 577843 403338 577889 403350
rect 578101 404326 578147 404338
rect 578101 403350 578107 404326
rect 578141 403350 578147 404326
rect 578101 403338 578147 403350
rect 578359 404326 578405 404338
rect 578359 403350 578365 404326
rect 578399 403350 578405 404326
rect 578359 403338 578405 403350
rect 578617 404326 578663 404338
rect 578617 403350 578623 404326
rect 578657 403350 578663 404326
rect 578617 403338 578663 403350
rect 578875 404326 578921 404338
rect 578875 403350 578881 404326
rect 578915 403350 578921 404326
rect 578875 403338 578921 403350
rect 579133 404326 579179 404338
rect 579133 403350 579139 404326
rect 579173 403350 579179 404326
rect 579133 403338 579179 403350
rect 579391 404326 579437 404338
rect 579391 403350 579397 404326
rect 579431 403350 579437 404326
rect 579391 403338 579437 403350
rect 579649 404326 579695 404338
rect 579649 403350 579655 404326
rect 579689 403350 579695 404326
rect 579649 403338 579695 403350
rect 573509 403107 573538 403312
rect 573510 402980 573538 403107
rect 573888 403120 574144 403312
rect 580076 403254 580180 405292
rect 579808 403242 580180 403254
rect 579808 403154 579820 403242
rect 579910 403154 580180 403242
rect 579808 403150 580180 403154
rect 579808 403148 579922 403150
rect 573888 403108 574312 403120
rect 573888 403004 574212 403108
rect 574304 403004 574312 403108
rect 573888 402992 574312 403004
rect 573888 402980 574196 402992
rect 573510 402956 574196 402980
rect 574448 402868 579834 402898
rect 560592 402828 565906 402858
rect 560592 402768 560860 402828
rect 560920 402768 561060 402828
rect 561120 402768 561260 402828
rect 561320 402768 561460 402828
rect 561520 402768 561660 402828
rect 561720 402768 561860 402828
rect 561920 402768 562060 402828
rect 562120 402768 562260 402828
rect 562320 402768 562460 402828
rect 562520 402768 562660 402828
rect 562720 402768 562860 402828
rect 562920 402768 563060 402828
rect 563120 402768 563260 402828
rect 563320 402768 563460 402828
rect 563520 402768 563660 402828
rect 563720 402768 563860 402828
rect 563920 402768 564060 402828
rect 564120 402768 564260 402828
rect 564320 402768 564460 402828
rect 564520 402768 564660 402828
rect 564720 402768 564860 402828
rect 564920 402768 565060 402828
rect 565120 402768 565260 402828
rect 565320 402768 565460 402828
rect 565520 402768 565660 402828
rect 565720 402768 565906 402828
rect 574448 402808 574506 402868
rect 574566 402808 574706 402868
rect 574766 402808 574906 402868
rect 574966 402808 575106 402868
rect 575166 402808 575306 402868
rect 575366 402808 575506 402868
rect 575566 402808 575706 402868
rect 575766 402808 575906 402868
rect 575966 402808 576106 402868
rect 576166 402808 576306 402868
rect 576366 402808 576506 402868
rect 576566 402808 576706 402868
rect 576766 402808 576906 402868
rect 576966 402808 577106 402868
rect 577166 402808 577306 402868
rect 577366 402808 577506 402868
rect 577566 402808 577706 402868
rect 577766 402808 577906 402868
rect 577966 402808 578106 402868
rect 578166 402808 578306 402868
rect 578366 402808 578506 402868
rect 578566 402808 578706 402868
rect 578766 402808 578906 402868
rect 578966 402808 579106 402868
rect 579166 402808 579306 402868
rect 579366 402808 579506 402868
rect 579566 402808 579834 402868
rect 574448 402778 579834 402808
rect 560592 402738 565906 402768
rect 537512 389450 537564 389456
rect 537512 389392 537564 389398
rect 537524 387432 537552 389392
rect 537512 387426 537564 387432
rect 537512 387368 537564 387374
rect 536288 370189 536331 370223
rect 536365 370189 536408 370223
rect 536288 370023 536408 370189
rect 536288 369989 536331 370023
rect 536365 369989 536408 370023
rect 534408 369789 534451 369823
rect 534485 369789 534528 369823
rect 534408 369623 534528 369789
rect 534408 369589 534451 369623
rect 534485 369589 534528 369623
rect 534408 369423 534528 369589
rect 534408 369389 534451 369423
rect 534485 369389 534528 369423
rect 532684 369302 532736 369308
rect 532684 369244 532736 369250
rect 531509 369171 532473 369182
rect 530947 369164 532473 369171
rect 530947 368770 530959 369164
rect 531497 368770 531919 369164
rect 532457 368770 532473 369164
rect 530947 368761 532473 368770
rect 531509 368750 532473 368761
rect 532528 369173 532571 369207
rect 532605 369173 532648 369207
rect 532528 369007 532648 369173
rect 532528 368973 532571 369007
rect 532605 368973 532648 369007
rect 530860 368618 531024 368646
rect 530996 368435 531024 368618
rect 530648 368229 530691 368263
rect 530725 368229 530768 368263
rect 530648 368063 530768 368229
rect 530648 368029 530691 368063
rect 530725 368029 530768 368063
rect 530648 367863 530768 368029
rect 530947 368427 531509 368435
rect 530947 368033 530959 368427
rect 531497 368033 531509 368427
rect 530947 368025 531509 368033
rect 531907 368427 532469 368435
rect 531907 368033 531919 368427
rect 532457 368033 532469 368427
rect 531907 368025 532469 368033
rect 532528 368263 532648 368973
rect 532528 368229 532571 368263
rect 532605 368229 532648 368263
rect 532528 368063 532648 368229
rect 532528 368029 532571 368063
rect 532605 368029 532648 368063
rect 530848 368014 530900 368020
rect 530848 367956 530900 367962
rect 530648 367829 530691 367863
rect 530725 367829 530768 367863
rect 530648 367663 530768 367829
rect 530648 367629 530691 367663
rect 530725 367629 530768 367663
rect 530648 367463 530768 367629
rect 530648 367429 530691 367463
rect 530725 367429 530768 367463
rect 530648 367263 530768 367429
rect 530648 367229 530691 367263
rect 530725 367229 530768 367263
rect 530648 367063 530768 367229
rect 530648 367029 530691 367063
rect 530725 367029 530768 367063
rect 530648 366863 530768 367029
rect 530648 366829 530691 366863
rect 530725 366829 530768 366863
rect 530648 366663 530768 366829
rect 530648 366629 530691 366663
rect 530725 366629 530768 366663
rect 530648 366463 530768 366629
rect 530648 366429 530691 366463
rect 530725 366429 530768 366463
rect 530648 366263 530768 366429
rect 530648 366229 530691 366263
rect 530725 366229 530768 366263
rect 530648 365519 530768 366229
rect 530860 365978 530888 367956
rect 532528 367863 532648 368029
rect 532528 367829 532571 367863
rect 532605 367829 532648 367863
rect 532528 367663 532648 367829
rect 532528 367629 532571 367663
rect 532605 367629 532648 367663
rect 532528 367463 532648 367629
rect 532528 367429 532571 367463
rect 532605 367429 532648 367463
rect 532528 367263 532648 367429
rect 532528 367229 532571 367263
rect 532605 367229 532648 367263
rect 532528 367063 532648 367229
rect 532528 367029 532571 367063
rect 532605 367029 532648 367063
rect 532528 366863 532648 367029
rect 532528 366829 532571 366863
rect 532605 366829 532648 366863
rect 532528 366663 532648 366829
rect 532528 366629 532571 366663
rect 532605 366629 532648 366663
rect 532528 366463 532648 366629
rect 531509 366427 532473 366438
rect 530947 366420 532473 366427
rect 530947 366026 530959 366420
rect 531497 366026 531919 366420
rect 532457 366026 532473 366420
rect 530947 366017 532473 366026
rect 531509 366006 532473 366017
rect 532528 366429 532571 366463
rect 532605 366429 532648 366463
rect 532528 366263 532648 366429
rect 532528 366229 532571 366263
rect 532605 366229 532648 366263
rect 530860 365950 531024 365978
rect 530996 365691 531024 365950
rect 531936 365898 531988 365904
rect 531936 365840 531988 365846
rect 531948 365691 531976 365840
rect 530648 365485 530691 365519
rect 530725 365485 530768 365519
rect 530648 365319 530768 365485
rect 530648 365285 530691 365319
rect 530725 365285 530768 365319
rect 530648 365119 530768 365285
rect 530947 365683 531509 365691
rect 530947 365289 530959 365683
rect 531497 365289 531509 365683
rect 530947 365281 531509 365289
rect 531907 365683 532469 365691
rect 531907 365289 531919 365683
rect 532457 365289 532469 365683
rect 531907 365281 532469 365289
rect 532528 365519 532648 366229
rect 532528 365485 532571 365519
rect 532605 365485 532648 365519
rect 532528 365319 532648 365485
rect 532528 365285 532571 365319
rect 532605 365285 532648 365319
rect 530648 365085 530691 365119
rect 530725 365085 530768 365119
rect 530648 364919 530768 365085
rect 530648 364885 530691 364919
rect 530725 364885 530768 364919
rect 530648 364719 530768 364885
rect 530648 364685 530691 364719
rect 530725 364685 530768 364719
rect 530648 364519 530768 364685
rect 530648 364485 530691 364519
rect 530725 364485 530768 364519
rect 530648 364319 530768 364485
rect 530648 364285 530691 364319
rect 530725 364285 530768 364319
rect 530648 364119 530768 364285
rect 530648 364085 530691 364119
rect 530725 364085 530768 364119
rect 530648 363919 530768 364085
rect 530648 363885 530691 363919
rect 530725 363885 530768 363919
rect 530648 363719 530768 363885
rect 530648 363685 530691 363719
rect 530725 363685 530768 363719
rect 532528 365119 532648 365285
rect 532528 365085 532571 365119
rect 532605 365085 532648 365119
rect 532528 364919 532648 365085
rect 532696 365076 532724 369244
rect 534408 369223 534528 369389
rect 534408 369189 534451 369223
rect 534485 369189 534528 369223
rect 534408 369023 534528 369189
rect 534408 368989 534451 369023
rect 534485 368989 534528 369023
rect 534408 368823 534528 368989
rect 534408 368789 534451 368823
rect 534485 368789 534528 368823
rect 534408 368623 534528 368789
rect 534408 368589 534451 368623
rect 534485 368589 534528 368623
rect 534408 368423 534528 368589
rect 534736 368462 534764 369985
rect 534408 368389 534451 368423
rect 534485 368389 534528 368423
rect 534408 368223 534528 368389
rect 534408 368189 534451 368223
rect 534485 368189 534528 368223
rect 534408 367479 534528 368189
rect 534408 367445 534451 367479
rect 534485 367445 534528 367479
rect 534408 367279 534528 367445
rect 534408 367245 534451 367279
rect 534485 367245 534528 367279
rect 534408 367079 534528 367245
rect 534408 367045 534451 367079
rect 534485 367045 534528 367079
rect 534408 366879 534528 367045
rect 534408 366845 534451 366879
rect 534485 366845 534528 366879
rect 534408 366679 534528 366845
rect 534408 366645 534451 366679
rect 534485 366645 534528 366679
rect 534408 366479 534528 366645
rect 534408 366445 534451 366479
rect 534485 366445 534528 366479
rect 534408 366279 534528 366445
rect 534408 366245 534451 366279
rect 534485 366245 534528 366279
rect 534408 366079 534528 366245
rect 534408 366045 534451 366079
rect 534485 366045 534528 366079
rect 534408 365879 534528 366045
rect 534408 365845 534451 365879
rect 534485 365845 534528 365879
rect 534408 365679 534528 365845
rect 534408 365645 534451 365679
rect 534485 365645 534528 365679
rect 534408 365479 534528 365645
rect 534408 365445 534451 365479
rect 534485 365445 534528 365479
rect 532684 365070 532736 365076
rect 532684 365012 532736 365018
rect 532528 364885 532571 364919
rect 532605 364885 532648 364919
rect 532528 364719 532648 364885
rect 532528 364685 532571 364719
rect 532605 364685 532648 364719
rect 532528 364519 532648 364685
rect 532528 364485 532571 364519
rect 532605 364485 532648 364519
rect 532528 364319 532648 364485
rect 532528 364285 532571 364319
rect 532605 364285 532648 364319
rect 532528 364119 532648 364285
rect 532528 364085 532571 364119
rect 532605 364085 532648 364119
rect 532528 363919 532648 364085
rect 532528 363885 532571 363919
rect 532605 363885 532648 363919
rect 532528 363719 532648 363885
rect 530648 363519 530768 363685
rect 531509 363683 532473 363694
rect 530648 363485 530691 363519
rect 530725 363485 530768 363519
rect 530648 361476 530768 363485
rect 530947 363676 532473 363683
rect 530947 363282 530959 363676
rect 531497 363282 531919 363676
rect 532457 363282 532473 363676
rect 530947 363273 532473 363282
rect 531509 363262 532473 363273
rect 532528 363685 532571 363719
rect 532605 363685 532648 363719
rect 532528 363519 532648 363685
rect 532528 363485 532571 363519
rect 532605 363485 532648 363519
rect 530648 359888 530650 361476
rect 530766 359888 530768 361476
rect 530648 359866 530768 359888
rect 528768 357440 528770 359028
rect 528886 357440 528888 359028
rect 528768 357418 528888 357440
rect 532528 359028 532648 363485
rect 534408 364735 534528 365445
rect 534600 368434 534764 368462
rect 536288 369823 536408 369989
rect 536288 369789 536331 369823
rect 536365 369789 536408 369823
rect 536288 369623 536408 369789
rect 536288 369589 536331 369623
rect 536365 369589 536408 369623
rect 536288 369423 536408 369589
rect 536288 369389 536331 369423
rect 536365 369389 536408 369423
rect 536288 369223 536408 369389
rect 536288 369189 536331 369223
rect 536365 369189 536408 369223
rect 536288 369023 536408 369189
rect 536288 368989 536331 369023
rect 536365 368989 536408 369023
rect 536288 368823 536408 368989
rect 536288 368789 536331 368823
rect 536365 368789 536408 368823
rect 536288 368623 536408 368789
rect 536288 368589 536331 368623
rect 536365 368589 536408 368623
rect 534600 365168 534628 368434
rect 536288 368423 536408 368589
rect 535269 368387 536233 368398
rect 534707 368380 536233 368387
rect 534707 367986 534719 368380
rect 535257 367986 535679 368380
rect 536217 367986 536233 368380
rect 534707 367977 536233 367986
rect 535269 367966 536233 367977
rect 536288 368389 536331 368423
rect 536365 368389 536408 368423
rect 536288 368223 536408 368389
rect 536288 368189 536331 368223
rect 536365 368189 536408 368223
rect 534707 367643 535269 367651
rect 534707 367249 534719 367643
rect 535257 367249 535269 367643
rect 534707 367241 535269 367249
rect 535667 367643 536229 367651
rect 535667 367249 535679 367643
rect 536217 367634 536229 367643
rect 536288 367634 536408 368189
rect 536217 367606 536408 367634
rect 536217 367249 536229 367606
rect 535667 367241 536229 367249
rect 536288 367479 536408 367606
rect 536288 367445 536331 367479
rect 536365 367445 536408 367479
rect 536288 367279 536408 367445
rect 536288 367245 536331 367279
rect 536365 367245 536408 367279
rect 534736 365812 534764 367241
rect 536288 367079 536408 367245
rect 536288 367045 536331 367079
rect 536365 367045 536408 367079
rect 536288 366879 536408 367045
rect 536288 366845 536331 366879
rect 536365 366845 536408 366879
rect 536288 366679 536408 366845
rect 536288 366645 536331 366679
rect 536365 366645 536408 366679
rect 536288 366479 536408 366645
rect 536288 366445 536331 366479
rect 536365 366445 536408 366479
rect 536288 366279 536408 366445
rect 536288 366245 536331 366279
rect 536365 366245 536408 366279
rect 536288 366079 536408 366245
rect 536288 366045 536331 366079
rect 536365 366045 536408 366079
rect 536288 365879 536408 366045
rect 536288 365845 536331 365879
rect 536365 365845 536408 365879
rect 534724 365806 534776 365812
rect 534724 365748 534776 365754
rect 536288 365679 536408 365845
rect 535269 365643 536233 365654
rect 534707 365636 536233 365643
rect 534707 365242 534719 365636
rect 535257 365242 535679 365636
rect 536217 365242 536233 365636
rect 534707 365233 536233 365242
rect 535269 365222 536233 365233
rect 536288 365645 536331 365679
rect 536365 365645 536408 365679
rect 536288 365479 536408 365645
rect 536288 365445 536331 365479
rect 536365 365445 536408 365479
rect 534588 365162 534640 365168
rect 534588 365104 534640 365110
rect 535676 365162 535728 365168
rect 535676 365104 535728 365110
rect 534724 365070 534776 365076
rect 534724 365012 534776 365018
rect 534736 364907 534764 365012
rect 535688 364907 535716 365104
rect 534408 364701 534451 364735
rect 534485 364701 534528 364735
rect 534408 364535 534528 364701
rect 534408 364501 534451 364535
rect 534485 364501 534528 364535
rect 534408 364335 534528 364501
rect 534707 364899 535269 364907
rect 534707 364505 534719 364899
rect 535257 364505 535269 364899
rect 534707 364497 535269 364505
rect 535667 364899 536229 364907
rect 535667 364505 535679 364899
rect 536217 364505 536229 364899
rect 535667 364497 536229 364505
rect 536288 364735 536408 365445
rect 536288 364701 536331 364735
rect 536365 364701 536408 364735
rect 536288 364535 536408 364701
rect 536288 364501 536331 364535
rect 536365 364501 536408 364535
rect 534408 364301 534451 364335
rect 534485 364301 534528 364335
rect 534408 364135 534528 364301
rect 534408 364101 534451 364135
rect 534485 364101 534528 364135
rect 534408 363935 534528 364101
rect 534408 363901 534451 363935
rect 534485 363901 534528 363935
rect 534408 363735 534528 363901
rect 534408 363701 534451 363735
rect 534485 363701 534528 363735
rect 534408 363535 534528 363701
rect 534408 363501 534451 363535
rect 534485 363501 534528 363535
rect 534408 363335 534528 363501
rect 534408 363301 534451 363335
rect 534485 363301 534528 363335
rect 534408 363135 534528 363301
rect 534408 363101 534451 363135
rect 534485 363101 534528 363135
rect 534408 362935 534528 363101
rect 534408 362901 534451 362935
rect 534485 362901 534528 362935
rect 536288 364335 536408 364501
rect 536288 364301 536331 364335
rect 536365 364301 536408 364335
rect 536288 364135 536408 364301
rect 536288 364101 536331 364135
rect 536365 364101 536408 364135
rect 536288 363935 536408 364101
rect 536288 363901 536331 363935
rect 536365 363901 536408 363935
rect 536288 363735 536408 363901
rect 536288 363701 536331 363735
rect 536365 363701 536408 363735
rect 536288 363535 536408 363701
rect 536288 363501 536331 363535
rect 536365 363501 536408 363535
rect 536288 363335 536408 363501
rect 536288 363301 536331 363335
rect 536365 363301 536408 363335
rect 536288 363135 536408 363301
rect 536288 363101 536331 363135
rect 536365 363101 536408 363135
rect 536288 362935 536408 363101
rect 534408 362735 534528 362901
rect 535269 362899 536233 362910
rect 534408 362701 534451 362735
rect 534485 362701 534528 362735
rect 534408 361476 534528 362701
rect 534707 362892 536233 362899
rect 534707 362498 534719 362892
rect 535257 362498 535679 362892
rect 536217 362498 536233 362892
rect 534707 362489 536233 362498
rect 535269 362478 536233 362489
rect 536288 362901 536331 362935
rect 536365 362901 536408 362935
rect 536288 362735 536408 362901
rect 536288 362701 536331 362735
rect 536365 362701 536408 362735
rect 534408 359888 534410 361476
rect 534526 359888 534528 361476
rect 534408 359866 534528 359888
rect 532528 357440 532530 359028
rect 532646 357440 532648 359028
rect 532528 357418 532648 357440
rect 536288 359028 536408 362701
rect 566270 359978 566494 360002
rect 566264 359786 566274 359978
rect 566500 359786 566510 359978
rect 580252 359906 580356 359934
rect 580242 359786 580252 359906
rect 580358 359786 580368 359906
rect 560542 359390 565856 359420
rect 560542 359330 560728 359390
rect 560788 359330 560928 359390
rect 560988 359330 561128 359390
rect 561188 359330 561328 359390
rect 561388 359330 561528 359390
rect 561588 359330 561728 359390
rect 561788 359330 561928 359390
rect 561988 359330 562128 359390
rect 562188 359330 562328 359390
rect 562388 359330 562528 359390
rect 562588 359330 562728 359390
rect 562788 359330 562928 359390
rect 562988 359330 563128 359390
rect 563188 359330 563328 359390
rect 563388 359330 563528 359390
rect 563588 359330 563728 359390
rect 563788 359330 563928 359390
rect 563988 359330 564128 359390
rect 564188 359330 564328 359390
rect 564388 359330 564528 359390
rect 564588 359330 564728 359390
rect 564788 359330 564928 359390
rect 564988 359330 565128 359390
rect 565188 359330 565328 359390
rect 565388 359330 565528 359390
rect 565588 359330 565856 359390
rect 560542 359300 565856 359330
rect 536288 357440 536290 359028
rect 536406 357440 536408 359028
rect 560547 358968 560593 358980
rect 559702 357844 559712 358052
rect 559920 358022 560378 358052
rect 559920 357872 560232 358022
rect 560364 357872 560378 358022
rect 560547 357992 560553 358968
rect 560587 357992 560593 358968
rect 560547 357980 560593 357992
rect 560805 358968 560851 358980
rect 560805 357992 560811 358968
rect 560845 357992 560851 358968
rect 560805 357980 560851 357992
rect 561063 358968 561109 358980
rect 561063 357992 561069 358968
rect 561103 357992 561109 358968
rect 561063 357980 561109 357992
rect 561321 358968 561367 358980
rect 561321 357992 561327 358968
rect 561361 357992 561367 358968
rect 561321 357980 561367 357992
rect 561579 358968 561625 358980
rect 561579 357992 561585 358968
rect 561619 357992 561625 358968
rect 561579 357980 561625 357992
rect 561837 358968 561883 358980
rect 561837 357992 561843 358968
rect 561877 357992 561883 358968
rect 561837 357980 561883 357992
rect 562095 358968 562141 358980
rect 562095 357992 562101 358968
rect 562135 357992 562141 358968
rect 562095 357980 562141 357992
rect 562353 358968 562399 358980
rect 562353 357992 562359 358968
rect 562393 357992 562399 358968
rect 562353 357980 562399 357992
rect 562611 358968 562657 358980
rect 562611 357992 562617 358968
rect 562651 357992 562657 358968
rect 562611 357980 562657 357992
rect 562869 358968 562915 358980
rect 562869 357992 562875 358968
rect 562909 357992 562915 358968
rect 562869 357980 562915 357992
rect 563127 358968 563173 358980
rect 563127 357992 563133 358968
rect 563167 357992 563173 358968
rect 563127 357980 563173 357992
rect 563385 358968 563431 358980
rect 563385 357992 563391 358968
rect 563425 357992 563431 358968
rect 563385 357980 563431 357992
rect 563643 358968 563689 358980
rect 563643 357992 563649 358968
rect 563683 357992 563689 358968
rect 563643 357980 563689 357992
rect 563901 358968 563947 358980
rect 563901 357992 563907 358968
rect 563941 357992 563947 358968
rect 563901 357980 563947 357992
rect 564159 358968 564205 358980
rect 564159 357992 564165 358968
rect 564199 357992 564205 358968
rect 564159 357980 564205 357992
rect 564417 358968 564463 358980
rect 564417 357992 564423 358968
rect 564457 357992 564463 358968
rect 564417 357980 564463 357992
rect 564675 358968 564721 358980
rect 564675 357992 564681 358968
rect 564715 357992 564721 358968
rect 564675 357980 564721 357992
rect 564933 358968 564979 358980
rect 564933 357992 564939 358968
rect 564973 357992 564979 358968
rect 564933 357980 564979 357992
rect 565191 358968 565237 358980
rect 565191 357992 565197 358968
rect 565231 357992 565237 358968
rect 565191 357980 565237 357992
rect 565449 358968 565495 358980
rect 565449 357992 565455 358968
rect 565489 357992 565495 358968
rect 565449 357980 565495 357992
rect 565707 358968 565753 358980
rect 565707 357992 565713 358968
rect 565747 357992 565753 358968
rect 566270 357992 566494 359786
rect 574644 359320 580030 359350
rect 574644 359260 574702 359320
rect 574762 359260 574902 359320
rect 574962 359260 575102 359320
rect 575162 359260 575302 359320
rect 575362 359260 575502 359320
rect 575562 359260 575702 359320
rect 575762 359260 575902 359320
rect 575962 359260 576102 359320
rect 576162 359260 576302 359320
rect 576362 359260 576502 359320
rect 576562 359260 576702 359320
rect 576762 359260 576902 359320
rect 576962 359260 577102 359320
rect 577162 359260 577302 359320
rect 577362 359260 577502 359320
rect 577562 359260 577702 359320
rect 577762 359260 577902 359320
rect 577962 359260 578102 359320
rect 578162 359260 578302 359320
rect 578362 359260 578502 359320
rect 578562 359260 578702 359320
rect 578762 359260 578902 359320
rect 578962 359260 579102 359320
rect 579162 359260 579302 359320
rect 579362 359260 579502 359320
rect 579562 359260 579702 359320
rect 579762 359260 580030 359320
rect 574644 359230 580030 359260
rect 565707 357980 565753 357992
rect 559920 357844 560378 357872
rect 565950 357968 566494 357992
rect 565950 357860 565966 357968
rect 566126 357860 566494 357968
rect 574685 358898 574731 358910
rect 565950 357846 566494 357860
rect 573509 357959 573755 357965
rect 573509 357920 573911 357959
rect 565950 357844 566418 357846
rect 573509 357594 573540 357920
rect 573878 357810 573911 357920
rect 574685 357922 574691 358898
rect 574725 357922 574731 358898
rect 574685 357910 574731 357922
rect 574943 358898 574989 358910
rect 574943 357922 574949 358898
rect 574983 357922 574989 358898
rect 574943 357910 574989 357922
rect 575201 358898 575247 358910
rect 575201 357922 575207 358898
rect 575241 357922 575247 358898
rect 575201 357910 575247 357922
rect 575459 358898 575505 358910
rect 575459 357922 575465 358898
rect 575499 357922 575505 358898
rect 575459 357910 575505 357922
rect 575717 358898 575763 358910
rect 575717 357922 575723 358898
rect 575757 357922 575763 358898
rect 575717 357910 575763 357922
rect 575975 358898 576021 358910
rect 575975 357922 575981 358898
rect 576015 357922 576021 358898
rect 575975 357910 576021 357922
rect 576233 358898 576279 358910
rect 576233 357922 576239 358898
rect 576273 357922 576279 358898
rect 576233 357910 576279 357922
rect 576491 358898 576537 358910
rect 576491 357922 576497 358898
rect 576531 357922 576537 358898
rect 576491 357910 576537 357922
rect 576749 358898 576795 358910
rect 576749 357922 576755 358898
rect 576789 357922 576795 358898
rect 576749 357910 576795 357922
rect 577007 358898 577053 358910
rect 577007 357922 577013 358898
rect 577047 357922 577053 358898
rect 577007 357910 577053 357922
rect 577265 358898 577311 358910
rect 577265 357922 577271 358898
rect 577305 357922 577311 358898
rect 577265 357910 577311 357922
rect 577523 358898 577569 358910
rect 577523 357922 577529 358898
rect 577563 357922 577569 358898
rect 577523 357910 577569 357922
rect 577781 358898 577827 358910
rect 577781 357922 577787 358898
rect 577821 357922 577827 358898
rect 577781 357910 577827 357922
rect 578039 358898 578085 358910
rect 578039 357922 578045 358898
rect 578079 357922 578085 358898
rect 578039 357910 578085 357922
rect 578297 358898 578343 358910
rect 578297 357922 578303 358898
rect 578337 357922 578343 358898
rect 578297 357910 578343 357922
rect 578555 358898 578601 358910
rect 578555 357922 578561 358898
rect 578595 357922 578601 358898
rect 578555 357910 578601 357922
rect 578813 358898 578859 358910
rect 578813 357922 578819 358898
rect 578853 357922 578859 358898
rect 578813 357910 578859 357922
rect 579071 358898 579117 358910
rect 579071 357922 579077 358898
rect 579111 357922 579117 358898
rect 579071 357910 579117 357922
rect 579329 358898 579375 358910
rect 579329 357922 579335 358898
rect 579369 357922 579375 358898
rect 579329 357910 579375 357922
rect 579587 358898 579633 358910
rect 579587 357922 579593 358898
rect 579627 357922 579633 358898
rect 579587 357910 579633 357922
rect 579845 358898 579891 358910
rect 579845 357922 579851 358898
rect 579885 357922 579891 358898
rect 579845 357910 579891 357922
rect 580252 357826 580356 359786
rect 580004 357814 580356 357826
rect 573878 357682 574512 357810
rect 580004 357726 580016 357814
rect 580106 357726 580356 357814
rect 580004 357722 580356 357726
rect 580004 357720 580118 357722
rect 573878 357680 574508 357682
rect 573878 357594 574408 357680
rect 573509 357576 574408 357594
rect 574500 357576 574508 357680
rect 573509 357564 574508 357576
rect 536288 357418 536408 357440
rect 560542 357510 565856 357540
rect 560542 357450 560728 357510
rect 560788 357450 560928 357510
rect 560988 357450 561128 357510
rect 561188 357450 561328 357510
rect 561388 357450 561528 357510
rect 561588 357450 561728 357510
rect 561788 357450 561928 357510
rect 561988 357450 562128 357510
rect 562188 357450 562328 357510
rect 562388 357450 562528 357510
rect 562588 357450 562728 357510
rect 562788 357450 562928 357510
rect 562988 357450 563128 357510
rect 563188 357450 563328 357510
rect 563388 357450 563528 357510
rect 563588 357450 563728 357510
rect 563788 357450 563928 357510
rect 563988 357450 564128 357510
rect 564188 357450 564328 357510
rect 564388 357450 564528 357510
rect 564588 357450 564728 357510
rect 564788 357450 564928 357510
rect 564988 357450 565128 357510
rect 565188 357450 565328 357510
rect 565388 357450 565528 357510
rect 565588 357450 565856 357510
rect 560542 357420 565856 357450
rect 574644 357440 580030 357470
rect 574644 357380 574702 357440
rect 574762 357380 574902 357440
rect 574962 357380 575102 357440
rect 575162 357380 575302 357440
rect 575362 357380 575502 357440
rect 575562 357380 575702 357440
rect 575762 357380 575902 357440
rect 575962 357380 576102 357440
rect 576162 357380 576302 357440
rect 576362 357380 576502 357440
rect 576562 357380 576702 357440
rect 576762 357380 576902 357440
rect 576962 357380 577102 357440
rect 577162 357380 577302 357440
rect 577362 357380 577502 357440
rect 577562 357380 577702 357440
rect 577762 357380 577902 357440
rect 577962 357380 578102 357440
rect 578162 357380 578302 357440
rect 578362 357380 578502 357440
rect 578562 357380 578702 357440
rect 578762 357380 578902 357440
rect 578962 357380 579102 357440
rect 579162 357380 579302 357440
rect 579362 357380 579502 357440
rect 579562 357380 579702 357440
rect 579762 357380 580030 357440
rect 574644 357350 580030 357380
rect 508352 356446 508362 356582
rect 508652 356446 508662 356582
rect 508622 356438 508658 356446
rect 566116 313610 566126 313804
rect 566346 313794 566356 313804
rect 566346 313610 566362 313794
rect 580844 313778 580948 313782
rect 580756 313770 580948 313778
rect 560404 313082 565718 313112
rect 560404 313022 560590 313082
rect 560650 313022 560790 313082
rect 560850 313022 560990 313082
rect 561050 313022 561190 313082
rect 561250 313022 561390 313082
rect 561450 313022 561590 313082
rect 561650 313022 561790 313082
rect 561850 313022 561990 313082
rect 562050 313022 562190 313082
rect 562250 313022 562390 313082
rect 562450 313022 562590 313082
rect 562650 313022 562790 313082
rect 562850 313022 562990 313082
rect 563050 313022 563190 313082
rect 563250 313022 563390 313082
rect 563450 313022 563590 313082
rect 563650 313022 563790 313082
rect 563850 313022 563990 313082
rect 564050 313022 564190 313082
rect 564250 313022 564390 313082
rect 564450 313022 564590 313082
rect 564650 313022 564790 313082
rect 564850 313022 564990 313082
rect 565050 313022 565190 313082
rect 565250 313022 565390 313082
rect 565450 313022 565718 313082
rect 560404 312992 565718 313022
rect 560409 312660 560455 312672
rect 559642 311536 559652 311744
rect 559860 311714 560240 311744
rect 559860 311564 560094 311714
rect 560226 311564 560240 311714
rect 560409 311684 560415 312660
rect 560449 311684 560455 312660
rect 560409 311672 560455 311684
rect 560667 312660 560713 312672
rect 560667 311684 560673 312660
rect 560707 311684 560713 312660
rect 560667 311672 560713 311684
rect 560925 312660 560971 312672
rect 560925 311684 560931 312660
rect 560965 311684 560971 312660
rect 560925 311672 560971 311684
rect 561183 312660 561229 312672
rect 561183 311684 561189 312660
rect 561223 311684 561229 312660
rect 561183 311672 561229 311684
rect 561441 312660 561487 312672
rect 561441 311684 561447 312660
rect 561481 311684 561487 312660
rect 561441 311672 561487 311684
rect 561699 312660 561745 312672
rect 561699 311684 561705 312660
rect 561739 311684 561745 312660
rect 561699 311672 561745 311684
rect 561957 312660 562003 312672
rect 561957 311684 561963 312660
rect 561997 311684 562003 312660
rect 561957 311672 562003 311684
rect 562215 312660 562261 312672
rect 562215 311684 562221 312660
rect 562255 311684 562261 312660
rect 562215 311672 562261 311684
rect 562473 312660 562519 312672
rect 562473 311684 562479 312660
rect 562513 311684 562519 312660
rect 562473 311672 562519 311684
rect 562731 312660 562777 312672
rect 562731 311684 562737 312660
rect 562771 311684 562777 312660
rect 562731 311672 562777 311684
rect 562989 312660 563035 312672
rect 562989 311684 562995 312660
rect 563029 311684 563035 312660
rect 562989 311672 563035 311684
rect 563247 312660 563293 312672
rect 563247 311684 563253 312660
rect 563287 311684 563293 312660
rect 563247 311672 563293 311684
rect 563505 312660 563551 312672
rect 563505 311684 563511 312660
rect 563545 311684 563551 312660
rect 563505 311672 563551 311684
rect 563763 312660 563809 312672
rect 563763 311684 563769 312660
rect 563803 311684 563809 312660
rect 563763 311672 563809 311684
rect 564021 312660 564067 312672
rect 564021 311684 564027 312660
rect 564061 311684 564067 312660
rect 564021 311672 564067 311684
rect 564279 312660 564325 312672
rect 564279 311684 564285 312660
rect 564319 311684 564325 312660
rect 564279 311672 564325 311684
rect 564537 312660 564583 312672
rect 564537 311684 564543 312660
rect 564577 311684 564583 312660
rect 564537 311672 564583 311684
rect 564795 312660 564841 312672
rect 564795 311684 564801 312660
rect 564835 311684 564841 312660
rect 564795 311672 564841 311684
rect 565053 312660 565099 312672
rect 565053 311684 565059 312660
rect 565093 311684 565099 312660
rect 565053 311672 565099 311684
rect 565311 312660 565357 312672
rect 565311 311684 565317 312660
rect 565351 311684 565357 312660
rect 565311 311672 565357 311684
rect 565569 312660 565615 312672
rect 565569 311684 565575 312660
rect 565609 311684 565615 312660
rect 566116 311684 566362 313610
rect 580748 313602 580758 313770
rect 580944 313602 580954 313770
rect 575092 313152 580478 313182
rect 575092 313092 575150 313152
rect 575210 313092 575350 313152
rect 575410 313092 575550 313152
rect 575610 313092 575750 313152
rect 575810 313092 575950 313152
rect 576010 313092 576150 313152
rect 576210 313092 576350 313152
rect 576410 313092 576550 313152
rect 576610 313092 576750 313152
rect 576810 313092 576950 313152
rect 577010 313092 577150 313152
rect 577210 313092 577350 313152
rect 577410 313092 577550 313152
rect 577610 313092 577750 313152
rect 577810 313092 577950 313152
rect 578010 313092 578150 313152
rect 578210 313092 578350 313152
rect 578410 313092 578550 313152
rect 578610 313092 578750 313152
rect 578810 313092 578950 313152
rect 579010 313092 579150 313152
rect 579210 313092 579350 313152
rect 579410 313092 579550 313152
rect 579610 313092 579750 313152
rect 579810 313092 579950 313152
rect 580010 313092 580150 313152
rect 580210 313092 580478 313152
rect 575092 313062 580478 313092
rect 575133 312730 575179 312742
rect 575133 311754 575139 312730
rect 575173 311754 575179 312730
rect 575133 311742 575179 311754
rect 575391 312730 575437 312742
rect 575391 311754 575397 312730
rect 575431 311754 575437 312730
rect 575391 311742 575437 311754
rect 575649 312730 575695 312742
rect 575649 311754 575655 312730
rect 575689 311754 575695 312730
rect 575649 311742 575695 311754
rect 575907 312730 575953 312742
rect 575907 311754 575913 312730
rect 575947 311754 575953 312730
rect 575907 311742 575953 311754
rect 576165 312730 576211 312742
rect 576165 311754 576171 312730
rect 576205 311754 576211 312730
rect 576165 311742 576211 311754
rect 576423 312730 576469 312742
rect 576423 311754 576429 312730
rect 576463 311754 576469 312730
rect 576423 311742 576469 311754
rect 576681 312730 576727 312742
rect 576681 311754 576687 312730
rect 576721 311754 576727 312730
rect 576681 311742 576727 311754
rect 576939 312730 576985 312742
rect 576939 311754 576945 312730
rect 576979 311754 576985 312730
rect 576939 311742 576985 311754
rect 577197 312730 577243 312742
rect 577197 311754 577203 312730
rect 577237 311754 577243 312730
rect 577197 311742 577243 311754
rect 577455 312730 577501 312742
rect 577455 311754 577461 312730
rect 577495 311754 577501 312730
rect 577455 311742 577501 311754
rect 577713 312730 577759 312742
rect 577713 311754 577719 312730
rect 577753 311754 577759 312730
rect 577713 311742 577759 311754
rect 577971 312730 578017 312742
rect 577971 311754 577977 312730
rect 578011 311754 578017 312730
rect 577971 311742 578017 311754
rect 578229 312730 578275 312742
rect 578229 311754 578235 312730
rect 578269 311754 578275 312730
rect 578229 311742 578275 311754
rect 578487 312730 578533 312742
rect 578487 311754 578493 312730
rect 578527 311754 578533 312730
rect 578487 311742 578533 311754
rect 578745 312730 578791 312742
rect 578745 311754 578751 312730
rect 578785 311754 578791 312730
rect 578745 311742 578791 311754
rect 579003 312730 579049 312742
rect 579003 311754 579009 312730
rect 579043 311754 579049 312730
rect 579003 311742 579049 311754
rect 579261 312730 579307 312742
rect 579261 311754 579267 312730
rect 579301 311754 579307 312730
rect 579261 311742 579307 311754
rect 579519 312730 579565 312742
rect 579519 311754 579525 312730
rect 579559 311754 579565 312730
rect 579519 311742 579565 311754
rect 579777 312730 579823 312742
rect 579777 311754 579783 312730
rect 579817 311754 579823 312730
rect 579777 311742 579823 311754
rect 580035 312730 580081 312742
rect 580035 311754 580041 312730
rect 580075 311754 580081 312730
rect 580035 311742 580081 311754
rect 580293 312730 580339 312742
rect 580293 311754 580299 312730
rect 580333 311754 580339 312730
rect 580293 311742 580339 311754
rect 565569 311672 565615 311684
rect 559860 311536 560240 311564
rect 565812 311660 566362 311684
rect 565812 311552 565828 311660
rect 565988 311552 566362 311660
rect 565812 311536 566362 311552
rect 573432 311700 574046 311742
rect 573432 311420 573492 311700
rect 573834 311590 574046 311700
rect 580756 311658 580948 313602
rect 580452 311646 580948 311658
rect 573834 311524 574952 311590
rect 580452 311558 580464 311646
rect 580554 311558 580948 311646
rect 580452 311554 580948 311558
rect 580452 311552 580566 311554
rect 573834 311512 574956 311524
rect 573834 311420 574856 311512
rect 573432 311408 574856 311420
rect 574948 311408 574956 311512
rect 573432 311396 574956 311408
rect 573432 311392 574952 311396
rect 573432 311382 574050 311392
rect 575092 311272 580478 311302
rect 560404 311202 565718 311232
rect 560404 311142 560590 311202
rect 560650 311142 560790 311202
rect 560850 311142 560990 311202
rect 561050 311142 561190 311202
rect 561250 311142 561390 311202
rect 561450 311142 561590 311202
rect 561650 311142 561790 311202
rect 561850 311142 561990 311202
rect 562050 311142 562190 311202
rect 562250 311142 562390 311202
rect 562450 311142 562590 311202
rect 562650 311142 562790 311202
rect 562850 311142 562990 311202
rect 563050 311142 563190 311202
rect 563250 311142 563390 311202
rect 563450 311142 563590 311202
rect 563650 311142 563790 311202
rect 563850 311142 563990 311202
rect 564050 311142 564190 311202
rect 564250 311142 564390 311202
rect 564450 311142 564590 311202
rect 564650 311142 564790 311202
rect 564850 311142 564990 311202
rect 565050 311142 565190 311202
rect 565250 311142 565390 311202
rect 565450 311142 565718 311202
rect 575092 311212 575150 311272
rect 575210 311212 575350 311272
rect 575410 311212 575550 311272
rect 575610 311212 575750 311272
rect 575810 311212 575950 311272
rect 576010 311212 576150 311272
rect 576210 311212 576350 311272
rect 576410 311212 576550 311272
rect 576610 311212 576750 311272
rect 576810 311212 576950 311272
rect 577010 311212 577150 311272
rect 577210 311212 577350 311272
rect 577410 311212 577550 311272
rect 577610 311212 577750 311272
rect 577810 311212 577950 311272
rect 578010 311212 578150 311272
rect 578210 311212 578350 311272
rect 578410 311212 578550 311272
rect 578610 311212 578750 311272
rect 578810 311212 578950 311272
rect 579010 311212 579150 311272
rect 579210 311212 579350 311272
rect 579410 311212 579550 311272
rect 579610 311212 579750 311272
rect 579810 311212 579950 311272
rect 580010 311212 580150 311272
rect 580210 311212 580478 311272
rect 575092 311182 580478 311212
rect 560404 311112 565718 311142
<< via1 >>
rect 566186 494126 566408 494310
rect 580856 494136 581040 494348
rect 559802 492324 560012 492536
rect 573564 491888 573874 492160
rect 491170 412444 491286 414032
rect 494930 412444 495046 414032
rect 493050 409996 493166 411584
rect 498690 412444 498806 414032
rect 494944 397218 494996 397270
rect 494740 395470 494792 395522
rect 493992 393906 494044 393958
rect 494808 391146 494860 391198
rect 494808 385485 494860 385494
rect 494808 385451 494817 385485
rect 494817 385451 494851 385485
rect 494851 385451 494860 385485
rect 494808 385442 494860 385451
rect 494536 366582 494588 366634
rect 493050 359888 493166 361476
rect 491170 357440 491286 359028
rect 496810 409996 496926 411584
rect 502450 412444 502566 414032
rect 498752 406602 498804 406654
rect 498344 400573 498396 400582
rect 498344 400539 498353 400573
rect 498353 400539 498387 400573
rect 498387 400539 498396 400573
rect 498344 400530 498396 400539
rect 498548 400389 498600 400398
rect 498548 400355 498557 400389
rect 498557 400355 498591 400389
rect 498591 400355 498600 400389
rect 498548 400346 498600 400355
rect 498480 399929 498532 399938
rect 498480 399895 498489 399929
rect 498489 399895 498523 399929
rect 498523 399895 498532 399929
rect 498480 399886 498532 399895
rect 498344 392710 498396 392762
rect 498582 385485 498634 385494
rect 498582 385451 498591 385485
rect 498591 385451 498625 385485
rect 498625 385451 498634 385485
rect 498582 385442 498634 385451
rect 497324 371660 497344 371694
rect 497344 371660 497376 371694
rect 497324 371642 497376 371660
rect 498752 371642 498804 371694
rect 498208 370814 498260 370866
rect 496810 359888 496926 361476
rect 494930 357440 495046 359028
rect 500570 409996 500686 411584
rect 506210 412444 506326 414032
rect 504330 409996 504446 411584
rect 509970 412444 510086 414032
rect 504872 402002 504924 402054
rect 506096 400990 506137 401042
rect 506137 400990 506148 401042
rect 503920 400530 503972 400582
rect 502492 399426 502544 399478
rect 502220 392710 502272 392762
rect 502220 391146 502272 391198
rect 505144 399334 505196 399386
rect 505620 398690 505672 398742
rect 505144 398322 505177 398374
rect 505177 398322 505196 398374
rect 504532 392618 504584 392670
rect 505620 392618 505672 392670
rect 505144 392526 505196 392578
rect 503988 389122 504040 389174
rect 502220 386865 502272 386874
rect 502220 386831 502229 386865
rect 502229 386831 502263 386865
rect 502263 386831 502272 386865
rect 502220 386822 502272 386831
rect 502288 386730 502340 386782
rect 502084 386546 502136 386598
rect 502356 385485 502408 385494
rect 502356 385451 502365 385485
rect 502365 385451 502399 385485
rect 502399 385451 502408 385485
rect 502356 385442 502408 385451
rect 504872 389122 504924 389174
rect 505892 386865 505944 386874
rect 505892 386831 505901 386865
rect 505901 386831 505935 386865
rect 505935 386831 505944 386865
rect 505892 386822 505944 386831
rect 505076 385442 505128 385494
rect 504396 381486 504448 381538
rect 504056 380474 504108 380526
rect 501948 379094 502000 379146
rect 504872 380474 504924 380526
rect 504056 379094 504108 379146
rect 501812 376334 501864 376386
rect 500928 372944 500980 372982
rect 500928 372930 500944 372944
rect 500944 372930 500978 372944
rect 500978 372930 500980 372944
rect 501132 372960 501184 372982
rect 501132 372930 501138 372960
rect 501138 372930 501184 372960
rect 501812 372774 501864 372798
rect 501812 372746 501842 372774
rect 501842 372746 501864 372774
rect 501268 370814 501320 370866
rect 502492 372953 502525 372982
rect 502525 372953 502544 372982
rect 502492 372930 502544 372953
rect 502152 366582 502204 366634
rect 500570 359888 500686 361476
rect 498690 357440 498806 359028
rect 506028 377389 506080 377398
rect 506028 377355 506037 377389
rect 506037 377355 506080 377389
rect 506028 377346 506080 377355
rect 506096 376377 506148 376386
rect 506096 376343 506105 376377
rect 506105 376343 506139 376377
rect 506139 376343 506148 376377
rect 506096 376334 506148 376343
rect 504872 372960 504924 372982
rect 504872 372930 504898 372960
rect 504898 372930 504924 372960
rect 506232 372953 506251 372982
rect 506251 372953 506284 372982
rect 506232 372930 506284 372953
rect 505552 372774 505604 372798
rect 505552 372746 505568 372774
rect 505568 372746 505602 372774
rect 505602 372746 505604 372774
rect 504330 359888 504446 361476
rect 502450 357440 502566 359028
rect 508090 409996 508206 411584
rect 509360 398322 509412 398374
rect 508408 395470 508460 395522
rect 513730 412444 513846 414032
rect 508884 390410 508936 390462
rect 508136 381486 508188 381538
rect 508476 373034 508528 373074
rect 508476 373022 508498 373034
rect 508498 373022 508528 373034
rect 508272 366214 508324 366266
rect 508090 359888 508206 361476
rect 506210 357440 506326 359028
rect 508816 372774 508868 372798
rect 508816 372746 508828 372774
rect 508828 372746 508862 372774
rect 508862 372746 508868 372774
rect 509360 372674 509412 372706
rect 509360 372654 509362 372674
rect 509362 372654 509412 372674
rect 511850 409996 511966 411584
rect 512624 398230 512676 398282
rect 517490 412444 517606 414032
rect 513100 396482 513152 396534
rect 512624 395838 512676 395890
rect 512012 393998 512064 394050
rect 513100 393998 513152 394050
rect 513100 393170 513152 393222
rect 512148 392710 512159 392762
rect 512159 392710 512200 392762
rect 512012 392526 512064 392578
rect 513100 390410 513152 390462
rect 512624 387466 512676 387518
rect 511876 381486 511928 381538
rect 513644 376377 513696 376386
rect 513644 376343 513653 376377
rect 513653 376343 513687 376377
rect 513687 376343 513696 376377
rect 513644 376334 513696 376343
rect 512352 372780 512404 372798
rect 512352 372746 512384 372780
rect 512384 372746 512404 372780
rect 512556 372674 512608 372706
rect 512556 372654 512588 372674
rect 512588 372654 512608 372674
rect 513100 366490 513152 366542
rect 513780 372787 513832 372798
rect 513780 372753 513805 372787
rect 513805 372753 513832 372787
rect 513780 372746 513832 372753
rect 511850 359888 511966 361476
rect 509970 357440 510086 359028
rect 515610 409996 515726 411584
rect 516160 400990 516212 401042
rect 521250 412444 521366 414032
rect 517384 391974 517436 392026
rect 516908 389524 516960 389542
rect 516908 389490 516925 389524
rect 516925 389490 516960 389524
rect 517180 387417 517232 387426
rect 517180 387383 517189 387417
rect 517189 387383 517223 387417
rect 517223 387383 517232 387417
rect 517180 387374 517232 387383
rect 516296 385442 516348 385494
rect 515616 381486 515668 381538
rect 519370 409996 519486 411584
rect 520648 398230 520700 398282
rect 519696 391974 519748 392026
rect 525010 412444 525126 414032
rect 520648 387466 520700 387518
rect 520172 385810 520224 385862
rect 520648 385166 520700 385218
rect 518608 383970 518660 384022
rect 517384 377541 517436 377582
rect 517384 377530 517417 377541
rect 517417 377530 517436 377541
rect 519696 383970 519748 384022
rect 519560 379922 519612 379974
rect 518608 377530 518660 377582
rect 517860 376610 517912 376662
rect 515820 374954 515872 375006
rect 516908 374954 516960 375006
rect 516432 374797 516484 374822
rect 516432 374770 516457 374797
rect 516457 374770 516484 374797
rect 515888 373482 515940 373534
rect 516364 372194 516416 372246
rect 517384 372053 517436 372062
rect 517384 372010 517417 372053
rect 517417 372010 517436 372053
rect 520648 379922 520700 379974
rect 520172 379830 520224 379882
rect 520648 379186 520700 379238
rect 519696 376610 519748 376662
rect 519560 374770 519612 374822
rect 517860 372010 517912 372062
rect 515820 368882 515872 368934
rect 516908 368915 516960 368934
rect 516908 368882 516960 368915
rect 515820 366398 515872 366450
rect 516432 366306 516457 366358
rect 516457 366306 516484 366358
rect 516908 366490 516960 366542
rect 515610 359888 515726 361476
rect 513730 357440 513846 359028
rect 520648 373482 520700 373534
rect 519560 372194 519612 372246
rect 519560 366398 519612 366450
rect 520648 366306 520700 366358
rect 519370 359888 519486 361476
rect 517490 357440 517606 359028
rect 523130 409996 523246 411584
rect 528770 412444 528886 414032
rect 524864 389533 524916 389542
rect 524864 389499 524907 389533
rect 524907 389499 524916 389533
rect 524864 389490 524916 389499
rect 524796 380609 524848 380618
rect 524796 380575 524805 380609
rect 524805 380575 524839 380609
rect 524839 380575 524848 380609
rect 524796 380566 524848 380575
rect 524660 370906 524712 370958
rect 523130 359888 523246 361476
rect 521250 357440 521366 359028
rect 526890 409996 527006 411584
rect 528196 370679 528248 370682
rect 528196 370630 528248 370679
rect 532530 412444 532646 414032
rect 527040 365846 527092 365898
rect 527176 370538 527228 370590
rect 527720 368238 527737 368290
rect 527737 368238 527772 368290
rect 528672 367962 528697 368014
rect 528697 367962 528724 368014
rect 528672 365386 528697 365438
rect 528697 365386 528724 365438
rect 526890 359888 527006 361476
rect 525010 357440 525126 359028
rect 530650 409996 530766 411584
rect 530984 370906 531036 370958
rect 536290 412444 536406 414032
rect 530848 370170 530900 370222
rect 532412 369250 532464 369302
rect 534410 409996 534526 411584
rect 535676 370170 535679 370222
rect 535679 370170 535728 370222
rect 566256 405258 566462 405476
rect 580074 405292 580182 405402
rect 559736 403192 559926 403368
rect 573538 402980 573888 403312
rect 537512 389398 537564 389450
rect 537512 387374 537564 387426
rect 532684 369250 532736 369302
rect 531936 368238 531988 368290
rect 530848 367962 530900 368014
rect 531936 365846 531988 365898
rect 532684 365018 532736 365070
rect 530650 359888 530766 361476
rect 528770 357440 528886 359028
rect 534724 365754 534776 365806
rect 534588 365110 534640 365162
rect 535676 365110 535728 365162
rect 534724 365018 534776 365070
rect 534410 359888 534526 361476
rect 532530 357440 532646 359028
rect 566274 359786 566500 359978
rect 580252 359786 580358 359906
rect 536290 357440 536406 359028
rect 559712 357844 559920 358052
rect 573540 357594 573878 357920
rect 508362 356446 508652 356582
rect 566126 313610 566346 313804
rect 559652 311536 559860 311744
rect 580758 313602 580944 313770
rect 573492 311420 573834 311700
<< metal2 >>
rect 580856 494348 581040 494358
rect 566186 494310 566408 494320
rect 580856 494126 581040 494136
rect 566186 494116 566408 494126
rect 559802 492536 560012 492546
rect 559802 492314 560012 492324
rect 573564 492160 573874 492170
rect 573564 491878 573874 491888
rect 491168 414032 491288 414054
rect 491168 412444 491170 414032
rect 491286 412444 491288 414032
rect 491168 412422 491288 412444
rect 494928 414032 495048 414054
rect 494928 412444 494930 414032
rect 495046 412444 495048 414032
rect 494928 412422 495048 412444
rect 498688 414032 498808 414054
rect 498688 412444 498690 414032
rect 498806 412444 498808 414032
rect 498688 412422 498808 412444
rect 502448 414032 502568 414054
rect 502448 412444 502450 414032
rect 502566 412444 502568 414032
rect 502448 412422 502568 412444
rect 506208 414032 506328 414054
rect 506208 412444 506210 414032
rect 506326 412444 506328 414032
rect 506208 412422 506328 412444
rect 509968 414032 510088 414054
rect 509968 412444 509970 414032
rect 510086 412444 510088 414032
rect 509968 412422 510088 412444
rect 513728 414032 513848 414054
rect 513728 412444 513730 414032
rect 513846 412444 513848 414032
rect 513728 412422 513848 412444
rect 517488 414032 517608 414054
rect 517488 412444 517490 414032
rect 517606 412444 517608 414032
rect 517488 412422 517608 412444
rect 521248 414032 521368 414054
rect 521248 412444 521250 414032
rect 521366 412444 521368 414032
rect 521248 412422 521368 412444
rect 525008 414032 525128 414054
rect 525008 412444 525010 414032
rect 525126 412444 525128 414032
rect 525008 412422 525128 412444
rect 528768 414032 528888 414054
rect 528768 412444 528770 414032
rect 528886 412444 528888 414032
rect 528768 412422 528888 412444
rect 532528 414032 532648 414054
rect 532528 412444 532530 414032
rect 532646 412444 532648 414032
rect 532528 412422 532648 412444
rect 536288 414032 536408 414054
rect 536288 412444 536290 414032
rect 536406 412444 536408 414032
rect 536288 412422 536408 412444
rect 493048 411584 493168 411606
rect 493048 409996 493050 411584
rect 493166 409996 493168 411584
rect 493048 409974 493168 409996
rect 496808 411584 496928 411606
rect 496808 409996 496810 411584
rect 496926 409996 496928 411584
rect 496808 409974 496928 409996
rect 500568 411584 500688 411606
rect 500568 409996 500570 411584
rect 500686 409996 500688 411584
rect 500568 409974 500688 409996
rect 504328 411584 504448 411606
rect 504328 409996 504330 411584
rect 504446 409996 504448 411584
rect 504328 409974 504448 409996
rect 508088 411584 508208 411606
rect 508088 409996 508090 411584
rect 508206 409996 508208 411584
rect 508088 409974 508208 409996
rect 511848 411584 511968 411606
rect 511848 409996 511850 411584
rect 511966 409996 511968 411584
rect 511848 409974 511968 409996
rect 515608 411584 515728 411606
rect 515608 409996 515610 411584
rect 515726 409996 515728 411584
rect 515608 409974 515728 409996
rect 519368 411584 519488 411606
rect 519368 409996 519370 411584
rect 519486 409996 519488 411584
rect 519368 409974 519488 409996
rect 523128 411584 523248 411606
rect 523128 409996 523130 411584
rect 523246 409996 523248 411584
rect 523128 409974 523248 409996
rect 526888 411584 527008 411606
rect 526888 409996 526890 411584
rect 527006 409996 527008 411584
rect 526888 409974 527008 409996
rect 530648 411584 530768 411606
rect 530648 409996 530650 411584
rect 530766 409996 530768 411584
rect 530648 409974 530768 409996
rect 534408 411584 534528 411606
rect 534408 409996 534410 411584
rect 534526 409996 534528 411584
rect 534408 409974 534528 409996
rect 493338 409006 493418 409038
rect 493338 408950 493350 409006
rect 493406 408950 493418 409006
rect 493338 408926 493418 408950
rect 493338 408870 493350 408926
rect 493406 408870 493418 408926
rect 493338 408838 493418 408870
rect 494748 408964 494848 409016
rect 494748 408908 494770 408964
rect 494826 408908 494848 408964
rect 494748 408856 494848 408908
rect 497098 409006 497178 409038
rect 497098 408950 497110 409006
rect 497166 408950 497178 409006
rect 497098 408926 497178 408950
rect 497098 408870 497110 408926
rect 497166 408870 497178 408926
rect 497098 408838 497178 408870
rect 498508 408964 498608 409016
rect 498508 408908 498530 408964
rect 498586 408908 498608 408964
rect 498508 408856 498608 408908
rect 500858 408614 500938 408646
rect 500858 408558 500870 408614
rect 500926 408558 500938 408614
rect 500858 408534 500938 408558
rect 500858 408478 500870 408534
rect 500926 408478 500938 408534
rect 500858 408446 500938 408478
rect 502268 408572 502368 408624
rect 502268 408516 502290 408572
rect 502346 408516 502368 408572
rect 502268 408464 502368 408516
rect 498701 406600 498710 406656
rect 498766 406654 498775 406656
rect 498804 406602 498810 406654
rect 498766 406600 498775 406602
rect 566256 405476 566462 405486
rect 580074 405402 580182 405412
rect 580074 405282 580182 405292
rect 566256 405248 566462 405258
rect 559736 403368 559926 403378
rect 559736 403182 559926 403192
rect 573538 403312 573888 403322
rect 573538 402970 573888 402980
rect 504801 402000 504810 402056
rect 504866 402054 504875 402056
rect 504866 402002 504872 402054
rect 504924 402002 504930 402054
rect 504866 402000 504875 402002
rect 493338 401558 493418 401590
rect 493338 401502 493350 401558
rect 493406 401502 493418 401558
rect 493338 401478 493418 401502
rect 493338 401422 493350 401478
rect 493406 401422 493418 401478
rect 493338 401390 493418 401422
rect 494748 401516 494848 401568
rect 494748 401460 494770 401516
rect 494826 401460 494848 401516
rect 494748 401408 494848 401460
rect 506090 400990 506096 401042
rect 506148 401030 506154 401042
rect 516154 401030 516160 401042
rect 506148 401002 516160 401030
rect 506148 400990 506154 401002
rect 516154 400990 516160 401002
rect 516212 400990 516218 401042
rect 498338 400530 498344 400582
rect 498396 400570 498402 400582
rect 503914 400570 503920 400582
rect 498396 400542 503920 400570
rect 498396 400530 498402 400542
rect 503914 400530 503920 400542
rect 503972 400530 503978 400582
rect 498579 400398 498588 400400
rect 498542 400346 498548 400398
rect 498579 400344 498588 400346
rect 498644 400344 498653 400400
rect 498213 399884 498222 399940
rect 498278 399926 498287 399940
rect 498474 399926 498480 399938
rect 498278 399898 498480 399926
rect 498278 399884 498287 399898
rect 498474 399886 498480 399898
rect 498532 399886 498538 399938
rect 500858 399794 500938 399826
rect 500858 399738 500870 399794
rect 500926 399738 500938 399794
rect 500858 399714 500938 399738
rect 500858 399658 500870 399714
rect 500926 399658 500938 399714
rect 500858 399626 500938 399658
rect 502268 399752 502368 399804
rect 502268 399696 502290 399752
rect 502346 399696 502368 399752
rect 502268 399644 502368 399696
rect 502361 399424 502370 399480
rect 502426 399466 502435 399480
rect 502486 399466 502492 399478
rect 502426 399438 502492 399466
rect 502426 399424 502435 399438
rect 502486 399426 502492 399438
rect 502544 399426 502550 399478
rect 505138 399334 505144 399386
rect 505196 399334 505202 399386
rect 505156 398730 505184 399334
rect 505614 398730 505620 398742
rect 505156 398702 505620 398730
rect 505614 398690 505620 398702
rect 505672 398690 505678 398742
rect 505138 398322 505144 398374
rect 505196 398362 505202 398374
rect 509354 398362 509360 398374
rect 505196 398334 509360 398362
rect 505196 398322 505202 398334
rect 509354 398322 509360 398334
rect 509412 398322 509418 398374
rect 512618 398230 512624 398282
rect 512676 398270 512682 398282
rect 520642 398270 520648 398282
rect 512676 398242 520648 398270
rect 512676 398230 512682 398242
rect 520642 398230 520648 398242
rect 520700 398230 520706 398282
rect 494919 397216 494928 397272
rect 494984 397270 494993 397272
rect 494996 397258 495002 397270
rect 494996 397230 495016 397258
rect 494996 397218 495002 397230
rect 494984 397216 494993 397218
rect 513094 396522 513100 396534
rect 512636 396494 513100 396522
rect 512636 395890 512664 396494
rect 513094 396482 513100 396494
rect 513152 396482 513158 396534
rect 512618 395838 512624 395890
rect 512676 395838 512682 395890
rect 494734 395470 494740 395522
rect 494792 395510 494798 395522
rect 508402 395510 508408 395522
rect 494792 395482 508408 395510
rect 494792 395470 494798 395482
rect 508402 395470 508408 395482
rect 508460 395470 508466 395522
rect 512006 393998 512012 394050
rect 512064 394038 512070 394050
rect 513094 394038 513100 394050
rect 512064 394010 513100 394038
rect 512064 393998 512070 394010
rect 513094 393998 513100 394010
rect 513152 393998 513158 394050
rect 493986 393906 493992 393958
rect 494044 393946 494050 393958
rect 494044 393918 512936 393946
rect 494044 393906 494050 393918
rect 512908 393210 512936 393918
rect 513094 393210 513100 393222
rect 512908 393182 513100 393210
rect 513094 393170 513100 393182
rect 513152 393170 513158 393222
rect 498338 392710 498344 392762
rect 498396 392750 498402 392762
rect 500653 392750 500662 392764
rect 498396 392722 500662 392750
rect 498396 392710 498402 392722
rect 500653 392708 500662 392722
rect 500718 392750 500727 392764
rect 502214 392750 502220 392762
rect 500718 392722 502220 392750
rect 500718 392708 500727 392722
rect 502214 392710 502220 392722
rect 502272 392750 502278 392762
rect 512142 392750 512148 392762
rect 502272 392722 512148 392750
rect 502272 392710 502278 392722
rect 512142 392710 512148 392722
rect 512200 392710 512206 392762
rect 504526 392618 504532 392670
rect 504584 392658 504590 392670
rect 505614 392658 505620 392670
rect 504584 392630 505620 392658
rect 504584 392618 504590 392630
rect 505614 392618 505620 392630
rect 505672 392618 505678 392670
rect 505138 392526 505144 392578
rect 505196 392566 505202 392578
rect 512006 392566 512012 392578
rect 505196 392538 512012 392566
rect 505196 392526 505202 392538
rect 512006 392526 512012 392538
rect 512064 392526 512070 392578
rect 517378 391974 517384 392026
rect 517436 392014 517442 392026
rect 519690 392014 519696 392026
rect 517436 391986 519696 392014
rect 517436 391974 517442 391986
rect 519690 391974 519696 391986
rect 519748 391974 519754 392026
rect 494802 391146 494808 391198
rect 494860 391186 494866 391198
rect 498579 391186 498588 391200
rect 494860 391158 498588 391186
rect 494860 391146 494866 391158
rect 498579 391144 498588 391158
rect 498644 391186 498653 391200
rect 502214 391186 502220 391198
rect 498644 391158 502220 391186
rect 498644 391144 498653 391158
rect 502214 391146 502220 391158
rect 502272 391146 502278 391198
rect 508878 390410 508884 390462
rect 508936 390450 508942 390462
rect 513094 390450 513100 390462
rect 508936 390422 513100 390450
rect 508936 390410 508942 390422
rect 513094 390410 513100 390422
rect 513152 390410 513158 390462
rect 516902 389490 516908 389542
rect 516960 389530 516966 389542
rect 524858 389530 524864 389542
rect 516960 389502 524864 389530
rect 516960 389490 516966 389502
rect 524858 389490 524864 389502
rect 524916 389490 524922 389542
rect 541952 389470 542058 389480
rect 537506 389398 537512 389450
rect 537564 389438 537570 389450
rect 537564 389410 541952 389438
rect 537564 389398 537570 389410
rect 542058 389410 542060 389438
rect 541952 389378 542058 389388
rect 503982 389122 503988 389174
rect 504040 389162 504046 389174
rect 504866 389162 504872 389174
rect 504040 389134 504872 389162
rect 504040 389122 504046 389134
rect 504866 389122 504872 389134
rect 504924 389122 504930 389174
rect 508378 388720 508458 388752
rect 508378 388664 508390 388720
rect 508446 388664 508458 388720
rect 508378 388640 508458 388664
rect 508378 388584 508390 388640
rect 508446 388584 508458 388640
rect 508378 388552 508458 388584
rect 509788 388678 509888 388730
rect 509788 388622 509810 388678
rect 509866 388622 509888 388678
rect 509788 388570 509888 388622
rect 512618 387466 512624 387518
rect 512676 387506 512682 387518
rect 520642 387506 520648 387518
rect 512676 387478 520648 387506
rect 512676 387466 512682 387478
rect 520642 387466 520648 387478
rect 520700 387466 520706 387518
rect 517174 387374 517180 387426
rect 517232 387414 517238 387426
rect 537506 387414 537512 387426
rect 517232 387386 537512 387414
rect 517232 387374 517238 387386
rect 537506 387374 537512 387386
rect 537564 387374 537570 387426
rect 502214 386822 502220 386874
rect 502272 386862 502278 386874
rect 505886 386862 505892 386874
rect 502272 386834 505892 386862
rect 502272 386822 502278 386834
rect 505886 386822 505892 386834
rect 505944 386822 505950 386874
rect 502282 386730 502288 386782
rect 502340 386730 502346 386782
rect 502078 386546 502084 386598
rect 502136 386586 502142 386598
rect 502300 386586 502328 386730
rect 502136 386558 502328 386586
rect 502136 386546 502142 386558
rect 520166 385810 520172 385862
rect 520224 385850 520230 385862
rect 520224 385822 520688 385850
rect 520224 385810 520230 385822
rect 494802 385442 494808 385494
rect 494860 385482 494866 385494
rect 498576 385482 498582 385494
rect 494860 385454 498582 385482
rect 494860 385442 494866 385454
rect 498576 385442 498582 385454
rect 498634 385482 498640 385494
rect 502350 385482 502356 385494
rect 498634 385454 502356 385482
rect 498634 385442 498640 385454
rect 502350 385442 502356 385454
rect 502408 385482 502414 385494
rect 505045 385482 505054 385496
rect 505110 385494 505119 385496
rect 502408 385454 505054 385482
rect 502408 385442 502414 385454
rect 505045 385440 505054 385454
rect 505128 385482 505134 385494
rect 505128 385454 505142 385482
rect 505128 385442 505134 385454
rect 505110 385440 505119 385442
rect 516269 385440 516278 385496
rect 516334 385494 516343 385496
rect 516348 385482 516354 385494
rect 516348 385454 516366 385482
rect 516348 385442 516354 385454
rect 516334 385440 516343 385442
rect 520660 385218 520688 385822
rect 520642 385166 520648 385218
rect 520700 385166 520706 385218
rect 504618 384996 504698 385028
rect 504618 384940 504630 384996
rect 504686 384940 504698 384996
rect 504618 384916 504698 384940
rect 504618 384860 504630 384916
rect 504686 384860 504698 384916
rect 504618 384828 504698 384860
rect 506028 384954 506128 385006
rect 506028 384898 506050 384954
rect 506106 384898 506128 384954
rect 506028 384846 506128 384898
rect 512138 384996 512218 385028
rect 512138 384940 512150 384996
rect 512206 384940 512218 384996
rect 512138 384916 512218 384940
rect 512138 384860 512150 384916
rect 512206 384860 512218 384916
rect 512138 384828 512218 384860
rect 513548 384954 513648 385006
rect 513548 384898 513570 384954
rect 513626 384898 513648 384954
rect 513548 384846 513648 384898
rect 515898 384996 515978 385028
rect 515898 384940 515910 384996
rect 515966 384940 515978 384996
rect 515898 384916 515978 384940
rect 515898 384860 515910 384916
rect 515966 384860 515978 384916
rect 515898 384828 515978 384860
rect 517308 384954 517408 385006
rect 517308 384898 517330 384954
rect 517386 384898 517408 384954
rect 517308 384846 517408 384898
rect 518602 383970 518608 384022
rect 518660 384010 518666 384022
rect 519690 384010 519696 384022
rect 518660 383982 519696 384010
rect 518660 383970 518666 383982
rect 519690 383970 519696 383982
rect 519748 383970 519754 384022
rect 504435 381538 504444 381540
rect 504390 381486 504396 381538
rect 504435 381484 504444 381486
rect 504500 381484 504509 381540
rect 508130 381538 508226 381540
rect 508130 381486 508136 381538
rect 508188 381486 508226 381538
rect 508130 381484 508226 381486
rect 508282 381484 508291 381540
rect 511877 381538 511886 381540
rect 511870 381486 511876 381538
rect 511942 381526 511951 381540
rect 515659 381538 515668 381540
rect 511942 381498 511967 381526
rect 511877 381484 511886 381486
rect 511942 381484 511951 381498
rect 515610 381486 515616 381538
rect 515659 381484 515668 381486
rect 515724 381484 515733 381540
rect 508378 381272 508458 381304
rect 508378 381216 508390 381272
rect 508446 381216 508458 381272
rect 508378 381192 508458 381216
rect 508378 381136 508390 381192
rect 508446 381136 508458 381192
rect 508378 381104 508458 381136
rect 509788 381230 509888 381282
rect 509788 381174 509810 381230
rect 509866 381174 509888 381230
rect 509788 381122 509888 381174
rect 541958 380644 542066 380654
rect 524790 380566 524796 380618
rect 524848 380606 524854 380618
rect 524848 380578 541958 380606
rect 524848 380566 524854 380578
rect 542066 380564 542068 380620
rect 541958 380562 542068 380564
rect 541958 380554 542066 380562
rect 504050 380474 504056 380526
rect 504108 380514 504114 380526
rect 504866 380514 504872 380526
rect 504108 380486 504872 380514
rect 504108 380474 504114 380486
rect 504866 380474 504872 380486
rect 504924 380474 504930 380526
rect 519554 379922 519560 379974
rect 519612 379962 519618 379974
rect 520642 379962 520648 379974
rect 519612 379934 520648 379962
rect 519612 379922 519618 379934
rect 520642 379922 520648 379934
rect 520700 379922 520706 379974
rect 520166 379830 520172 379882
rect 520224 379870 520230 379882
rect 520224 379842 520688 379870
rect 520224 379830 520230 379842
rect 520660 379238 520688 379842
rect 520642 379186 520648 379238
rect 520700 379186 520706 379238
rect 501942 379094 501948 379146
rect 502000 379134 502006 379146
rect 504050 379134 504056 379146
rect 502000 379106 504056 379134
rect 502000 379094 502006 379106
rect 504050 379094 504056 379106
rect 504108 379094 504114 379146
rect 517378 377530 517384 377582
rect 517436 377570 517442 377582
rect 518602 377570 518608 377582
rect 517436 377542 518608 377570
rect 517436 377530 517442 377542
rect 518602 377530 518608 377542
rect 518660 377530 518666 377582
rect 506021 377398 506030 377400
rect 506021 377346 506028 377398
rect 506086 377386 506095 377400
rect 506086 377358 506118 377386
rect 506021 377344 506030 377346
rect 506086 377344 506095 377358
rect 517854 376610 517860 376662
rect 517912 376650 517918 376662
rect 519690 376650 519696 376662
rect 517912 376622 519696 376650
rect 517912 376610 517918 376622
rect 519690 376610 519696 376622
rect 519748 376610 519754 376662
rect 501806 376334 501812 376386
rect 501864 376374 501870 376386
rect 506090 376374 506096 376386
rect 501864 376346 506096 376374
rect 501864 376334 501870 376346
rect 506090 376334 506096 376346
rect 506148 376374 506154 376386
rect 513638 376374 513644 376386
rect 506148 376346 513644 376374
rect 506148 376334 506154 376346
rect 513638 376334 513644 376346
rect 513696 376334 513702 376386
rect 515814 374954 515820 375006
rect 515872 374994 515878 375006
rect 516902 374994 516908 375006
rect 515872 374966 516908 374994
rect 515872 374954 515878 374966
rect 516902 374954 516908 374966
rect 516960 374954 516966 375006
rect 516426 374770 516432 374822
rect 516484 374810 516490 374822
rect 519554 374810 519560 374822
rect 516484 374782 519560 374810
rect 516484 374770 516490 374782
rect 519554 374770 519560 374782
rect 519612 374770 519618 374822
rect 515882 373482 515888 373534
rect 515940 373522 515946 373534
rect 520642 373522 520648 373534
rect 515940 373494 520648 373522
rect 515940 373482 515946 373494
rect 520642 373482 520648 373494
rect 520700 373482 520706 373534
rect 508470 373062 508476 373074
rect 508284 373034 508476 373062
rect 500922 372930 500928 372982
rect 500980 372970 500986 372982
rect 501126 372970 501132 372982
rect 500980 372942 501132 372970
rect 500980 372930 500986 372942
rect 501126 372930 501132 372942
rect 501184 372970 501190 372982
rect 502486 372970 502492 372982
rect 501184 372942 502492 372970
rect 501184 372930 501190 372942
rect 502486 372930 502492 372942
rect 502544 372930 502550 372982
rect 504866 372930 504872 372982
rect 504924 372970 504930 372982
rect 506226 372970 506232 372982
rect 504924 372942 506232 372970
rect 504924 372930 504930 372942
rect 506226 372930 506232 372942
rect 506284 372970 506290 372982
rect 508284 372970 508312 373034
rect 508470 373022 508476 373034
rect 508528 373022 508534 373074
rect 506284 372942 508312 372970
rect 506284 372930 506290 372942
rect 501806 372746 501812 372798
rect 501864 372786 501870 372798
rect 505546 372786 505552 372798
rect 501864 372758 505552 372786
rect 501864 372746 501870 372758
rect 505546 372746 505552 372758
rect 505604 372786 505610 372798
rect 508810 372786 508816 372798
rect 505604 372758 508816 372786
rect 505604 372746 505610 372758
rect 508810 372746 508816 372758
rect 508868 372746 508874 372798
rect 512346 372746 512352 372798
rect 512404 372786 512410 372798
rect 513774 372786 513780 372798
rect 512404 372758 513780 372786
rect 512404 372746 512410 372758
rect 513774 372746 513780 372758
rect 513832 372746 513838 372798
rect 509354 372654 509360 372706
rect 509412 372694 509418 372706
rect 512550 372694 512556 372706
rect 509412 372666 512556 372694
rect 509412 372654 509418 372666
rect 512550 372654 512556 372666
rect 512608 372654 512614 372706
rect 516358 372194 516364 372246
rect 516416 372234 516422 372246
rect 519554 372234 519560 372246
rect 516416 372206 519560 372234
rect 516416 372194 516422 372206
rect 519554 372194 519560 372206
rect 519612 372194 519618 372246
rect 517378 372010 517384 372062
rect 517436 372050 517442 372062
rect 517854 372050 517860 372062
rect 517436 372022 517860 372050
rect 517436 372010 517442 372022
rect 517854 372010 517860 372022
rect 517912 372010 517918 372062
rect 497318 371642 497324 371694
rect 497376 371682 497382 371694
rect 498746 371682 498752 371694
rect 497376 371654 498752 371682
rect 497376 371642 497382 371654
rect 498746 371642 498752 371654
rect 498804 371642 498810 371694
rect 524654 370906 524660 370958
rect 524712 370946 524718 370958
rect 530978 370946 530984 370958
rect 524712 370918 530984 370946
rect 524712 370906 524718 370918
rect 530978 370906 530984 370918
rect 531036 370906 531042 370958
rect 498202 370814 498208 370866
rect 498260 370854 498266 370866
rect 501262 370854 501268 370866
rect 498260 370826 501268 370854
rect 498260 370814 498266 370826
rect 501262 370814 501268 370826
rect 501320 370814 501326 370866
rect 528190 370670 528196 370682
rect 527188 370642 528196 370670
rect 527188 370590 527216 370642
rect 528190 370630 528196 370642
rect 528248 370630 528254 370682
rect 527170 370538 527176 370590
rect 527228 370538 527234 370590
rect 530842 370170 530848 370222
rect 530900 370210 530906 370222
rect 535670 370210 535676 370222
rect 530900 370182 535676 370210
rect 530900 370170 530906 370182
rect 535670 370170 535676 370182
rect 535728 370170 535734 370222
rect 532406 369250 532412 369302
rect 532464 369290 532470 369302
rect 532678 369290 532684 369302
rect 532464 369262 532684 369290
rect 532464 369250 532470 369262
rect 532678 369250 532684 369262
rect 532736 369250 532742 369302
rect 515814 368882 515820 368934
rect 515872 368922 515878 368934
rect 516902 368922 516908 368934
rect 515872 368894 516908 368922
rect 515872 368882 515878 368894
rect 516902 368882 516908 368894
rect 516960 368882 516966 368934
rect 527714 368238 527720 368290
rect 527772 368278 527778 368290
rect 531930 368278 531936 368290
rect 527772 368250 531936 368278
rect 527772 368238 527778 368250
rect 531930 368238 531936 368250
rect 531988 368238 531994 368290
rect 528666 367962 528672 368014
rect 528724 368002 528730 368014
rect 530842 368002 530848 368014
rect 528724 367974 530848 368002
rect 528724 367962 528730 367974
rect 530842 367962 530848 367974
rect 530900 367962 530906 368014
rect 494530 366582 494536 366634
rect 494588 366622 494594 366634
rect 502146 366622 502152 366634
rect 494588 366594 502152 366622
rect 494588 366582 494594 366594
rect 502146 366582 502152 366594
rect 502204 366622 502210 366634
rect 502204 366594 504912 366622
rect 502204 366582 502210 366594
rect 504884 366438 504912 366594
rect 513094 366490 513100 366542
rect 513152 366530 513158 366542
rect 516902 366530 516908 366542
rect 513152 366502 516908 366530
rect 513152 366490 513158 366502
rect 516902 366490 516908 366502
rect 516960 366490 516966 366542
rect 515814 366438 515820 366450
rect 504884 366410 515820 366438
rect 508284 366266 508312 366410
rect 515814 366398 515820 366410
rect 515872 366438 515878 366450
rect 519554 366438 519560 366450
rect 515872 366410 519560 366438
rect 515872 366398 515878 366410
rect 519554 366398 519560 366410
rect 519612 366398 519618 366450
rect 516426 366306 516432 366358
rect 516484 366346 516490 366358
rect 520642 366346 520648 366358
rect 516484 366318 520648 366346
rect 516484 366306 516490 366318
rect 520642 366306 520648 366318
rect 520700 366306 520706 366358
rect 508266 366214 508272 366266
rect 508324 366214 508330 366266
rect 527034 365846 527040 365898
rect 527092 365886 527098 365898
rect 531930 365886 531936 365898
rect 527092 365858 531936 365886
rect 527092 365846 527098 365858
rect 531930 365846 531936 365858
rect 531988 365846 531994 365898
rect 534718 365794 534724 365806
rect 534532 365766 534724 365794
rect 528666 365386 528672 365438
rect 528724 365426 528730 365438
rect 534532 365426 534560 365766
rect 534718 365754 534724 365766
rect 534776 365754 534782 365806
rect 528724 365398 534560 365426
rect 528724 365386 528730 365398
rect 534582 365110 534588 365162
rect 534640 365150 534646 365162
rect 535670 365150 535676 365162
rect 534640 365122 535676 365150
rect 534640 365110 534646 365122
rect 535670 365110 535676 365122
rect 535728 365110 535734 365162
rect 532678 365018 532684 365070
rect 532736 365058 532742 365070
rect 534718 365058 534724 365070
rect 532736 365030 534724 365058
rect 532736 365018 532742 365030
rect 534718 365018 534724 365030
rect 534776 365018 534782 365070
rect 493048 361476 493168 361498
rect 493048 359888 493050 361476
rect 493166 359888 493168 361476
rect 493048 359866 493168 359888
rect 496808 361476 496928 361498
rect 496808 359888 496810 361476
rect 496926 359888 496928 361476
rect 496808 359866 496928 359888
rect 500568 361476 500688 361498
rect 500568 359888 500570 361476
rect 500686 359888 500688 361476
rect 500568 359866 500688 359888
rect 504328 361476 504448 361498
rect 504328 359888 504330 361476
rect 504446 359888 504448 361476
rect 504328 359866 504448 359888
rect 508088 361476 508208 361498
rect 508088 359888 508090 361476
rect 508206 359888 508208 361476
rect 508088 359866 508208 359888
rect 511848 361476 511968 361498
rect 511848 359888 511850 361476
rect 511966 359888 511968 361476
rect 511848 359866 511968 359888
rect 515608 361476 515728 361498
rect 515608 359888 515610 361476
rect 515726 359888 515728 361476
rect 515608 359866 515728 359888
rect 519368 361476 519488 361498
rect 519368 359888 519370 361476
rect 519486 359888 519488 361476
rect 519368 359866 519488 359888
rect 523128 361476 523248 361498
rect 523128 359888 523130 361476
rect 523246 359888 523248 361476
rect 523128 359866 523248 359888
rect 526888 361476 527008 361498
rect 526888 359888 526890 361476
rect 527006 359888 527008 361476
rect 526888 359866 527008 359888
rect 530648 361476 530768 361498
rect 530648 359888 530650 361476
rect 530766 359888 530768 361476
rect 530648 359866 530768 359888
rect 534408 361476 534528 361498
rect 534408 359888 534410 361476
rect 534526 359888 534528 361476
rect 534408 359866 534528 359888
rect 566274 359978 566500 359988
rect 566274 359776 566500 359786
rect 580252 359906 580358 359916
rect 580252 359776 580358 359786
rect 491168 359028 491288 359050
rect 491168 357440 491170 359028
rect 491286 357440 491288 359028
rect 491168 357418 491288 357440
rect 494928 359028 495048 359050
rect 494928 357440 494930 359028
rect 495046 357440 495048 359028
rect 494928 357418 495048 357440
rect 498688 359028 498808 359050
rect 498688 357440 498690 359028
rect 498806 357440 498808 359028
rect 498688 357418 498808 357440
rect 502448 359028 502568 359050
rect 502448 357440 502450 359028
rect 502566 357440 502568 359028
rect 502448 357418 502568 357440
rect 506208 359028 506328 359050
rect 506208 357440 506210 359028
rect 506326 357440 506328 359028
rect 506208 357418 506328 357440
rect 509968 359028 510088 359050
rect 509968 357440 509970 359028
rect 510086 357440 510088 359028
rect 509968 357418 510088 357440
rect 513728 359028 513848 359050
rect 513728 357440 513730 359028
rect 513846 357440 513848 359028
rect 513728 357418 513848 357440
rect 517488 359028 517608 359050
rect 517488 357440 517490 359028
rect 517606 357440 517608 359028
rect 517488 357418 517608 357440
rect 521248 359028 521368 359050
rect 521248 357440 521250 359028
rect 521366 357440 521368 359028
rect 521248 357418 521368 357440
rect 525008 359028 525128 359050
rect 525008 357440 525010 359028
rect 525126 357440 525128 359028
rect 525008 357418 525128 357440
rect 528768 359028 528888 359050
rect 528768 357440 528770 359028
rect 528886 357440 528888 359028
rect 528768 357418 528888 357440
rect 532528 359028 532648 359050
rect 532528 357440 532530 359028
rect 532646 357440 532648 359028
rect 532528 357418 532648 357440
rect 536288 359028 536408 359050
rect 536288 357440 536290 359028
rect 536406 357440 536408 359028
rect 559712 358052 559920 358062
rect 559712 357834 559920 357844
rect 573540 357920 573878 357930
rect 573540 357584 573878 357594
rect 536288 357418 536408 357440
rect 508362 356582 508652 356592
rect 508362 356436 508652 356446
rect 566126 313804 566346 313814
rect 566126 313600 566346 313610
rect 580758 313770 580944 313780
rect 580758 313592 580944 313602
rect 559652 311744 559860 311754
rect 559652 311526 559860 311536
rect 573492 311700 573834 311710
rect 573492 311410 573834 311420
<< via2 >>
rect 566186 494126 566408 494310
rect 580856 494136 581040 494348
rect 559802 492324 560012 492536
rect 573564 491888 573874 492160
rect 491200 413970 491256 414026
rect 491200 413890 491256 413946
rect 491200 413810 491256 413866
rect 491200 413730 491256 413786
rect 491200 413650 491256 413706
rect 491200 413570 491256 413626
rect 491200 413490 491256 413546
rect 491200 413410 491256 413466
rect 491200 413330 491256 413386
rect 491200 413250 491256 413306
rect 491200 413170 491256 413226
rect 491200 413090 491256 413146
rect 491200 413010 491256 413066
rect 491200 412930 491256 412986
rect 491200 412850 491256 412906
rect 491200 412770 491256 412826
rect 491200 412690 491256 412746
rect 491200 412610 491256 412666
rect 491200 412530 491256 412586
rect 491200 412450 491256 412506
rect 494960 413970 495016 414026
rect 494960 413890 495016 413946
rect 494960 413810 495016 413866
rect 494960 413730 495016 413786
rect 494960 413650 495016 413706
rect 494960 413570 495016 413626
rect 494960 413490 495016 413546
rect 494960 413410 495016 413466
rect 494960 413330 495016 413386
rect 494960 413250 495016 413306
rect 494960 413170 495016 413226
rect 494960 413090 495016 413146
rect 494960 413010 495016 413066
rect 494960 412930 495016 412986
rect 494960 412850 495016 412906
rect 494960 412770 495016 412826
rect 494960 412690 495016 412746
rect 494960 412610 495016 412666
rect 494960 412530 495016 412586
rect 494960 412450 495016 412506
rect 498720 413970 498776 414026
rect 498720 413890 498776 413946
rect 498720 413810 498776 413866
rect 498720 413730 498776 413786
rect 498720 413650 498776 413706
rect 498720 413570 498776 413626
rect 498720 413490 498776 413546
rect 498720 413410 498776 413466
rect 498720 413330 498776 413386
rect 498720 413250 498776 413306
rect 498720 413170 498776 413226
rect 498720 413090 498776 413146
rect 498720 413010 498776 413066
rect 498720 412930 498776 412986
rect 498720 412850 498776 412906
rect 498720 412770 498776 412826
rect 498720 412690 498776 412746
rect 498720 412610 498776 412666
rect 498720 412530 498776 412586
rect 498720 412450 498776 412506
rect 502480 413970 502536 414026
rect 502480 413890 502536 413946
rect 502480 413810 502536 413866
rect 502480 413730 502536 413786
rect 502480 413650 502536 413706
rect 502480 413570 502536 413626
rect 502480 413490 502536 413546
rect 502480 413410 502536 413466
rect 502480 413330 502536 413386
rect 502480 413250 502536 413306
rect 502480 413170 502536 413226
rect 502480 413090 502536 413146
rect 502480 413010 502536 413066
rect 502480 412930 502536 412986
rect 502480 412850 502536 412906
rect 502480 412770 502536 412826
rect 502480 412690 502536 412746
rect 502480 412610 502536 412666
rect 502480 412530 502536 412586
rect 502480 412450 502536 412506
rect 506240 413970 506296 414026
rect 506240 413890 506296 413946
rect 506240 413810 506296 413866
rect 506240 413730 506296 413786
rect 506240 413650 506296 413706
rect 506240 413570 506296 413626
rect 506240 413490 506296 413546
rect 506240 413410 506296 413466
rect 506240 413330 506296 413386
rect 506240 413250 506296 413306
rect 506240 413170 506296 413226
rect 506240 413090 506296 413146
rect 506240 413010 506296 413066
rect 506240 412930 506296 412986
rect 506240 412850 506296 412906
rect 506240 412770 506296 412826
rect 506240 412690 506296 412746
rect 506240 412610 506296 412666
rect 506240 412530 506296 412586
rect 506240 412450 506296 412506
rect 510000 413970 510056 414026
rect 510000 413890 510056 413946
rect 510000 413810 510056 413866
rect 510000 413730 510056 413786
rect 510000 413650 510056 413706
rect 510000 413570 510056 413626
rect 510000 413490 510056 413546
rect 510000 413410 510056 413466
rect 510000 413330 510056 413386
rect 510000 413250 510056 413306
rect 510000 413170 510056 413226
rect 510000 413090 510056 413146
rect 510000 413010 510056 413066
rect 510000 412930 510056 412986
rect 510000 412850 510056 412906
rect 510000 412770 510056 412826
rect 510000 412690 510056 412746
rect 510000 412610 510056 412666
rect 510000 412530 510056 412586
rect 510000 412450 510056 412506
rect 513760 413970 513816 414026
rect 513760 413890 513816 413946
rect 513760 413810 513816 413866
rect 513760 413730 513816 413786
rect 513760 413650 513816 413706
rect 513760 413570 513816 413626
rect 513760 413490 513816 413546
rect 513760 413410 513816 413466
rect 513760 413330 513816 413386
rect 513760 413250 513816 413306
rect 513760 413170 513816 413226
rect 513760 413090 513816 413146
rect 513760 413010 513816 413066
rect 513760 412930 513816 412986
rect 513760 412850 513816 412906
rect 513760 412770 513816 412826
rect 513760 412690 513816 412746
rect 513760 412610 513816 412666
rect 513760 412530 513816 412586
rect 513760 412450 513816 412506
rect 517520 413970 517576 414026
rect 517520 413890 517576 413946
rect 517520 413810 517576 413866
rect 517520 413730 517576 413786
rect 517520 413650 517576 413706
rect 517520 413570 517576 413626
rect 517520 413490 517576 413546
rect 517520 413410 517576 413466
rect 517520 413330 517576 413386
rect 517520 413250 517576 413306
rect 517520 413170 517576 413226
rect 517520 413090 517576 413146
rect 517520 413010 517576 413066
rect 517520 412930 517576 412986
rect 517520 412850 517576 412906
rect 517520 412770 517576 412826
rect 517520 412690 517576 412746
rect 517520 412610 517576 412666
rect 517520 412530 517576 412586
rect 517520 412450 517576 412506
rect 521280 413970 521336 414026
rect 521280 413890 521336 413946
rect 521280 413810 521336 413866
rect 521280 413730 521336 413786
rect 521280 413650 521336 413706
rect 521280 413570 521336 413626
rect 521280 413490 521336 413546
rect 521280 413410 521336 413466
rect 521280 413330 521336 413386
rect 521280 413250 521336 413306
rect 521280 413170 521336 413226
rect 521280 413090 521336 413146
rect 521280 413010 521336 413066
rect 521280 412930 521336 412986
rect 521280 412850 521336 412906
rect 521280 412770 521336 412826
rect 521280 412690 521336 412746
rect 521280 412610 521336 412666
rect 521280 412530 521336 412586
rect 521280 412450 521336 412506
rect 525040 413970 525096 414026
rect 525040 413890 525096 413946
rect 525040 413810 525096 413866
rect 525040 413730 525096 413786
rect 525040 413650 525096 413706
rect 525040 413570 525096 413626
rect 525040 413490 525096 413546
rect 525040 413410 525096 413466
rect 525040 413330 525096 413386
rect 525040 413250 525096 413306
rect 525040 413170 525096 413226
rect 525040 413090 525096 413146
rect 525040 413010 525096 413066
rect 525040 412930 525096 412986
rect 525040 412850 525096 412906
rect 525040 412770 525096 412826
rect 525040 412690 525096 412746
rect 525040 412610 525096 412666
rect 525040 412530 525096 412586
rect 525040 412450 525096 412506
rect 528800 413970 528856 414026
rect 528800 413890 528856 413946
rect 528800 413810 528856 413866
rect 528800 413730 528856 413786
rect 528800 413650 528856 413706
rect 528800 413570 528856 413626
rect 528800 413490 528856 413546
rect 528800 413410 528856 413466
rect 528800 413330 528856 413386
rect 528800 413250 528856 413306
rect 528800 413170 528856 413226
rect 528800 413090 528856 413146
rect 528800 413010 528856 413066
rect 528800 412930 528856 412986
rect 528800 412850 528856 412906
rect 528800 412770 528856 412826
rect 528800 412690 528856 412746
rect 528800 412610 528856 412666
rect 528800 412530 528856 412586
rect 528800 412450 528856 412506
rect 532560 413970 532616 414026
rect 532560 413890 532616 413946
rect 532560 413810 532616 413866
rect 532560 413730 532616 413786
rect 532560 413650 532616 413706
rect 532560 413570 532616 413626
rect 532560 413490 532616 413546
rect 532560 413410 532616 413466
rect 532560 413330 532616 413386
rect 532560 413250 532616 413306
rect 532560 413170 532616 413226
rect 532560 413090 532616 413146
rect 532560 413010 532616 413066
rect 532560 412930 532616 412986
rect 532560 412850 532616 412906
rect 532560 412770 532616 412826
rect 532560 412690 532616 412746
rect 532560 412610 532616 412666
rect 532560 412530 532616 412586
rect 532560 412450 532616 412506
rect 536320 413970 536376 414026
rect 536320 413890 536376 413946
rect 536320 413810 536376 413866
rect 536320 413730 536376 413786
rect 536320 413650 536376 413706
rect 536320 413570 536376 413626
rect 536320 413490 536376 413546
rect 536320 413410 536376 413466
rect 536320 413330 536376 413386
rect 536320 413250 536376 413306
rect 536320 413170 536376 413226
rect 536320 413090 536376 413146
rect 536320 413010 536376 413066
rect 536320 412930 536376 412986
rect 536320 412850 536376 412906
rect 536320 412770 536376 412826
rect 536320 412690 536376 412746
rect 536320 412610 536376 412666
rect 536320 412530 536376 412586
rect 536320 412450 536376 412506
rect 493080 411522 493136 411578
rect 493080 411442 493136 411498
rect 493080 411362 493136 411418
rect 493080 411282 493136 411338
rect 493080 411202 493136 411258
rect 493080 411122 493136 411178
rect 493080 411042 493136 411098
rect 493080 410962 493136 411018
rect 493080 410882 493136 410938
rect 493080 410802 493136 410858
rect 493080 410722 493136 410778
rect 493080 410642 493136 410698
rect 493080 410562 493136 410618
rect 493080 410482 493136 410538
rect 493080 410402 493136 410458
rect 493080 410322 493136 410378
rect 493080 410242 493136 410298
rect 493080 410162 493136 410218
rect 493080 410082 493136 410138
rect 493080 410002 493136 410058
rect 496840 411522 496896 411578
rect 496840 411442 496896 411498
rect 496840 411362 496896 411418
rect 496840 411282 496896 411338
rect 496840 411202 496896 411258
rect 496840 411122 496896 411178
rect 496840 411042 496896 411098
rect 496840 410962 496896 411018
rect 496840 410882 496896 410938
rect 496840 410802 496896 410858
rect 496840 410722 496896 410778
rect 496840 410642 496896 410698
rect 496840 410562 496896 410618
rect 496840 410482 496896 410538
rect 496840 410402 496896 410458
rect 496840 410322 496896 410378
rect 496840 410242 496896 410298
rect 496840 410162 496896 410218
rect 496840 410082 496896 410138
rect 496840 410002 496896 410058
rect 500600 411522 500656 411578
rect 500600 411442 500656 411498
rect 500600 411362 500656 411418
rect 500600 411282 500656 411338
rect 500600 411202 500656 411258
rect 500600 411122 500656 411178
rect 500600 411042 500656 411098
rect 500600 410962 500656 411018
rect 500600 410882 500656 410938
rect 500600 410802 500656 410858
rect 500600 410722 500656 410778
rect 500600 410642 500656 410698
rect 500600 410562 500656 410618
rect 500600 410482 500656 410538
rect 500600 410402 500656 410458
rect 500600 410322 500656 410378
rect 500600 410242 500656 410298
rect 500600 410162 500656 410218
rect 500600 410082 500656 410138
rect 500600 410002 500656 410058
rect 504360 411522 504416 411578
rect 504360 411442 504416 411498
rect 504360 411362 504416 411418
rect 504360 411282 504416 411338
rect 504360 411202 504416 411258
rect 504360 411122 504416 411178
rect 504360 411042 504416 411098
rect 504360 410962 504416 411018
rect 504360 410882 504416 410938
rect 504360 410802 504416 410858
rect 504360 410722 504416 410778
rect 504360 410642 504416 410698
rect 504360 410562 504416 410618
rect 504360 410482 504416 410538
rect 504360 410402 504416 410458
rect 504360 410322 504416 410378
rect 504360 410242 504416 410298
rect 504360 410162 504416 410218
rect 504360 410082 504416 410138
rect 504360 410002 504416 410058
rect 508120 411522 508176 411578
rect 508120 411442 508176 411498
rect 508120 411362 508176 411418
rect 508120 411282 508176 411338
rect 508120 411202 508176 411258
rect 508120 411122 508176 411178
rect 508120 411042 508176 411098
rect 508120 410962 508176 411018
rect 508120 410882 508176 410938
rect 508120 410802 508176 410858
rect 508120 410722 508176 410778
rect 508120 410642 508176 410698
rect 508120 410562 508176 410618
rect 508120 410482 508176 410538
rect 508120 410402 508176 410458
rect 508120 410322 508176 410378
rect 508120 410242 508176 410298
rect 508120 410162 508176 410218
rect 508120 410082 508176 410138
rect 508120 410002 508176 410058
rect 511880 411522 511936 411578
rect 511880 411442 511936 411498
rect 511880 411362 511936 411418
rect 511880 411282 511936 411338
rect 511880 411202 511936 411258
rect 511880 411122 511936 411178
rect 511880 411042 511936 411098
rect 511880 410962 511936 411018
rect 511880 410882 511936 410938
rect 511880 410802 511936 410858
rect 511880 410722 511936 410778
rect 511880 410642 511936 410698
rect 511880 410562 511936 410618
rect 511880 410482 511936 410538
rect 511880 410402 511936 410458
rect 511880 410322 511936 410378
rect 511880 410242 511936 410298
rect 511880 410162 511936 410218
rect 511880 410082 511936 410138
rect 511880 410002 511936 410058
rect 515640 411522 515696 411578
rect 515640 411442 515696 411498
rect 515640 411362 515696 411418
rect 515640 411282 515696 411338
rect 515640 411202 515696 411258
rect 515640 411122 515696 411178
rect 515640 411042 515696 411098
rect 515640 410962 515696 411018
rect 515640 410882 515696 410938
rect 515640 410802 515696 410858
rect 515640 410722 515696 410778
rect 515640 410642 515696 410698
rect 515640 410562 515696 410618
rect 515640 410482 515696 410538
rect 515640 410402 515696 410458
rect 515640 410322 515696 410378
rect 515640 410242 515696 410298
rect 515640 410162 515696 410218
rect 515640 410082 515696 410138
rect 515640 410002 515696 410058
rect 519400 411522 519456 411578
rect 519400 411442 519456 411498
rect 519400 411362 519456 411418
rect 519400 411282 519456 411338
rect 519400 411202 519456 411258
rect 519400 411122 519456 411178
rect 519400 411042 519456 411098
rect 519400 410962 519456 411018
rect 519400 410882 519456 410938
rect 519400 410802 519456 410858
rect 519400 410722 519456 410778
rect 519400 410642 519456 410698
rect 519400 410562 519456 410618
rect 519400 410482 519456 410538
rect 519400 410402 519456 410458
rect 519400 410322 519456 410378
rect 519400 410242 519456 410298
rect 519400 410162 519456 410218
rect 519400 410082 519456 410138
rect 519400 410002 519456 410058
rect 523160 411522 523216 411578
rect 523160 411442 523216 411498
rect 523160 411362 523216 411418
rect 523160 411282 523216 411338
rect 523160 411202 523216 411258
rect 523160 411122 523216 411178
rect 523160 411042 523216 411098
rect 523160 410962 523216 411018
rect 523160 410882 523216 410938
rect 523160 410802 523216 410858
rect 523160 410722 523216 410778
rect 523160 410642 523216 410698
rect 523160 410562 523216 410618
rect 523160 410482 523216 410538
rect 523160 410402 523216 410458
rect 523160 410322 523216 410378
rect 523160 410242 523216 410298
rect 523160 410162 523216 410218
rect 523160 410082 523216 410138
rect 523160 410002 523216 410058
rect 526920 411522 526976 411578
rect 526920 411442 526976 411498
rect 526920 411362 526976 411418
rect 526920 411282 526976 411338
rect 526920 411202 526976 411258
rect 526920 411122 526976 411178
rect 526920 411042 526976 411098
rect 526920 410962 526976 411018
rect 526920 410882 526976 410938
rect 526920 410802 526976 410858
rect 526920 410722 526976 410778
rect 526920 410642 526976 410698
rect 526920 410562 526976 410618
rect 526920 410482 526976 410538
rect 526920 410402 526976 410458
rect 526920 410322 526976 410378
rect 526920 410242 526976 410298
rect 526920 410162 526976 410218
rect 526920 410082 526976 410138
rect 526920 410002 526976 410058
rect 530680 411522 530736 411578
rect 530680 411442 530736 411498
rect 530680 411362 530736 411418
rect 530680 411282 530736 411338
rect 530680 411202 530736 411258
rect 530680 411122 530736 411178
rect 530680 411042 530736 411098
rect 530680 410962 530736 411018
rect 530680 410882 530736 410938
rect 530680 410802 530736 410858
rect 530680 410722 530736 410778
rect 530680 410642 530736 410698
rect 530680 410562 530736 410618
rect 530680 410482 530736 410538
rect 530680 410402 530736 410458
rect 530680 410322 530736 410378
rect 530680 410242 530736 410298
rect 530680 410162 530736 410218
rect 530680 410082 530736 410138
rect 530680 410002 530736 410058
rect 534440 411522 534496 411578
rect 534440 411442 534496 411498
rect 534440 411362 534496 411418
rect 534440 411282 534496 411338
rect 534440 411202 534496 411258
rect 534440 411122 534496 411178
rect 534440 411042 534496 411098
rect 534440 410962 534496 411018
rect 534440 410882 534496 410938
rect 534440 410802 534496 410858
rect 534440 410722 534496 410778
rect 534440 410642 534496 410698
rect 534440 410562 534496 410618
rect 534440 410482 534496 410538
rect 534440 410402 534496 410458
rect 534440 410322 534496 410378
rect 534440 410242 534496 410298
rect 534440 410162 534496 410218
rect 534440 410082 534496 410138
rect 534440 410002 534496 410058
rect 493350 408950 493406 409006
rect 493350 408870 493406 408926
rect 494770 408908 494826 408964
rect 497110 408950 497166 409006
rect 497110 408870 497166 408926
rect 498530 408908 498586 408964
rect 500870 408558 500926 408614
rect 500870 408478 500926 408534
rect 502290 408516 502346 408572
rect 498710 406654 498766 406656
rect 498710 406602 498752 406654
rect 498752 406602 498766 406654
rect 498710 406600 498766 406602
rect 566256 405258 566462 405476
rect 580074 405292 580182 405402
rect 559736 403192 559926 403368
rect 573538 402980 573888 403312
rect 504810 402000 504866 402056
rect 493350 401502 493406 401558
rect 493350 401422 493406 401478
rect 494770 401460 494826 401516
rect 498588 400398 498644 400400
rect 498588 400346 498600 400398
rect 498600 400346 498644 400398
rect 498588 400344 498644 400346
rect 498222 399884 498278 399940
rect 500870 399738 500926 399794
rect 500870 399658 500926 399714
rect 502290 399696 502346 399752
rect 502370 399424 502426 399480
rect 494928 397270 494984 397272
rect 494928 397218 494944 397270
rect 494944 397218 494984 397270
rect 494928 397216 494984 397218
rect 500662 392708 500718 392764
rect 498588 391144 498644 391200
rect 541952 389388 542058 389470
rect 508390 388664 508446 388720
rect 508390 388584 508446 388640
rect 509810 388622 509866 388678
rect 505054 385494 505110 385496
rect 505054 385442 505076 385494
rect 505076 385442 505110 385494
rect 505054 385440 505110 385442
rect 516278 385494 516334 385496
rect 516278 385442 516296 385494
rect 516296 385442 516334 385494
rect 516278 385440 516334 385442
rect 504630 384940 504686 384996
rect 504630 384860 504686 384916
rect 506050 384898 506106 384954
rect 512150 384940 512206 384996
rect 512150 384860 512206 384916
rect 513570 384898 513626 384954
rect 515910 384940 515966 384996
rect 515910 384860 515966 384916
rect 517330 384898 517386 384954
rect 504444 381538 504500 381540
rect 504444 381486 504448 381538
rect 504448 381486 504500 381538
rect 504444 381484 504500 381486
rect 508226 381484 508282 381540
rect 511886 381538 511942 381540
rect 511886 381486 511928 381538
rect 511928 381486 511942 381538
rect 511886 381484 511942 381486
rect 515668 381484 515724 381540
rect 508390 381216 508446 381272
rect 508390 381136 508446 381192
rect 509810 381174 509866 381230
rect 541958 380564 542066 380644
rect 506030 377398 506086 377400
rect 506030 377346 506080 377398
rect 506080 377346 506086 377398
rect 506030 377344 506086 377346
rect 493080 361414 493136 361470
rect 493080 361334 493136 361390
rect 493080 361254 493136 361310
rect 493080 361174 493136 361230
rect 493080 361094 493136 361150
rect 493080 361014 493136 361070
rect 493080 360934 493136 360990
rect 493080 360854 493136 360910
rect 493080 360774 493136 360830
rect 493080 360694 493136 360750
rect 493080 360614 493136 360670
rect 493080 360534 493136 360590
rect 493080 360454 493136 360510
rect 493080 360374 493136 360430
rect 493080 360294 493136 360350
rect 493080 360214 493136 360270
rect 493080 360134 493136 360190
rect 493080 360054 493136 360110
rect 493080 359974 493136 360030
rect 493080 359894 493136 359950
rect 496840 361414 496896 361470
rect 496840 361334 496896 361390
rect 496840 361254 496896 361310
rect 496840 361174 496896 361230
rect 496840 361094 496896 361150
rect 496840 361014 496896 361070
rect 496840 360934 496896 360990
rect 496840 360854 496896 360910
rect 496840 360774 496896 360830
rect 496840 360694 496896 360750
rect 496840 360614 496896 360670
rect 496840 360534 496896 360590
rect 496840 360454 496896 360510
rect 496840 360374 496896 360430
rect 496840 360294 496896 360350
rect 496840 360214 496896 360270
rect 496840 360134 496896 360190
rect 496840 360054 496896 360110
rect 496840 359974 496896 360030
rect 496840 359894 496896 359950
rect 500600 361414 500656 361470
rect 500600 361334 500656 361390
rect 500600 361254 500656 361310
rect 500600 361174 500656 361230
rect 500600 361094 500656 361150
rect 500600 361014 500656 361070
rect 500600 360934 500656 360990
rect 500600 360854 500656 360910
rect 500600 360774 500656 360830
rect 500600 360694 500656 360750
rect 500600 360614 500656 360670
rect 500600 360534 500656 360590
rect 500600 360454 500656 360510
rect 500600 360374 500656 360430
rect 500600 360294 500656 360350
rect 500600 360214 500656 360270
rect 500600 360134 500656 360190
rect 500600 360054 500656 360110
rect 500600 359974 500656 360030
rect 500600 359894 500656 359950
rect 504360 361414 504416 361470
rect 504360 361334 504416 361390
rect 504360 361254 504416 361310
rect 504360 361174 504416 361230
rect 504360 361094 504416 361150
rect 504360 361014 504416 361070
rect 504360 360934 504416 360990
rect 504360 360854 504416 360910
rect 504360 360774 504416 360830
rect 504360 360694 504416 360750
rect 504360 360614 504416 360670
rect 504360 360534 504416 360590
rect 504360 360454 504416 360510
rect 504360 360374 504416 360430
rect 504360 360294 504416 360350
rect 504360 360214 504416 360270
rect 504360 360134 504416 360190
rect 504360 360054 504416 360110
rect 504360 359974 504416 360030
rect 504360 359894 504416 359950
rect 508120 361414 508176 361470
rect 508120 361334 508176 361390
rect 508120 361254 508176 361310
rect 508120 361174 508176 361230
rect 508120 361094 508176 361150
rect 508120 361014 508176 361070
rect 508120 360934 508176 360990
rect 508120 360854 508176 360910
rect 508120 360774 508176 360830
rect 508120 360694 508176 360750
rect 508120 360614 508176 360670
rect 508120 360534 508176 360590
rect 508120 360454 508176 360510
rect 508120 360374 508176 360430
rect 508120 360294 508176 360350
rect 508120 360214 508176 360270
rect 508120 360134 508176 360190
rect 508120 360054 508176 360110
rect 508120 359974 508176 360030
rect 508120 359894 508176 359950
rect 511880 361414 511936 361470
rect 511880 361334 511936 361390
rect 511880 361254 511936 361310
rect 511880 361174 511936 361230
rect 511880 361094 511936 361150
rect 511880 361014 511936 361070
rect 511880 360934 511936 360990
rect 511880 360854 511936 360910
rect 511880 360774 511936 360830
rect 511880 360694 511936 360750
rect 511880 360614 511936 360670
rect 511880 360534 511936 360590
rect 511880 360454 511936 360510
rect 511880 360374 511936 360430
rect 511880 360294 511936 360350
rect 511880 360214 511936 360270
rect 511880 360134 511936 360190
rect 511880 360054 511936 360110
rect 511880 359974 511936 360030
rect 511880 359894 511936 359950
rect 515640 361414 515696 361470
rect 515640 361334 515696 361390
rect 515640 361254 515696 361310
rect 515640 361174 515696 361230
rect 515640 361094 515696 361150
rect 515640 361014 515696 361070
rect 515640 360934 515696 360990
rect 515640 360854 515696 360910
rect 515640 360774 515696 360830
rect 515640 360694 515696 360750
rect 515640 360614 515696 360670
rect 515640 360534 515696 360590
rect 515640 360454 515696 360510
rect 515640 360374 515696 360430
rect 515640 360294 515696 360350
rect 515640 360214 515696 360270
rect 515640 360134 515696 360190
rect 515640 360054 515696 360110
rect 515640 359974 515696 360030
rect 515640 359894 515696 359950
rect 519400 361414 519456 361470
rect 519400 361334 519456 361390
rect 519400 361254 519456 361310
rect 519400 361174 519456 361230
rect 519400 361094 519456 361150
rect 519400 361014 519456 361070
rect 519400 360934 519456 360990
rect 519400 360854 519456 360910
rect 519400 360774 519456 360830
rect 519400 360694 519456 360750
rect 519400 360614 519456 360670
rect 519400 360534 519456 360590
rect 519400 360454 519456 360510
rect 519400 360374 519456 360430
rect 519400 360294 519456 360350
rect 519400 360214 519456 360270
rect 519400 360134 519456 360190
rect 519400 360054 519456 360110
rect 519400 359974 519456 360030
rect 519400 359894 519456 359950
rect 523160 361414 523216 361470
rect 523160 361334 523216 361390
rect 523160 361254 523216 361310
rect 523160 361174 523216 361230
rect 523160 361094 523216 361150
rect 523160 361014 523216 361070
rect 523160 360934 523216 360990
rect 523160 360854 523216 360910
rect 523160 360774 523216 360830
rect 523160 360694 523216 360750
rect 523160 360614 523216 360670
rect 523160 360534 523216 360590
rect 523160 360454 523216 360510
rect 523160 360374 523216 360430
rect 523160 360294 523216 360350
rect 523160 360214 523216 360270
rect 523160 360134 523216 360190
rect 523160 360054 523216 360110
rect 523160 359974 523216 360030
rect 523160 359894 523216 359950
rect 526920 361414 526976 361470
rect 526920 361334 526976 361390
rect 526920 361254 526976 361310
rect 526920 361174 526976 361230
rect 526920 361094 526976 361150
rect 526920 361014 526976 361070
rect 526920 360934 526976 360990
rect 526920 360854 526976 360910
rect 526920 360774 526976 360830
rect 526920 360694 526976 360750
rect 526920 360614 526976 360670
rect 526920 360534 526976 360590
rect 526920 360454 526976 360510
rect 526920 360374 526976 360430
rect 526920 360294 526976 360350
rect 526920 360214 526976 360270
rect 526920 360134 526976 360190
rect 526920 360054 526976 360110
rect 526920 359974 526976 360030
rect 526920 359894 526976 359950
rect 530680 361414 530736 361470
rect 530680 361334 530736 361390
rect 530680 361254 530736 361310
rect 530680 361174 530736 361230
rect 530680 361094 530736 361150
rect 530680 361014 530736 361070
rect 530680 360934 530736 360990
rect 530680 360854 530736 360910
rect 530680 360774 530736 360830
rect 530680 360694 530736 360750
rect 530680 360614 530736 360670
rect 530680 360534 530736 360590
rect 530680 360454 530736 360510
rect 530680 360374 530736 360430
rect 530680 360294 530736 360350
rect 530680 360214 530736 360270
rect 530680 360134 530736 360190
rect 530680 360054 530736 360110
rect 530680 359974 530736 360030
rect 530680 359894 530736 359950
rect 534440 361414 534496 361470
rect 534440 361334 534496 361390
rect 534440 361254 534496 361310
rect 534440 361174 534496 361230
rect 534440 361094 534496 361150
rect 534440 361014 534496 361070
rect 534440 360934 534496 360990
rect 534440 360854 534496 360910
rect 534440 360774 534496 360830
rect 534440 360694 534496 360750
rect 534440 360614 534496 360670
rect 534440 360534 534496 360590
rect 534440 360454 534496 360510
rect 534440 360374 534496 360430
rect 534440 360294 534496 360350
rect 534440 360214 534496 360270
rect 534440 360134 534496 360190
rect 534440 360054 534496 360110
rect 534440 359974 534496 360030
rect 534440 359894 534496 359950
rect 566274 359786 566500 359978
rect 580252 359786 580358 359906
rect 491200 358966 491256 359022
rect 491200 358886 491256 358942
rect 491200 358806 491256 358862
rect 491200 358726 491256 358782
rect 491200 358646 491256 358702
rect 491200 358566 491256 358622
rect 491200 358486 491256 358542
rect 491200 358406 491256 358462
rect 491200 358326 491256 358382
rect 491200 358246 491256 358302
rect 491200 358166 491256 358222
rect 491200 358086 491256 358142
rect 491200 358006 491256 358062
rect 491200 357926 491256 357982
rect 491200 357846 491256 357902
rect 491200 357766 491256 357822
rect 491200 357686 491256 357742
rect 491200 357606 491256 357662
rect 491200 357526 491256 357582
rect 491200 357446 491256 357502
rect 494960 358966 495016 359022
rect 494960 358886 495016 358942
rect 494960 358806 495016 358862
rect 494960 358726 495016 358782
rect 494960 358646 495016 358702
rect 494960 358566 495016 358622
rect 494960 358486 495016 358542
rect 494960 358406 495016 358462
rect 494960 358326 495016 358382
rect 494960 358246 495016 358302
rect 494960 358166 495016 358222
rect 494960 358086 495016 358142
rect 494960 358006 495016 358062
rect 494960 357926 495016 357982
rect 494960 357846 495016 357902
rect 494960 357766 495016 357822
rect 494960 357686 495016 357742
rect 494960 357606 495016 357662
rect 494960 357526 495016 357582
rect 494960 357446 495016 357502
rect 498720 358966 498776 359022
rect 498720 358886 498776 358942
rect 498720 358806 498776 358862
rect 498720 358726 498776 358782
rect 498720 358646 498776 358702
rect 498720 358566 498776 358622
rect 498720 358486 498776 358542
rect 498720 358406 498776 358462
rect 498720 358326 498776 358382
rect 498720 358246 498776 358302
rect 498720 358166 498776 358222
rect 498720 358086 498776 358142
rect 498720 358006 498776 358062
rect 498720 357926 498776 357982
rect 498720 357846 498776 357902
rect 498720 357766 498776 357822
rect 498720 357686 498776 357742
rect 498720 357606 498776 357662
rect 498720 357526 498776 357582
rect 498720 357446 498776 357502
rect 502480 358966 502536 359022
rect 502480 358886 502536 358942
rect 502480 358806 502536 358862
rect 502480 358726 502536 358782
rect 502480 358646 502536 358702
rect 502480 358566 502536 358622
rect 502480 358486 502536 358542
rect 502480 358406 502536 358462
rect 502480 358326 502536 358382
rect 502480 358246 502536 358302
rect 502480 358166 502536 358222
rect 502480 358086 502536 358142
rect 502480 358006 502536 358062
rect 502480 357926 502536 357982
rect 502480 357846 502536 357902
rect 502480 357766 502536 357822
rect 502480 357686 502536 357742
rect 502480 357606 502536 357662
rect 502480 357526 502536 357582
rect 502480 357446 502536 357502
rect 506240 358966 506296 359022
rect 506240 358886 506296 358942
rect 506240 358806 506296 358862
rect 506240 358726 506296 358782
rect 506240 358646 506296 358702
rect 506240 358566 506296 358622
rect 506240 358486 506296 358542
rect 506240 358406 506296 358462
rect 506240 358326 506296 358382
rect 506240 358246 506296 358302
rect 506240 358166 506296 358222
rect 506240 358086 506296 358142
rect 506240 358006 506296 358062
rect 506240 357926 506296 357982
rect 506240 357846 506296 357902
rect 506240 357766 506296 357822
rect 506240 357686 506296 357742
rect 506240 357606 506296 357662
rect 506240 357526 506296 357582
rect 506240 357446 506296 357502
rect 510000 358966 510056 359022
rect 510000 358886 510056 358942
rect 510000 358806 510056 358862
rect 510000 358726 510056 358782
rect 510000 358646 510056 358702
rect 510000 358566 510056 358622
rect 510000 358486 510056 358542
rect 510000 358406 510056 358462
rect 510000 358326 510056 358382
rect 510000 358246 510056 358302
rect 510000 358166 510056 358222
rect 510000 358086 510056 358142
rect 510000 358006 510056 358062
rect 510000 357926 510056 357982
rect 510000 357846 510056 357902
rect 510000 357766 510056 357822
rect 510000 357686 510056 357742
rect 510000 357606 510056 357662
rect 510000 357526 510056 357582
rect 510000 357446 510056 357502
rect 513760 358966 513816 359022
rect 513760 358886 513816 358942
rect 513760 358806 513816 358862
rect 513760 358726 513816 358782
rect 513760 358646 513816 358702
rect 513760 358566 513816 358622
rect 513760 358486 513816 358542
rect 513760 358406 513816 358462
rect 513760 358326 513816 358382
rect 513760 358246 513816 358302
rect 513760 358166 513816 358222
rect 513760 358086 513816 358142
rect 513760 358006 513816 358062
rect 513760 357926 513816 357982
rect 513760 357846 513816 357902
rect 513760 357766 513816 357822
rect 513760 357686 513816 357742
rect 513760 357606 513816 357662
rect 513760 357526 513816 357582
rect 513760 357446 513816 357502
rect 517520 358966 517576 359022
rect 517520 358886 517576 358942
rect 517520 358806 517576 358862
rect 517520 358726 517576 358782
rect 517520 358646 517576 358702
rect 517520 358566 517576 358622
rect 517520 358486 517576 358542
rect 517520 358406 517576 358462
rect 517520 358326 517576 358382
rect 517520 358246 517576 358302
rect 517520 358166 517576 358222
rect 517520 358086 517576 358142
rect 517520 358006 517576 358062
rect 517520 357926 517576 357982
rect 517520 357846 517576 357902
rect 517520 357766 517576 357822
rect 517520 357686 517576 357742
rect 517520 357606 517576 357662
rect 517520 357526 517576 357582
rect 517520 357446 517576 357502
rect 521280 358966 521336 359022
rect 521280 358886 521336 358942
rect 521280 358806 521336 358862
rect 521280 358726 521336 358782
rect 521280 358646 521336 358702
rect 521280 358566 521336 358622
rect 521280 358486 521336 358542
rect 521280 358406 521336 358462
rect 521280 358326 521336 358382
rect 521280 358246 521336 358302
rect 521280 358166 521336 358222
rect 521280 358086 521336 358142
rect 521280 358006 521336 358062
rect 521280 357926 521336 357982
rect 521280 357846 521336 357902
rect 521280 357766 521336 357822
rect 521280 357686 521336 357742
rect 521280 357606 521336 357662
rect 521280 357526 521336 357582
rect 521280 357446 521336 357502
rect 525040 358966 525096 359022
rect 525040 358886 525096 358942
rect 525040 358806 525096 358862
rect 525040 358726 525096 358782
rect 525040 358646 525096 358702
rect 525040 358566 525096 358622
rect 525040 358486 525096 358542
rect 525040 358406 525096 358462
rect 525040 358326 525096 358382
rect 525040 358246 525096 358302
rect 525040 358166 525096 358222
rect 525040 358086 525096 358142
rect 525040 358006 525096 358062
rect 525040 357926 525096 357982
rect 525040 357846 525096 357902
rect 525040 357766 525096 357822
rect 525040 357686 525096 357742
rect 525040 357606 525096 357662
rect 525040 357526 525096 357582
rect 525040 357446 525096 357502
rect 528800 358966 528856 359022
rect 528800 358886 528856 358942
rect 528800 358806 528856 358862
rect 528800 358726 528856 358782
rect 528800 358646 528856 358702
rect 528800 358566 528856 358622
rect 528800 358486 528856 358542
rect 528800 358406 528856 358462
rect 528800 358326 528856 358382
rect 528800 358246 528856 358302
rect 528800 358166 528856 358222
rect 528800 358086 528856 358142
rect 528800 358006 528856 358062
rect 528800 357926 528856 357982
rect 528800 357846 528856 357902
rect 528800 357766 528856 357822
rect 528800 357686 528856 357742
rect 528800 357606 528856 357662
rect 528800 357526 528856 357582
rect 528800 357446 528856 357502
rect 532560 358966 532616 359022
rect 532560 358886 532616 358942
rect 532560 358806 532616 358862
rect 532560 358726 532616 358782
rect 532560 358646 532616 358702
rect 532560 358566 532616 358622
rect 532560 358486 532616 358542
rect 532560 358406 532616 358462
rect 532560 358326 532616 358382
rect 532560 358246 532616 358302
rect 532560 358166 532616 358222
rect 532560 358086 532616 358142
rect 532560 358006 532616 358062
rect 532560 357926 532616 357982
rect 532560 357846 532616 357902
rect 532560 357766 532616 357822
rect 532560 357686 532616 357742
rect 532560 357606 532616 357662
rect 532560 357526 532616 357582
rect 532560 357446 532616 357502
rect 536320 358966 536376 359022
rect 536320 358886 536376 358942
rect 536320 358806 536376 358862
rect 536320 358726 536376 358782
rect 536320 358646 536376 358702
rect 536320 358566 536376 358622
rect 536320 358486 536376 358542
rect 536320 358406 536376 358462
rect 536320 358326 536376 358382
rect 536320 358246 536376 358302
rect 536320 358166 536376 358222
rect 536320 358086 536376 358142
rect 536320 358006 536376 358062
rect 536320 357926 536376 357982
rect 536320 357846 536376 357902
rect 536320 357766 536376 357822
rect 536320 357686 536376 357742
rect 536320 357606 536376 357662
rect 536320 357526 536376 357582
rect 536320 357446 536376 357502
rect 559712 357844 559920 358052
rect 573540 357594 573878 357920
rect 508362 356446 508652 356582
rect 566126 313610 566346 313804
rect 580758 313602 580944 313770
rect 559652 311536 559860 311744
rect 573492 311420 573834 311700
<< metal3 >>
rect 413300 698232 418436 703282
rect 465296 698476 470432 703526
rect 510560 701276 515394 703604
rect 510552 701180 515394 701276
rect 510552 700092 515386 701180
rect 510552 699264 515392 700092
rect 510538 697668 515392 699264
rect 510538 697378 515372 697668
rect 510538 696840 510704 697378
rect 510560 689882 510704 696840
rect 515202 689882 515372 697378
rect 510560 689666 515372 689882
rect 520554 697354 525388 703122
rect 566500 698354 571636 703404
rect 520554 689858 520704 697354
rect 525202 689858 525388 697354
rect 520554 689727 525388 689858
rect 577256 677954 582392 683004
rect 567105 644596 581232 644606
rect 567105 644324 582918 644596
rect 567105 640080 567306 644324
rect 573722 640080 582918 644324
rect 567105 639760 582918 640080
rect 567308 634256 583176 634588
rect 567296 630012 567306 634256
rect 573722 630012 583176 634256
rect 567308 629752 583176 630012
rect 580846 494348 581050 494353
rect 566148 494310 566454 494332
rect 566148 494248 566186 494310
rect 501828 494126 566186 494248
rect 566408 494248 566454 494310
rect 580846 494248 580856 494348
rect 566408 494136 580856 494248
rect 581040 494248 581050 494348
rect 581040 494136 583862 494248
rect 566408 494126 583862 494136
rect 501828 494124 583862 494126
rect 501828 415012 501952 494124
rect 566148 494090 566454 494124
rect 559792 492536 560022 492541
rect 559792 492324 559802 492536
rect 560012 492324 560022 492536
rect 559792 492319 560022 492324
rect 573554 492160 573884 492165
rect 573554 491888 573564 492160
rect 573874 491888 573884 492160
rect 573554 491883 573884 491888
rect 501026 414806 501952 415012
rect 491168 414030 491288 414054
rect 491168 413966 491196 414030
rect 491260 413966 491288 414030
rect 491168 413950 491288 413966
rect 491168 413886 491196 413950
rect 491260 413886 491288 413950
rect 491168 413870 491288 413886
rect 491168 413806 491196 413870
rect 491260 413806 491288 413870
rect 491168 413790 491288 413806
rect 491168 413726 491196 413790
rect 491260 413726 491288 413790
rect 491168 413710 491288 413726
rect 491168 413646 491196 413710
rect 491260 413646 491288 413710
rect 491168 413630 491288 413646
rect 491168 413566 491196 413630
rect 491260 413566 491288 413630
rect 491168 413550 491288 413566
rect 491168 413486 491196 413550
rect 491260 413486 491288 413550
rect 491168 413470 491288 413486
rect 491168 413406 491196 413470
rect 491260 413406 491288 413470
rect 491168 413390 491288 413406
rect 491168 413326 491196 413390
rect 491260 413326 491288 413390
rect 491168 413310 491288 413326
rect 491168 413246 491196 413310
rect 491260 413246 491288 413310
rect 491168 413230 491288 413246
rect 491168 413166 491196 413230
rect 491260 413166 491288 413230
rect 491168 413150 491288 413166
rect 491168 413086 491196 413150
rect 491260 413086 491288 413150
rect 491168 413070 491288 413086
rect 491168 413006 491196 413070
rect 491260 413006 491288 413070
rect 491168 412990 491288 413006
rect 491168 412926 491196 412990
rect 491260 412926 491288 412990
rect 491168 412910 491288 412926
rect 491168 412846 491196 412910
rect 491260 412846 491288 412910
rect 491168 412830 491288 412846
rect 491168 412766 491196 412830
rect 491260 412766 491288 412830
rect 491168 412750 491288 412766
rect 491168 412686 491196 412750
rect 491260 412686 491288 412750
rect 491168 412670 491288 412686
rect 491168 412606 491196 412670
rect 491260 412606 491288 412670
rect 491168 412590 491288 412606
rect 491168 412526 491196 412590
rect 491260 412526 491288 412590
rect 491168 412510 491288 412526
rect 491168 412446 491196 412510
rect 491260 412446 491288 412510
rect 491168 412422 491288 412446
rect 494928 414030 495048 414054
rect 494928 413966 494956 414030
rect 495020 413966 495048 414030
rect 494928 413950 495048 413966
rect 494928 413886 494956 413950
rect 495020 413886 495048 413950
rect 494928 413870 495048 413886
rect 494928 413806 494956 413870
rect 495020 413806 495048 413870
rect 494928 413790 495048 413806
rect 494928 413726 494956 413790
rect 495020 413726 495048 413790
rect 494928 413710 495048 413726
rect 494928 413646 494956 413710
rect 495020 413646 495048 413710
rect 494928 413630 495048 413646
rect 494928 413566 494956 413630
rect 495020 413566 495048 413630
rect 494928 413550 495048 413566
rect 494928 413486 494956 413550
rect 495020 413486 495048 413550
rect 494928 413470 495048 413486
rect 494928 413406 494956 413470
rect 495020 413406 495048 413470
rect 494928 413390 495048 413406
rect 494928 413326 494956 413390
rect 495020 413326 495048 413390
rect 494928 413310 495048 413326
rect 494928 413246 494956 413310
rect 495020 413246 495048 413310
rect 494928 413230 495048 413246
rect 494928 413166 494956 413230
rect 495020 413166 495048 413230
rect 494928 413150 495048 413166
rect 494928 413086 494956 413150
rect 495020 413086 495048 413150
rect 494928 413070 495048 413086
rect 494928 413006 494956 413070
rect 495020 413006 495048 413070
rect 494928 412990 495048 413006
rect 494928 412926 494956 412990
rect 495020 412926 495048 412990
rect 494928 412910 495048 412926
rect 494928 412846 494956 412910
rect 495020 412846 495048 412910
rect 494928 412830 495048 412846
rect 494928 412766 494956 412830
rect 495020 412766 495048 412830
rect 494928 412750 495048 412766
rect 494928 412686 494956 412750
rect 495020 412686 495048 412750
rect 494928 412670 495048 412686
rect 494928 412606 494956 412670
rect 495020 412606 495048 412670
rect 494928 412590 495048 412606
rect 494928 412526 494956 412590
rect 495020 412526 495048 412590
rect 494928 412510 495048 412526
rect 494928 412446 494956 412510
rect 495020 412446 495048 412510
rect 494928 412422 495048 412446
rect 498688 414030 498808 414054
rect 498688 413966 498716 414030
rect 498780 413966 498808 414030
rect 498688 413950 498808 413966
rect 498688 413886 498716 413950
rect 498780 413886 498808 413950
rect 498688 413870 498808 413886
rect 498688 413806 498716 413870
rect 498780 413806 498808 413870
rect 498688 413790 498808 413806
rect 498688 413726 498716 413790
rect 498780 413726 498808 413790
rect 498688 413710 498808 413726
rect 498688 413646 498716 413710
rect 498780 413646 498808 413710
rect 498688 413630 498808 413646
rect 498688 413566 498716 413630
rect 498780 413566 498808 413630
rect 498688 413550 498808 413566
rect 498688 413486 498716 413550
rect 498780 413486 498808 413550
rect 498688 413470 498808 413486
rect 498688 413406 498716 413470
rect 498780 413406 498808 413470
rect 498688 413390 498808 413406
rect 498688 413326 498716 413390
rect 498780 413326 498808 413390
rect 498688 413310 498808 413326
rect 498688 413246 498716 413310
rect 498780 413246 498808 413310
rect 498688 413230 498808 413246
rect 498688 413166 498716 413230
rect 498780 413166 498808 413230
rect 498688 413150 498808 413166
rect 498688 413086 498716 413150
rect 498780 413086 498808 413150
rect 498688 413070 498808 413086
rect 498688 413006 498716 413070
rect 498780 413006 498808 413070
rect 498688 412990 498808 413006
rect 498688 412926 498716 412990
rect 498780 412926 498808 412990
rect 498688 412910 498808 412926
rect 498688 412846 498716 412910
rect 498780 412846 498808 412910
rect 498688 412830 498808 412846
rect 498688 412766 498716 412830
rect 498780 412766 498808 412830
rect 498688 412750 498808 412766
rect 498688 412686 498716 412750
rect 498780 412686 498808 412750
rect 498688 412670 498808 412686
rect 498688 412606 498716 412670
rect 498780 412606 498808 412670
rect 498688 412590 498808 412606
rect 498688 412526 498716 412590
rect 498780 412526 498808 412590
rect 498688 412510 498808 412526
rect 498688 412446 498716 412510
rect 498780 412446 498808 412510
rect 498688 412422 498808 412446
rect 493048 411582 493168 411606
rect 493048 411518 493076 411582
rect 493140 411518 493168 411582
rect 493048 411502 493168 411518
rect 493048 411438 493076 411502
rect 493140 411438 493168 411502
rect 493048 411422 493168 411438
rect 493048 411358 493076 411422
rect 493140 411358 493168 411422
rect 493048 411342 493168 411358
rect 493048 411278 493076 411342
rect 493140 411278 493168 411342
rect 493048 411262 493168 411278
rect 493048 411198 493076 411262
rect 493140 411198 493168 411262
rect 493048 411182 493168 411198
rect 493048 411118 493076 411182
rect 493140 411118 493168 411182
rect 493048 411102 493168 411118
rect 493048 411038 493076 411102
rect 493140 411038 493168 411102
rect 493048 411022 493168 411038
rect 493048 410958 493076 411022
rect 493140 410958 493168 411022
rect 493048 410942 493168 410958
rect 493048 410878 493076 410942
rect 493140 410878 493168 410942
rect 493048 410862 493168 410878
rect 493048 410798 493076 410862
rect 493140 410798 493168 410862
rect 493048 410782 493168 410798
rect 493048 410718 493076 410782
rect 493140 410718 493168 410782
rect 493048 410702 493168 410718
rect 493048 410638 493076 410702
rect 493140 410638 493168 410702
rect 493048 410622 493168 410638
rect 493048 410558 493076 410622
rect 493140 410558 493168 410622
rect 493048 410542 493168 410558
rect 493048 410478 493076 410542
rect 493140 410478 493168 410542
rect 493048 410462 493168 410478
rect 493048 410398 493076 410462
rect 493140 410398 493168 410462
rect 493048 410382 493168 410398
rect 493048 410318 493076 410382
rect 493140 410318 493168 410382
rect 493048 410302 493168 410318
rect 493048 410238 493076 410302
rect 493140 410238 493168 410302
rect 493048 410222 493168 410238
rect 493048 410158 493076 410222
rect 493140 410158 493168 410222
rect 493048 410142 493168 410158
rect 493048 410078 493076 410142
rect 493140 410078 493168 410142
rect 493048 410062 493168 410078
rect 493048 409998 493076 410062
rect 493140 409998 493168 410062
rect 493048 409974 493168 409998
rect 496808 411582 496928 411606
rect 496808 411518 496836 411582
rect 496900 411518 496928 411582
rect 496808 411502 496928 411518
rect 496808 411438 496836 411502
rect 496900 411438 496928 411502
rect 496808 411422 496928 411438
rect 496808 411358 496836 411422
rect 496900 411358 496928 411422
rect 496808 411342 496928 411358
rect 496808 411278 496836 411342
rect 496900 411278 496928 411342
rect 496808 411262 496928 411278
rect 496808 411198 496836 411262
rect 496900 411198 496928 411262
rect 496808 411182 496928 411198
rect 496808 411118 496836 411182
rect 496900 411118 496928 411182
rect 496808 411102 496928 411118
rect 496808 411038 496836 411102
rect 496900 411038 496928 411102
rect 496808 411022 496928 411038
rect 496808 410958 496836 411022
rect 496900 410958 496928 411022
rect 496808 410942 496928 410958
rect 496808 410878 496836 410942
rect 496900 410878 496928 410942
rect 496808 410862 496928 410878
rect 496808 410798 496836 410862
rect 496900 410798 496928 410862
rect 496808 410782 496928 410798
rect 496808 410718 496836 410782
rect 496900 410718 496928 410782
rect 496808 410702 496928 410718
rect 496808 410638 496836 410702
rect 496900 410638 496928 410702
rect 496808 410622 496928 410638
rect 496808 410558 496836 410622
rect 496900 410558 496928 410622
rect 496808 410542 496928 410558
rect 496808 410478 496836 410542
rect 496900 410478 496928 410542
rect 496808 410462 496928 410478
rect 496808 410398 496836 410462
rect 496900 410398 496928 410462
rect 496808 410382 496928 410398
rect 496808 410318 496836 410382
rect 496900 410318 496928 410382
rect 496808 410302 496928 410318
rect 496808 410238 496836 410302
rect 496900 410238 496928 410302
rect 496808 410222 496928 410238
rect 496808 410158 496836 410222
rect 496900 410158 496928 410222
rect 496808 410142 496928 410158
rect 496808 410078 496836 410142
rect 496900 410078 496928 410142
rect 496808 410062 496928 410078
rect 496808 409998 496836 410062
rect 496900 409998 496928 410062
rect 496808 409974 496928 409998
rect 500568 411582 500688 411606
rect 500568 411518 500596 411582
rect 500660 411518 500688 411582
rect 500568 411502 500688 411518
rect 500568 411438 500596 411502
rect 500660 411438 500688 411502
rect 500568 411422 500688 411438
rect 500568 411358 500596 411422
rect 500660 411358 500688 411422
rect 500568 411342 500688 411358
rect 500568 411278 500596 411342
rect 500660 411278 500688 411342
rect 500568 411262 500688 411278
rect 500568 411198 500596 411262
rect 500660 411198 500688 411262
rect 500568 411182 500688 411198
rect 500568 411118 500596 411182
rect 500660 411118 500688 411182
rect 500568 411102 500688 411118
rect 500568 411038 500596 411102
rect 500660 411038 500688 411102
rect 500568 411022 500688 411038
rect 500568 410958 500596 411022
rect 500660 410958 500688 411022
rect 500568 410942 500688 410958
rect 500568 410878 500596 410942
rect 500660 410878 500688 410942
rect 500568 410862 500688 410878
rect 500568 410798 500596 410862
rect 500660 410798 500688 410862
rect 500568 410782 500688 410798
rect 500568 410718 500596 410782
rect 500660 410718 500688 410782
rect 500568 410702 500688 410718
rect 500568 410638 500596 410702
rect 500660 410638 500688 410702
rect 500568 410622 500688 410638
rect 500568 410558 500596 410622
rect 500660 410558 500688 410622
rect 500568 410542 500688 410558
rect 500568 410478 500596 410542
rect 500660 410478 500688 410542
rect 500568 410462 500688 410478
rect 500568 410398 500596 410462
rect 500660 410398 500688 410462
rect 500568 410382 500688 410398
rect 500568 410318 500596 410382
rect 500660 410318 500688 410382
rect 500568 410302 500688 410318
rect 500568 410238 500596 410302
rect 500660 410238 500688 410302
rect 500568 410222 500688 410238
rect 500568 410158 500596 410222
rect 500660 410158 500688 410222
rect 500568 410142 500688 410158
rect 500568 410078 500596 410142
rect 500660 410078 500688 410142
rect 500568 410062 500688 410078
rect 500568 409998 500596 410062
rect 500660 409998 500688 410062
rect 500568 409974 500688 409998
rect 501026 409786 501086 414806
rect 502448 414030 502568 414054
rect 502448 413966 502476 414030
rect 502540 413966 502568 414030
rect 502448 413950 502568 413966
rect 502448 413886 502476 413950
rect 502540 413886 502568 413950
rect 502448 413870 502568 413886
rect 502448 413806 502476 413870
rect 502540 413806 502568 413870
rect 502448 413790 502568 413806
rect 502448 413726 502476 413790
rect 502540 413726 502568 413790
rect 502448 413710 502568 413726
rect 502448 413646 502476 413710
rect 502540 413646 502568 413710
rect 502448 413630 502568 413646
rect 502448 413566 502476 413630
rect 502540 413566 502568 413630
rect 502448 413550 502568 413566
rect 502448 413486 502476 413550
rect 502540 413486 502568 413550
rect 502448 413470 502568 413486
rect 502448 413406 502476 413470
rect 502540 413406 502568 413470
rect 502448 413390 502568 413406
rect 502448 413326 502476 413390
rect 502540 413326 502568 413390
rect 502448 413310 502568 413326
rect 502448 413246 502476 413310
rect 502540 413246 502568 413310
rect 502448 413230 502568 413246
rect 502448 413166 502476 413230
rect 502540 413166 502568 413230
rect 502448 413150 502568 413166
rect 502448 413086 502476 413150
rect 502540 413086 502568 413150
rect 502448 413070 502568 413086
rect 502448 413006 502476 413070
rect 502540 413006 502568 413070
rect 502448 412990 502568 413006
rect 502448 412926 502476 412990
rect 502540 412926 502568 412990
rect 502448 412910 502568 412926
rect 502448 412846 502476 412910
rect 502540 412846 502568 412910
rect 502448 412830 502568 412846
rect 502448 412766 502476 412830
rect 502540 412766 502568 412830
rect 502448 412750 502568 412766
rect 502448 412686 502476 412750
rect 502540 412686 502568 412750
rect 502448 412670 502568 412686
rect 502448 412606 502476 412670
rect 502540 412606 502568 412670
rect 502448 412590 502568 412606
rect 502448 412526 502476 412590
rect 502540 412526 502568 412590
rect 502448 412510 502568 412526
rect 502448 412446 502476 412510
rect 502540 412446 502568 412510
rect 502448 412422 502568 412446
rect 506208 414030 506328 414054
rect 506208 413966 506236 414030
rect 506300 413966 506328 414030
rect 506208 413950 506328 413966
rect 506208 413886 506236 413950
rect 506300 413886 506328 413950
rect 506208 413870 506328 413886
rect 506208 413806 506236 413870
rect 506300 413806 506328 413870
rect 506208 413790 506328 413806
rect 506208 413726 506236 413790
rect 506300 413726 506328 413790
rect 506208 413710 506328 413726
rect 506208 413646 506236 413710
rect 506300 413646 506328 413710
rect 506208 413630 506328 413646
rect 506208 413566 506236 413630
rect 506300 413566 506328 413630
rect 506208 413550 506328 413566
rect 506208 413486 506236 413550
rect 506300 413486 506328 413550
rect 506208 413470 506328 413486
rect 506208 413406 506236 413470
rect 506300 413406 506328 413470
rect 506208 413390 506328 413406
rect 506208 413326 506236 413390
rect 506300 413326 506328 413390
rect 506208 413310 506328 413326
rect 506208 413246 506236 413310
rect 506300 413246 506328 413310
rect 506208 413230 506328 413246
rect 506208 413166 506236 413230
rect 506300 413166 506328 413230
rect 506208 413150 506328 413166
rect 506208 413086 506236 413150
rect 506300 413086 506328 413150
rect 506208 413070 506328 413086
rect 506208 413006 506236 413070
rect 506300 413006 506328 413070
rect 506208 412990 506328 413006
rect 506208 412926 506236 412990
rect 506300 412926 506328 412990
rect 506208 412910 506328 412926
rect 506208 412846 506236 412910
rect 506300 412846 506328 412910
rect 506208 412830 506328 412846
rect 506208 412766 506236 412830
rect 506300 412766 506328 412830
rect 506208 412750 506328 412766
rect 506208 412686 506236 412750
rect 506300 412686 506328 412750
rect 506208 412670 506328 412686
rect 506208 412606 506236 412670
rect 506300 412606 506328 412670
rect 506208 412590 506328 412606
rect 506208 412526 506236 412590
rect 506300 412526 506328 412590
rect 506208 412510 506328 412526
rect 506208 412446 506236 412510
rect 506300 412446 506328 412510
rect 506208 412422 506328 412446
rect 509968 414030 510088 414054
rect 509968 413966 509996 414030
rect 510060 413966 510088 414030
rect 509968 413950 510088 413966
rect 509968 413886 509996 413950
rect 510060 413886 510088 413950
rect 509968 413870 510088 413886
rect 509968 413806 509996 413870
rect 510060 413806 510088 413870
rect 509968 413790 510088 413806
rect 509968 413726 509996 413790
rect 510060 413726 510088 413790
rect 509968 413710 510088 413726
rect 509968 413646 509996 413710
rect 510060 413646 510088 413710
rect 509968 413630 510088 413646
rect 509968 413566 509996 413630
rect 510060 413566 510088 413630
rect 509968 413550 510088 413566
rect 509968 413486 509996 413550
rect 510060 413486 510088 413550
rect 509968 413470 510088 413486
rect 509968 413406 509996 413470
rect 510060 413406 510088 413470
rect 509968 413390 510088 413406
rect 509968 413326 509996 413390
rect 510060 413326 510088 413390
rect 509968 413310 510088 413326
rect 509968 413246 509996 413310
rect 510060 413246 510088 413310
rect 509968 413230 510088 413246
rect 509968 413166 509996 413230
rect 510060 413166 510088 413230
rect 509968 413150 510088 413166
rect 509968 413086 509996 413150
rect 510060 413086 510088 413150
rect 509968 413070 510088 413086
rect 509968 413006 509996 413070
rect 510060 413006 510088 413070
rect 509968 412990 510088 413006
rect 509968 412926 509996 412990
rect 510060 412926 510088 412990
rect 509968 412910 510088 412926
rect 509968 412846 509996 412910
rect 510060 412846 510088 412910
rect 509968 412830 510088 412846
rect 509968 412766 509996 412830
rect 510060 412766 510088 412830
rect 509968 412750 510088 412766
rect 509968 412686 509996 412750
rect 510060 412686 510088 412750
rect 509968 412670 510088 412686
rect 509968 412606 509996 412670
rect 510060 412606 510088 412670
rect 509968 412590 510088 412606
rect 509968 412526 509996 412590
rect 510060 412526 510088 412590
rect 509968 412510 510088 412526
rect 509968 412446 509996 412510
rect 510060 412446 510088 412510
rect 509968 412422 510088 412446
rect 513728 414030 513848 414054
rect 513728 413966 513756 414030
rect 513820 413966 513848 414030
rect 513728 413950 513848 413966
rect 513728 413886 513756 413950
rect 513820 413886 513848 413950
rect 513728 413870 513848 413886
rect 513728 413806 513756 413870
rect 513820 413806 513848 413870
rect 513728 413790 513848 413806
rect 513728 413726 513756 413790
rect 513820 413726 513848 413790
rect 513728 413710 513848 413726
rect 513728 413646 513756 413710
rect 513820 413646 513848 413710
rect 513728 413630 513848 413646
rect 513728 413566 513756 413630
rect 513820 413566 513848 413630
rect 513728 413550 513848 413566
rect 513728 413486 513756 413550
rect 513820 413486 513848 413550
rect 513728 413470 513848 413486
rect 513728 413406 513756 413470
rect 513820 413406 513848 413470
rect 513728 413390 513848 413406
rect 513728 413326 513756 413390
rect 513820 413326 513848 413390
rect 513728 413310 513848 413326
rect 513728 413246 513756 413310
rect 513820 413246 513848 413310
rect 513728 413230 513848 413246
rect 513728 413166 513756 413230
rect 513820 413166 513848 413230
rect 513728 413150 513848 413166
rect 513728 413086 513756 413150
rect 513820 413086 513848 413150
rect 513728 413070 513848 413086
rect 513728 413006 513756 413070
rect 513820 413006 513848 413070
rect 513728 412990 513848 413006
rect 513728 412926 513756 412990
rect 513820 412926 513848 412990
rect 513728 412910 513848 412926
rect 513728 412846 513756 412910
rect 513820 412846 513848 412910
rect 513728 412830 513848 412846
rect 513728 412766 513756 412830
rect 513820 412766 513848 412830
rect 513728 412750 513848 412766
rect 513728 412686 513756 412750
rect 513820 412686 513848 412750
rect 513728 412670 513848 412686
rect 513728 412606 513756 412670
rect 513820 412606 513848 412670
rect 513728 412590 513848 412606
rect 513728 412526 513756 412590
rect 513820 412526 513848 412590
rect 513728 412510 513848 412526
rect 513728 412446 513756 412510
rect 513820 412446 513848 412510
rect 513728 412422 513848 412446
rect 517488 414030 517608 414054
rect 517488 413966 517516 414030
rect 517580 413966 517608 414030
rect 517488 413950 517608 413966
rect 517488 413886 517516 413950
rect 517580 413886 517608 413950
rect 517488 413870 517608 413886
rect 517488 413806 517516 413870
rect 517580 413806 517608 413870
rect 517488 413790 517608 413806
rect 517488 413726 517516 413790
rect 517580 413726 517608 413790
rect 517488 413710 517608 413726
rect 517488 413646 517516 413710
rect 517580 413646 517608 413710
rect 517488 413630 517608 413646
rect 517488 413566 517516 413630
rect 517580 413566 517608 413630
rect 517488 413550 517608 413566
rect 517488 413486 517516 413550
rect 517580 413486 517608 413550
rect 517488 413470 517608 413486
rect 517488 413406 517516 413470
rect 517580 413406 517608 413470
rect 517488 413390 517608 413406
rect 517488 413326 517516 413390
rect 517580 413326 517608 413390
rect 517488 413310 517608 413326
rect 517488 413246 517516 413310
rect 517580 413246 517608 413310
rect 517488 413230 517608 413246
rect 517488 413166 517516 413230
rect 517580 413166 517608 413230
rect 517488 413150 517608 413166
rect 517488 413086 517516 413150
rect 517580 413086 517608 413150
rect 517488 413070 517608 413086
rect 517488 413006 517516 413070
rect 517580 413006 517608 413070
rect 517488 412990 517608 413006
rect 517488 412926 517516 412990
rect 517580 412926 517608 412990
rect 517488 412910 517608 412926
rect 517488 412846 517516 412910
rect 517580 412846 517608 412910
rect 517488 412830 517608 412846
rect 517488 412766 517516 412830
rect 517580 412766 517608 412830
rect 517488 412750 517608 412766
rect 517488 412686 517516 412750
rect 517580 412686 517608 412750
rect 517488 412670 517608 412686
rect 517488 412606 517516 412670
rect 517580 412606 517608 412670
rect 517488 412590 517608 412606
rect 517488 412526 517516 412590
rect 517580 412526 517608 412590
rect 517488 412510 517608 412526
rect 517488 412446 517516 412510
rect 517580 412446 517608 412510
rect 517488 412422 517608 412446
rect 521248 414030 521368 414054
rect 521248 413966 521276 414030
rect 521340 413966 521368 414030
rect 521248 413950 521368 413966
rect 521248 413886 521276 413950
rect 521340 413886 521368 413950
rect 521248 413870 521368 413886
rect 521248 413806 521276 413870
rect 521340 413806 521368 413870
rect 521248 413790 521368 413806
rect 521248 413726 521276 413790
rect 521340 413726 521368 413790
rect 521248 413710 521368 413726
rect 521248 413646 521276 413710
rect 521340 413646 521368 413710
rect 521248 413630 521368 413646
rect 521248 413566 521276 413630
rect 521340 413566 521368 413630
rect 521248 413550 521368 413566
rect 521248 413486 521276 413550
rect 521340 413486 521368 413550
rect 521248 413470 521368 413486
rect 521248 413406 521276 413470
rect 521340 413406 521368 413470
rect 521248 413390 521368 413406
rect 521248 413326 521276 413390
rect 521340 413326 521368 413390
rect 521248 413310 521368 413326
rect 521248 413246 521276 413310
rect 521340 413246 521368 413310
rect 521248 413230 521368 413246
rect 521248 413166 521276 413230
rect 521340 413166 521368 413230
rect 521248 413150 521368 413166
rect 521248 413086 521276 413150
rect 521340 413086 521368 413150
rect 521248 413070 521368 413086
rect 521248 413006 521276 413070
rect 521340 413006 521368 413070
rect 521248 412990 521368 413006
rect 521248 412926 521276 412990
rect 521340 412926 521368 412990
rect 521248 412910 521368 412926
rect 521248 412846 521276 412910
rect 521340 412846 521368 412910
rect 521248 412830 521368 412846
rect 521248 412766 521276 412830
rect 521340 412766 521368 412830
rect 521248 412750 521368 412766
rect 521248 412686 521276 412750
rect 521340 412686 521368 412750
rect 521248 412670 521368 412686
rect 521248 412606 521276 412670
rect 521340 412606 521368 412670
rect 521248 412590 521368 412606
rect 521248 412526 521276 412590
rect 521340 412526 521368 412590
rect 521248 412510 521368 412526
rect 521248 412446 521276 412510
rect 521340 412446 521368 412510
rect 521248 412422 521368 412446
rect 525008 414030 525128 414054
rect 525008 413966 525036 414030
rect 525100 413966 525128 414030
rect 525008 413950 525128 413966
rect 525008 413886 525036 413950
rect 525100 413886 525128 413950
rect 525008 413870 525128 413886
rect 525008 413806 525036 413870
rect 525100 413806 525128 413870
rect 525008 413790 525128 413806
rect 525008 413726 525036 413790
rect 525100 413726 525128 413790
rect 525008 413710 525128 413726
rect 525008 413646 525036 413710
rect 525100 413646 525128 413710
rect 525008 413630 525128 413646
rect 525008 413566 525036 413630
rect 525100 413566 525128 413630
rect 525008 413550 525128 413566
rect 525008 413486 525036 413550
rect 525100 413486 525128 413550
rect 525008 413470 525128 413486
rect 525008 413406 525036 413470
rect 525100 413406 525128 413470
rect 525008 413390 525128 413406
rect 525008 413326 525036 413390
rect 525100 413326 525128 413390
rect 525008 413310 525128 413326
rect 525008 413246 525036 413310
rect 525100 413246 525128 413310
rect 525008 413230 525128 413246
rect 525008 413166 525036 413230
rect 525100 413166 525128 413230
rect 525008 413150 525128 413166
rect 525008 413086 525036 413150
rect 525100 413086 525128 413150
rect 525008 413070 525128 413086
rect 525008 413006 525036 413070
rect 525100 413006 525128 413070
rect 525008 412990 525128 413006
rect 525008 412926 525036 412990
rect 525100 412926 525128 412990
rect 525008 412910 525128 412926
rect 525008 412846 525036 412910
rect 525100 412846 525128 412910
rect 525008 412830 525128 412846
rect 525008 412766 525036 412830
rect 525100 412766 525128 412830
rect 525008 412750 525128 412766
rect 525008 412686 525036 412750
rect 525100 412686 525128 412750
rect 525008 412670 525128 412686
rect 525008 412606 525036 412670
rect 525100 412606 525128 412670
rect 525008 412590 525128 412606
rect 525008 412526 525036 412590
rect 525100 412526 525128 412590
rect 525008 412510 525128 412526
rect 525008 412446 525036 412510
rect 525100 412446 525128 412510
rect 525008 412422 525128 412446
rect 528768 414030 528888 414054
rect 528768 413966 528796 414030
rect 528860 413966 528888 414030
rect 528768 413950 528888 413966
rect 528768 413886 528796 413950
rect 528860 413886 528888 413950
rect 528768 413870 528888 413886
rect 528768 413806 528796 413870
rect 528860 413806 528888 413870
rect 528768 413790 528888 413806
rect 528768 413726 528796 413790
rect 528860 413726 528888 413790
rect 528768 413710 528888 413726
rect 528768 413646 528796 413710
rect 528860 413646 528888 413710
rect 528768 413630 528888 413646
rect 528768 413566 528796 413630
rect 528860 413566 528888 413630
rect 528768 413550 528888 413566
rect 528768 413486 528796 413550
rect 528860 413486 528888 413550
rect 528768 413470 528888 413486
rect 528768 413406 528796 413470
rect 528860 413406 528888 413470
rect 528768 413390 528888 413406
rect 528768 413326 528796 413390
rect 528860 413326 528888 413390
rect 528768 413310 528888 413326
rect 528768 413246 528796 413310
rect 528860 413246 528888 413310
rect 528768 413230 528888 413246
rect 528768 413166 528796 413230
rect 528860 413166 528888 413230
rect 528768 413150 528888 413166
rect 528768 413086 528796 413150
rect 528860 413086 528888 413150
rect 528768 413070 528888 413086
rect 528768 413006 528796 413070
rect 528860 413006 528888 413070
rect 528768 412990 528888 413006
rect 528768 412926 528796 412990
rect 528860 412926 528888 412990
rect 528768 412910 528888 412926
rect 528768 412846 528796 412910
rect 528860 412846 528888 412910
rect 528768 412830 528888 412846
rect 528768 412766 528796 412830
rect 528860 412766 528888 412830
rect 528768 412750 528888 412766
rect 528768 412686 528796 412750
rect 528860 412686 528888 412750
rect 528768 412670 528888 412686
rect 528768 412606 528796 412670
rect 528860 412606 528888 412670
rect 528768 412590 528888 412606
rect 528768 412526 528796 412590
rect 528860 412526 528888 412590
rect 528768 412510 528888 412526
rect 528768 412446 528796 412510
rect 528860 412446 528888 412510
rect 528768 412422 528888 412446
rect 532528 414030 532648 414054
rect 532528 413966 532556 414030
rect 532620 413966 532648 414030
rect 532528 413950 532648 413966
rect 532528 413886 532556 413950
rect 532620 413886 532648 413950
rect 532528 413870 532648 413886
rect 532528 413806 532556 413870
rect 532620 413806 532648 413870
rect 532528 413790 532648 413806
rect 532528 413726 532556 413790
rect 532620 413726 532648 413790
rect 532528 413710 532648 413726
rect 532528 413646 532556 413710
rect 532620 413646 532648 413710
rect 532528 413630 532648 413646
rect 532528 413566 532556 413630
rect 532620 413566 532648 413630
rect 532528 413550 532648 413566
rect 532528 413486 532556 413550
rect 532620 413486 532648 413550
rect 532528 413470 532648 413486
rect 532528 413406 532556 413470
rect 532620 413406 532648 413470
rect 532528 413390 532648 413406
rect 532528 413326 532556 413390
rect 532620 413326 532648 413390
rect 532528 413310 532648 413326
rect 532528 413246 532556 413310
rect 532620 413246 532648 413310
rect 532528 413230 532648 413246
rect 532528 413166 532556 413230
rect 532620 413166 532648 413230
rect 532528 413150 532648 413166
rect 532528 413086 532556 413150
rect 532620 413086 532648 413150
rect 532528 413070 532648 413086
rect 532528 413006 532556 413070
rect 532620 413006 532648 413070
rect 532528 412990 532648 413006
rect 532528 412926 532556 412990
rect 532620 412926 532648 412990
rect 532528 412910 532648 412926
rect 532528 412846 532556 412910
rect 532620 412846 532648 412910
rect 532528 412830 532648 412846
rect 532528 412766 532556 412830
rect 532620 412766 532648 412830
rect 532528 412750 532648 412766
rect 532528 412686 532556 412750
rect 532620 412686 532648 412750
rect 532528 412670 532648 412686
rect 532528 412606 532556 412670
rect 532620 412606 532648 412670
rect 532528 412590 532648 412606
rect 532528 412526 532556 412590
rect 532620 412526 532648 412590
rect 532528 412510 532648 412526
rect 532528 412446 532556 412510
rect 532620 412446 532648 412510
rect 532528 412422 532648 412446
rect 536288 414030 536408 414054
rect 536288 413966 536316 414030
rect 536380 413966 536408 414030
rect 536288 413950 536408 413966
rect 536288 413886 536316 413950
rect 536380 413886 536408 413950
rect 536288 413870 536408 413886
rect 536288 413806 536316 413870
rect 536380 413806 536408 413870
rect 536288 413790 536408 413806
rect 536288 413726 536316 413790
rect 536380 413726 536408 413790
rect 536288 413710 536408 413726
rect 536288 413646 536316 413710
rect 536380 413646 536408 413710
rect 536288 413630 536408 413646
rect 536288 413566 536316 413630
rect 536380 413566 536408 413630
rect 536288 413550 536408 413566
rect 536288 413486 536316 413550
rect 536380 413486 536408 413550
rect 536288 413470 536408 413486
rect 536288 413406 536316 413470
rect 536380 413406 536408 413470
rect 536288 413390 536408 413406
rect 536288 413326 536316 413390
rect 536380 413326 536408 413390
rect 536288 413310 536408 413326
rect 536288 413246 536316 413310
rect 536380 413246 536408 413310
rect 536288 413230 536408 413246
rect 536288 413166 536316 413230
rect 536380 413166 536408 413230
rect 536288 413150 536408 413166
rect 536288 413086 536316 413150
rect 536380 413086 536408 413150
rect 536288 413070 536408 413086
rect 536288 413006 536316 413070
rect 536380 413006 536408 413070
rect 536288 412990 536408 413006
rect 536288 412926 536316 412990
rect 536380 412926 536408 412990
rect 536288 412910 536408 412926
rect 536288 412846 536316 412910
rect 536380 412846 536408 412910
rect 536288 412830 536408 412846
rect 536288 412766 536316 412830
rect 536380 412766 536408 412830
rect 536288 412750 536408 412766
rect 536288 412686 536316 412750
rect 536380 412686 536408 412750
rect 536288 412670 536408 412686
rect 536288 412606 536316 412670
rect 536380 412606 536408 412670
rect 536288 412590 536408 412606
rect 536288 412526 536316 412590
rect 536380 412526 536408 412590
rect 536288 412510 536408 412526
rect 536288 412446 536316 412510
rect 536380 412446 536408 412510
rect 536288 412422 536408 412446
rect 504328 411582 504448 411606
rect 504328 411518 504356 411582
rect 504420 411518 504448 411582
rect 504328 411502 504448 411518
rect 504328 411438 504356 411502
rect 504420 411438 504448 411502
rect 504328 411422 504448 411438
rect 504328 411358 504356 411422
rect 504420 411358 504448 411422
rect 504328 411342 504448 411358
rect 504328 411278 504356 411342
rect 504420 411278 504448 411342
rect 504328 411262 504448 411278
rect 504328 411198 504356 411262
rect 504420 411198 504448 411262
rect 504328 411182 504448 411198
rect 504328 411118 504356 411182
rect 504420 411118 504448 411182
rect 504328 411102 504448 411118
rect 504328 411038 504356 411102
rect 504420 411038 504448 411102
rect 504328 411022 504448 411038
rect 504328 410958 504356 411022
rect 504420 410958 504448 411022
rect 504328 410942 504448 410958
rect 504328 410878 504356 410942
rect 504420 410878 504448 410942
rect 504328 410862 504448 410878
rect 504328 410798 504356 410862
rect 504420 410798 504448 410862
rect 504328 410782 504448 410798
rect 504328 410718 504356 410782
rect 504420 410718 504448 410782
rect 504328 410702 504448 410718
rect 504328 410638 504356 410702
rect 504420 410638 504448 410702
rect 504328 410622 504448 410638
rect 504328 410558 504356 410622
rect 504420 410558 504448 410622
rect 504328 410542 504448 410558
rect 504328 410478 504356 410542
rect 504420 410478 504448 410542
rect 504328 410462 504448 410478
rect 504328 410398 504356 410462
rect 504420 410398 504448 410462
rect 504328 410382 504448 410398
rect 504328 410318 504356 410382
rect 504420 410318 504448 410382
rect 504328 410302 504448 410318
rect 504328 410238 504356 410302
rect 504420 410238 504448 410302
rect 504328 410222 504448 410238
rect 504328 410158 504356 410222
rect 504420 410158 504448 410222
rect 504328 410142 504448 410158
rect 504328 410078 504356 410142
rect 504420 410078 504448 410142
rect 504328 410062 504448 410078
rect 504328 409998 504356 410062
rect 504420 409998 504448 410062
rect 504328 409974 504448 409998
rect 508088 411582 508208 411606
rect 508088 411518 508116 411582
rect 508180 411518 508208 411582
rect 508088 411502 508208 411518
rect 508088 411438 508116 411502
rect 508180 411438 508208 411502
rect 508088 411422 508208 411438
rect 508088 411358 508116 411422
rect 508180 411358 508208 411422
rect 508088 411342 508208 411358
rect 508088 411278 508116 411342
rect 508180 411278 508208 411342
rect 508088 411262 508208 411278
rect 508088 411198 508116 411262
rect 508180 411198 508208 411262
rect 508088 411182 508208 411198
rect 508088 411118 508116 411182
rect 508180 411118 508208 411182
rect 508088 411102 508208 411118
rect 508088 411038 508116 411102
rect 508180 411038 508208 411102
rect 508088 411022 508208 411038
rect 508088 410958 508116 411022
rect 508180 410958 508208 411022
rect 508088 410942 508208 410958
rect 508088 410878 508116 410942
rect 508180 410878 508208 410942
rect 508088 410862 508208 410878
rect 508088 410798 508116 410862
rect 508180 410798 508208 410862
rect 508088 410782 508208 410798
rect 508088 410718 508116 410782
rect 508180 410718 508208 410782
rect 508088 410702 508208 410718
rect 508088 410638 508116 410702
rect 508180 410638 508208 410702
rect 508088 410622 508208 410638
rect 508088 410558 508116 410622
rect 508180 410558 508208 410622
rect 508088 410542 508208 410558
rect 508088 410478 508116 410542
rect 508180 410478 508208 410542
rect 508088 410462 508208 410478
rect 508088 410398 508116 410462
rect 508180 410398 508208 410462
rect 508088 410382 508208 410398
rect 508088 410318 508116 410382
rect 508180 410318 508208 410382
rect 508088 410302 508208 410318
rect 508088 410238 508116 410302
rect 508180 410238 508208 410302
rect 508088 410222 508208 410238
rect 508088 410158 508116 410222
rect 508180 410158 508208 410222
rect 508088 410142 508208 410158
rect 508088 410078 508116 410142
rect 508180 410078 508208 410142
rect 508088 410062 508208 410078
rect 508088 409998 508116 410062
rect 508180 409998 508208 410062
rect 508088 409974 508208 409998
rect 511848 411582 511968 411606
rect 511848 411518 511876 411582
rect 511940 411518 511968 411582
rect 511848 411502 511968 411518
rect 511848 411438 511876 411502
rect 511940 411438 511968 411502
rect 511848 411422 511968 411438
rect 511848 411358 511876 411422
rect 511940 411358 511968 411422
rect 511848 411342 511968 411358
rect 511848 411278 511876 411342
rect 511940 411278 511968 411342
rect 511848 411262 511968 411278
rect 511848 411198 511876 411262
rect 511940 411198 511968 411262
rect 511848 411182 511968 411198
rect 511848 411118 511876 411182
rect 511940 411118 511968 411182
rect 511848 411102 511968 411118
rect 511848 411038 511876 411102
rect 511940 411038 511968 411102
rect 511848 411022 511968 411038
rect 511848 410958 511876 411022
rect 511940 410958 511968 411022
rect 511848 410942 511968 410958
rect 511848 410878 511876 410942
rect 511940 410878 511968 410942
rect 511848 410862 511968 410878
rect 511848 410798 511876 410862
rect 511940 410798 511968 410862
rect 511848 410782 511968 410798
rect 511848 410718 511876 410782
rect 511940 410718 511968 410782
rect 511848 410702 511968 410718
rect 511848 410638 511876 410702
rect 511940 410638 511968 410702
rect 511848 410622 511968 410638
rect 511848 410558 511876 410622
rect 511940 410558 511968 410622
rect 511848 410542 511968 410558
rect 511848 410478 511876 410542
rect 511940 410478 511968 410542
rect 511848 410462 511968 410478
rect 511848 410398 511876 410462
rect 511940 410398 511968 410462
rect 511848 410382 511968 410398
rect 511848 410318 511876 410382
rect 511940 410318 511968 410382
rect 511848 410302 511968 410318
rect 511848 410238 511876 410302
rect 511940 410238 511968 410302
rect 511848 410222 511968 410238
rect 511848 410158 511876 410222
rect 511940 410158 511968 410222
rect 511848 410142 511968 410158
rect 511848 410078 511876 410142
rect 511940 410078 511968 410142
rect 511848 410062 511968 410078
rect 511848 409998 511876 410062
rect 511940 409998 511968 410062
rect 511848 409974 511968 409998
rect 515608 411582 515728 411606
rect 515608 411518 515636 411582
rect 515700 411518 515728 411582
rect 515608 411502 515728 411518
rect 515608 411438 515636 411502
rect 515700 411438 515728 411502
rect 515608 411422 515728 411438
rect 515608 411358 515636 411422
rect 515700 411358 515728 411422
rect 515608 411342 515728 411358
rect 515608 411278 515636 411342
rect 515700 411278 515728 411342
rect 515608 411262 515728 411278
rect 515608 411198 515636 411262
rect 515700 411198 515728 411262
rect 515608 411182 515728 411198
rect 515608 411118 515636 411182
rect 515700 411118 515728 411182
rect 515608 411102 515728 411118
rect 515608 411038 515636 411102
rect 515700 411038 515728 411102
rect 515608 411022 515728 411038
rect 515608 410958 515636 411022
rect 515700 410958 515728 411022
rect 515608 410942 515728 410958
rect 515608 410878 515636 410942
rect 515700 410878 515728 410942
rect 515608 410862 515728 410878
rect 515608 410798 515636 410862
rect 515700 410798 515728 410862
rect 515608 410782 515728 410798
rect 515608 410718 515636 410782
rect 515700 410718 515728 410782
rect 515608 410702 515728 410718
rect 515608 410638 515636 410702
rect 515700 410638 515728 410702
rect 515608 410622 515728 410638
rect 515608 410558 515636 410622
rect 515700 410558 515728 410622
rect 515608 410542 515728 410558
rect 515608 410478 515636 410542
rect 515700 410478 515728 410542
rect 515608 410462 515728 410478
rect 515608 410398 515636 410462
rect 515700 410398 515728 410462
rect 515608 410382 515728 410398
rect 515608 410318 515636 410382
rect 515700 410318 515728 410382
rect 515608 410302 515728 410318
rect 515608 410238 515636 410302
rect 515700 410238 515728 410302
rect 515608 410222 515728 410238
rect 515608 410158 515636 410222
rect 515700 410158 515728 410222
rect 515608 410142 515728 410158
rect 515608 410078 515636 410142
rect 515700 410078 515728 410142
rect 515608 410062 515728 410078
rect 515608 409998 515636 410062
rect 515700 409998 515728 410062
rect 515608 409974 515728 409998
rect 519368 411582 519488 411606
rect 519368 411518 519396 411582
rect 519460 411518 519488 411582
rect 519368 411502 519488 411518
rect 519368 411438 519396 411502
rect 519460 411438 519488 411502
rect 519368 411422 519488 411438
rect 519368 411358 519396 411422
rect 519460 411358 519488 411422
rect 519368 411342 519488 411358
rect 519368 411278 519396 411342
rect 519460 411278 519488 411342
rect 519368 411262 519488 411278
rect 519368 411198 519396 411262
rect 519460 411198 519488 411262
rect 519368 411182 519488 411198
rect 519368 411118 519396 411182
rect 519460 411118 519488 411182
rect 519368 411102 519488 411118
rect 519368 411038 519396 411102
rect 519460 411038 519488 411102
rect 519368 411022 519488 411038
rect 519368 410958 519396 411022
rect 519460 410958 519488 411022
rect 519368 410942 519488 410958
rect 519368 410878 519396 410942
rect 519460 410878 519488 410942
rect 519368 410862 519488 410878
rect 519368 410798 519396 410862
rect 519460 410798 519488 410862
rect 519368 410782 519488 410798
rect 519368 410718 519396 410782
rect 519460 410718 519488 410782
rect 519368 410702 519488 410718
rect 519368 410638 519396 410702
rect 519460 410638 519488 410702
rect 519368 410622 519488 410638
rect 519368 410558 519396 410622
rect 519460 410558 519488 410622
rect 519368 410542 519488 410558
rect 519368 410478 519396 410542
rect 519460 410478 519488 410542
rect 519368 410462 519488 410478
rect 519368 410398 519396 410462
rect 519460 410398 519488 410462
rect 519368 410382 519488 410398
rect 519368 410318 519396 410382
rect 519460 410318 519488 410382
rect 519368 410302 519488 410318
rect 519368 410238 519396 410302
rect 519460 410238 519488 410302
rect 519368 410222 519488 410238
rect 519368 410158 519396 410222
rect 519460 410158 519488 410222
rect 519368 410142 519488 410158
rect 519368 410078 519396 410142
rect 519460 410078 519488 410142
rect 519368 410062 519488 410078
rect 519368 409998 519396 410062
rect 519460 409998 519488 410062
rect 519368 409974 519488 409998
rect 523128 411582 523248 411606
rect 523128 411518 523156 411582
rect 523220 411518 523248 411582
rect 523128 411502 523248 411518
rect 523128 411438 523156 411502
rect 523220 411438 523248 411502
rect 523128 411422 523248 411438
rect 523128 411358 523156 411422
rect 523220 411358 523248 411422
rect 523128 411342 523248 411358
rect 523128 411278 523156 411342
rect 523220 411278 523248 411342
rect 523128 411262 523248 411278
rect 523128 411198 523156 411262
rect 523220 411198 523248 411262
rect 523128 411182 523248 411198
rect 523128 411118 523156 411182
rect 523220 411118 523248 411182
rect 523128 411102 523248 411118
rect 523128 411038 523156 411102
rect 523220 411038 523248 411102
rect 523128 411022 523248 411038
rect 523128 410958 523156 411022
rect 523220 410958 523248 411022
rect 523128 410942 523248 410958
rect 523128 410878 523156 410942
rect 523220 410878 523248 410942
rect 523128 410862 523248 410878
rect 523128 410798 523156 410862
rect 523220 410798 523248 410862
rect 523128 410782 523248 410798
rect 523128 410718 523156 410782
rect 523220 410718 523248 410782
rect 523128 410702 523248 410718
rect 523128 410638 523156 410702
rect 523220 410638 523248 410702
rect 523128 410622 523248 410638
rect 523128 410558 523156 410622
rect 523220 410558 523248 410622
rect 523128 410542 523248 410558
rect 523128 410478 523156 410542
rect 523220 410478 523248 410542
rect 523128 410462 523248 410478
rect 523128 410398 523156 410462
rect 523220 410398 523248 410462
rect 523128 410382 523248 410398
rect 523128 410318 523156 410382
rect 523220 410318 523248 410382
rect 523128 410302 523248 410318
rect 523128 410238 523156 410302
rect 523220 410238 523248 410302
rect 523128 410222 523248 410238
rect 523128 410158 523156 410222
rect 523220 410158 523248 410222
rect 523128 410142 523248 410158
rect 523128 410078 523156 410142
rect 523220 410078 523248 410142
rect 523128 410062 523248 410078
rect 523128 409998 523156 410062
rect 523220 409998 523248 410062
rect 523128 409974 523248 409998
rect 526888 411582 527008 411606
rect 526888 411518 526916 411582
rect 526980 411518 527008 411582
rect 526888 411502 527008 411518
rect 526888 411438 526916 411502
rect 526980 411438 527008 411502
rect 526888 411422 527008 411438
rect 526888 411358 526916 411422
rect 526980 411358 527008 411422
rect 526888 411342 527008 411358
rect 526888 411278 526916 411342
rect 526980 411278 527008 411342
rect 526888 411262 527008 411278
rect 526888 411198 526916 411262
rect 526980 411198 527008 411262
rect 526888 411182 527008 411198
rect 526888 411118 526916 411182
rect 526980 411118 527008 411182
rect 526888 411102 527008 411118
rect 526888 411038 526916 411102
rect 526980 411038 527008 411102
rect 526888 411022 527008 411038
rect 526888 410958 526916 411022
rect 526980 410958 527008 411022
rect 526888 410942 527008 410958
rect 526888 410878 526916 410942
rect 526980 410878 527008 410942
rect 526888 410862 527008 410878
rect 526888 410798 526916 410862
rect 526980 410798 527008 410862
rect 526888 410782 527008 410798
rect 526888 410718 526916 410782
rect 526980 410718 527008 410782
rect 526888 410702 527008 410718
rect 526888 410638 526916 410702
rect 526980 410638 527008 410702
rect 526888 410622 527008 410638
rect 526888 410558 526916 410622
rect 526980 410558 527008 410622
rect 526888 410542 527008 410558
rect 526888 410478 526916 410542
rect 526980 410478 527008 410542
rect 526888 410462 527008 410478
rect 526888 410398 526916 410462
rect 526980 410398 527008 410462
rect 526888 410382 527008 410398
rect 526888 410318 526916 410382
rect 526980 410318 527008 410382
rect 526888 410302 527008 410318
rect 526888 410238 526916 410302
rect 526980 410238 527008 410302
rect 526888 410222 527008 410238
rect 526888 410158 526916 410222
rect 526980 410158 527008 410222
rect 526888 410142 527008 410158
rect 526888 410078 526916 410142
rect 526980 410078 527008 410142
rect 526888 410062 527008 410078
rect 526888 409998 526916 410062
rect 526980 409998 527008 410062
rect 526888 409974 527008 409998
rect 530648 411582 530768 411606
rect 530648 411518 530676 411582
rect 530740 411518 530768 411582
rect 530648 411502 530768 411518
rect 530648 411438 530676 411502
rect 530740 411438 530768 411502
rect 530648 411422 530768 411438
rect 530648 411358 530676 411422
rect 530740 411358 530768 411422
rect 530648 411342 530768 411358
rect 530648 411278 530676 411342
rect 530740 411278 530768 411342
rect 530648 411262 530768 411278
rect 530648 411198 530676 411262
rect 530740 411198 530768 411262
rect 530648 411182 530768 411198
rect 530648 411118 530676 411182
rect 530740 411118 530768 411182
rect 530648 411102 530768 411118
rect 530648 411038 530676 411102
rect 530740 411038 530768 411102
rect 530648 411022 530768 411038
rect 530648 410958 530676 411022
rect 530740 410958 530768 411022
rect 530648 410942 530768 410958
rect 530648 410878 530676 410942
rect 530740 410878 530768 410942
rect 530648 410862 530768 410878
rect 530648 410798 530676 410862
rect 530740 410798 530768 410862
rect 530648 410782 530768 410798
rect 530648 410718 530676 410782
rect 530740 410718 530768 410782
rect 530648 410702 530768 410718
rect 530648 410638 530676 410702
rect 530740 410638 530768 410702
rect 530648 410622 530768 410638
rect 530648 410558 530676 410622
rect 530740 410558 530768 410622
rect 530648 410542 530768 410558
rect 530648 410478 530676 410542
rect 530740 410478 530768 410542
rect 530648 410462 530768 410478
rect 530648 410398 530676 410462
rect 530740 410398 530768 410462
rect 530648 410382 530768 410398
rect 530648 410318 530676 410382
rect 530740 410318 530768 410382
rect 530648 410302 530768 410318
rect 530648 410238 530676 410302
rect 530740 410238 530768 410302
rect 530648 410222 530768 410238
rect 530648 410158 530676 410222
rect 530740 410158 530768 410222
rect 530648 410142 530768 410158
rect 530648 410078 530676 410142
rect 530740 410078 530768 410142
rect 530648 410062 530768 410078
rect 530648 409998 530676 410062
rect 530740 409998 530768 410062
rect 530648 409974 530768 409998
rect 534408 411582 534528 411606
rect 534408 411518 534436 411582
rect 534500 411518 534528 411582
rect 534408 411502 534528 411518
rect 534408 411438 534436 411502
rect 534500 411438 534528 411502
rect 534408 411422 534528 411438
rect 534408 411358 534436 411422
rect 534500 411358 534528 411422
rect 534408 411342 534528 411358
rect 534408 411278 534436 411342
rect 534500 411278 534528 411342
rect 534408 411262 534528 411278
rect 534408 411198 534436 411262
rect 534500 411198 534528 411262
rect 534408 411182 534528 411198
rect 534408 411118 534436 411182
rect 534500 411118 534528 411182
rect 534408 411102 534528 411118
rect 534408 411038 534436 411102
rect 534500 411038 534528 411102
rect 534408 411022 534528 411038
rect 534408 410958 534436 411022
rect 534500 410958 534528 411022
rect 534408 410942 534528 410958
rect 534408 410878 534436 410942
rect 534500 410878 534528 410942
rect 534408 410862 534528 410878
rect 534408 410798 534436 410862
rect 534500 410798 534528 410862
rect 534408 410782 534528 410798
rect 534408 410718 534436 410782
rect 534500 410718 534528 410782
rect 534408 410702 534528 410718
rect 534408 410638 534436 410702
rect 534500 410638 534528 410702
rect 534408 410622 534528 410638
rect 534408 410558 534436 410622
rect 534500 410558 534528 410622
rect 534408 410542 534528 410558
rect 534408 410478 534436 410542
rect 534500 410478 534528 410542
rect 534408 410462 534528 410478
rect 534408 410398 534436 410462
rect 534500 410398 534528 410462
rect 534408 410382 534528 410398
rect 534408 410318 534436 410382
rect 534500 410318 534528 410382
rect 534408 410302 534528 410318
rect 534408 410238 534436 410302
rect 534500 410238 534528 410302
rect 534408 410222 534528 410238
rect 534408 410158 534436 410222
rect 534500 410158 534528 410222
rect 534408 410142 534528 410158
rect 534408 410078 534436 410142
rect 534500 410078 534528 410142
rect 534408 410062 534528 410078
rect 534408 409998 534436 410062
rect 534500 409998 534528 410062
rect 534408 409974 534528 409998
rect 500660 409726 501086 409786
rect 493338 409006 494638 409038
rect 493338 408950 493350 409006
rect 493406 408950 494638 409006
rect 493338 408926 494638 408950
rect 493338 408870 493350 408926
rect 493406 408870 494638 408926
rect 493338 408422 494638 408870
rect 494738 409008 494858 409036
rect 494738 408944 494766 409008
rect 494830 408944 494858 409008
rect 494738 408928 494770 408944
rect 494826 408928 494858 408944
rect 494738 408864 494766 408928
rect 494830 408864 494858 408928
rect 494738 408836 494858 408864
rect 497098 409006 498398 409038
rect 497098 408950 497110 409006
rect 497166 408950 498398 409006
rect 497098 408926 498398 408950
rect 497098 408870 497110 408926
rect 497166 408870 498398 408926
rect 493338 408358 493366 408422
rect 493430 408358 493446 408422
rect 493510 408358 493526 408422
rect 493590 408358 493606 408422
rect 493670 408358 493686 408422
rect 493750 408358 493766 408422
rect 493830 408358 493846 408422
rect 493910 408358 494066 408422
rect 494130 408358 494146 408422
rect 494210 408358 494226 408422
rect 494290 408358 494306 408422
rect 494370 408358 494386 408422
rect 494450 408358 494466 408422
rect 494530 408358 494546 408422
rect 494610 408358 494638 408422
rect 493338 407703 494638 408358
rect 493338 407639 493366 407703
rect 493430 407639 493446 407703
rect 493510 407639 493526 407703
rect 493590 407639 493606 407703
rect 493670 407639 493686 407703
rect 493750 407639 493766 407703
rect 493830 407639 493846 407703
rect 493910 407639 494066 407703
rect 494130 407639 494146 407703
rect 494210 407639 494226 407703
rect 494290 407639 494306 407703
rect 494370 407639 494386 407703
rect 494450 407639 494466 407703
rect 494530 407639 494546 407703
rect 494610 407639 494638 407703
rect 493338 406984 494638 407639
rect 493338 406920 493366 406984
rect 493430 406920 493446 406984
rect 493510 406920 493526 406984
rect 493590 406920 493606 406984
rect 493670 406920 493686 406984
rect 493750 406920 493766 406984
rect 493830 406920 493846 406984
rect 493910 406920 494066 406984
rect 494130 406920 494146 406984
rect 494210 406920 494226 406984
rect 494290 406920 494306 406984
rect 494370 406920 494386 406984
rect 494450 406920 494466 406984
rect 494530 406920 494546 406984
rect 494610 406920 494638 406984
rect 493338 406265 494638 406920
rect 493338 406201 493366 406265
rect 493430 406201 493446 406265
rect 493510 406201 493526 406265
rect 493590 406201 493606 406265
rect 493670 406201 493686 406265
rect 493750 406201 493766 406265
rect 493830 406201 493846 406265
rect 493910 406201 494066 406265
rect 494130 406201 494146 406265
rect 494210 406201 494226 406265
rect 494290 406201 494306 406265
rect 494370 406201 494386 406265
rect 494450 406201 494466 406265
rect 494530 406201 494546 406265
rect 494610 406201 494638 406265
rect 493338 405546 494638 406201
rect 493338 405482 493366 405546
rect 493430 405482 493446 405546
rect 493510 405482 493526 405546
rect 493590 405482 493606 405546
rect 493670 405482 493686 405546
rect 493750 405482 493766 405546
rect 493830 405482 493846 405546
rect 493910 405482 494066 405546
rect 494130 405482 494146 405546
rect 494210 405482 494226 405546
rect 494290 405482 494306 405546
rect 494370 405482 494386 405546
rect 494450 405482 494466 405546
rect 494530 405482 494546 405546
rect 494610 405482 494638 405546
rect 493338 404827 494638 405482
rect 493338 404763 493366 404827
rect 493430 404763 493446 404827
rect 493510 404763 493526 404827
rect 493590 404763 493606 404827
rect 493670 404763 493686 404827
rect 493750 404763 493766 404827
rect 493830 404763 493846 404827
rect 493910 404763 494066 404827
rect 494130 404763 494146 404827
rect 494210 404763 494226 404827
rect 494290 404763 494306 404827
rect 494370 404763 494386 404827
rect 494450 404763 494466 404827
rect 494530 404763 494546 404827
rect 494610 404763 494638 404827
rect 493338 404108 494638 404763
rect 493338 404044 493366 404108
rect 493430 404044 493446 404108
rect 493510 404044 493526 404108
rect 493590 404044 493606 404108
rect 493670 404044 493686 404108
rect 493750 404044 493766 404108
rect 493830 404044 493846 404108
rect 493910 404044 494066 404108
rect 494130 404044 494146 404108
rect 494210 404044 494226 404108
rect 494290 404044 494306 404108
rect 494370 404044 494386 404108
rect 494450 404044 494466 404108
rect 494530 404044 494546 404108
rect 494610 404044 494638 404108
rect 493338 403389 494638 404044
rect 493338 403325 493366 403389
rect 493430 403325 493446 403389
rect 493510 403325 493526 403389
rect 493590 403325 493606 403389
rect 493670 403325 493686 403389
rect 493750 403325 493766 403389
rect 493830 403325 493846 403389
rect 493910 403325 494066 403389
rect 494130 403325 494146 403389
rect 494210 403325 494226 403389
rect 494290 403325 494306 403389
rect 494370 403325 494386 403389
rect 494450 403325 494466 403389
rect 494530 403325 494546 403389
rect 494610 403325 494638 403389
rect 493338 402670 494638 403325
rect 493338 402606 493366 402670
rect 493430 402606 493446 402670
rect 493510 402606 493526 402670
rect 493590 402606 493606 402670
rect 493670 402606 493686 402670
rect 493750 402606 493766 402670
rect 493830 402606 493846 402670
rect 493910 402606 494066 402670
rect 494130 402606 494146 402670
rect 494210 402606 494226 402670
rect 494290 402606 494306 402670
rect 494370 402606 494386 402670
rect 494450 402606 494466 402670
rect 494530 402606 494546 402670
rect 494610 402606 494638 402670
rect 493338 401951 494638 402606
rect 493338 401887 493366 401951
rect 493430 401887 493446 401951
rect 493510 401887 493526 401951
rect 493590 401887 493606 401951
rect 493670 401887 493686 401951
rect 493750 401887 493766 401951
rect 493830 401887 493846 401951
rect 493910 401887 494066 401951
rect 494130 401887 494146 401951
rect 494210 401887 494226 401951
rect 494290 401887 494306 401951
rect 494370 401887 494386 401951
rect 494450 401887 494466 401951
rect 494530 401887 494546 401951
rect 494610 401887 494638 401951
rect 493338 401866 494638 401887
rect 497098 408422 498398 408870
rect 498498 409008 498618 409036
rect 498498 408944 498526 409008
rect 498590 408944 498618 409008
rect 498498 408928 498530 408944
rect 498586 408928 498618 408944
rect 498498 408864 498526 408928
rect 498590 408864 498618 408928
rect 498498 408836 498618 408864
rect 497098 408358 497126 408422
rect 497190 408358 497206 408422
rect 497270 408358 497286 408422
rect 497350 408358 497366 408422
rect 497430 408358 497446 408422
rect 497510 408358 497526 408422
rect 497590 408358 497606 408422
rect 497670 408358 497826 408422
rect 497890 408358 497906 408422
rect 497970 408358 497986 408422
rect 498050 408358 498066 408422
rect 498130 408358 498146 408422
rect 498210 408358 498226 408422
rect 498290 408358 498306 408422
rect 498370 408358 498398 408422
rect 497098 407703 498398 408358
rect 500660 408046 500720 409726
rect 500858 408614 502158 408646
rect 500858 408558 500870 408614
rect 500926 408558 502158 408614
rect 500858 408534 502158 408558
rect 500858 408478 500870 408534
rect 500926 408478 502158 408534
rect 500658 408040 500722 408046
rect 500658 407970 500722 407976
rect 500858 408030 502158 408478
rect 502258 408616 502378 408644
rect 502258 408552 502286 408616
rect 502350 408552 502378 408616
rect 502258 408536 502290 408552
rect 502346 408536 502378 408552
rect 502258 408472 502286 408536
rect 502350 408472 502378 408536
rect 502258 408444 502378 408472
rect 497098 407639 497126 407703
rect 497190 407639 497206 407703
rect 497270 407639 497286 407703
rect 497350 407639 497366 407703
rect 497430 407639 497446 407703
rect 497510 407639 497526 407703
rect 497590 407639 497606 407703
rect 497670 407639 497826 407703
rect 497890 407639 497906 407703
rect 497970 407639 497986 407703
rect 498050 407639 498066 407703
rect 498130 407639 498146 407703
rect 498210 407639 498226 407703
rect 498290 407639 498306 407703
rect 498370 407639 498398 407703
rect 497098 406984 498398 407639
rect 497098 406920 497126 406984
rect 497190 406920 497206 406984
rect 497270 406920 497286 406984
rect 497350 406920 497366 406984
rect 497430 406920 497446 406984
rect 497510 406920 497526 406984
rect 497590 406920 497606 406984
rect 497670 406920 497826 406984
rect 497890 406920 497906 406984
rect 497970 406920 497986 406984
rect 498050 406920 498066 406984
rect 498130 406920 498146 406984
rect 498210 406920 498226 406984
rect 498290 406920 498306 406984
rect 498370 406920 498398 406984
rect 497098 406265 498398 406920
rect 500858 407966 500886 408030
rect 500950 407966 500966 408030
rect 501030 407966 501046 408030
rect 501110 407966 501126 408030
rect 501190 407966 501206 408030
rect 501270 407966 501286 408030
rect 501350 407966 501366 408030
rect 501430 407966 501586 408030
rect 501650 407966 501666 408030
rect 501730 407966 501746 408030
rect 501810 407966 501826 408030
rect 501890 407966 501906 408030
rect 501970 407966 501986 408030
rect 502050 407966 502066 408030
rect 502130 407966 502158 408030
rect 500858 407311 502158 407966
rect 500858 407247 500886 407311
rect 500950 407247 500966 407311
rect 501030 407247 501046 407311
rect 501110 407247 501126 407311
rect 501190 407247 501206 407311
rect 501270 407247 501286 407311
rect 501350 407247 501366 407311
rect 501430 407247 501586 407311
rect 501650 407247 501666 407311
rect 501730 407247 501746 407311
rect 501810 407247 501826 407311
rect 501890 407247 501906 407311
rect 501970 407247 501986 407311
rect 502050 407247 502066 407311
rect 502130 407247 502158 407311
rect 498706 406661 498770 406666
rect 498705 406660 498771 406661
rect 498705 406596 498706 406660
rect 498770 406596 498771 406660
rect 498705 406595 498771 406596
rect 498706 406590 498770 406595
rect 500858 406592 502158 407247
rect 498708 406506 498768 406590
rect 500858 406528 500886 406592
rect 500950 406528 500966 406592
rect 501030 406528 501046 406592
rect 501110 406528 501126 406592
rect 501190 406528 501206 406592
rect 501270 406528 501286 406592
rect 501350 406528 501366 406592
rect 501430 406528 501586 406592
rect 501650 406528 501666 406592
rect 501730 406528 501746 406592
rect 501810 406528 501826 406592
rect 501890 406528 501906 406592
rect 501970 406528 501986 406592
rect 502050 406528 502066 406592
rect 502130 406528 502158 406592
rect 497098 406201 497126 406265
rect 497190 406201 497206 406265
rect 497270 406201 497286 406265
rect 497350 406201 497366 406265
rect 497430 406201 497446 406265
rect 497510 406201 497526 406265
rect 497590 406201 497606 406265
rect 497670 406201 497826 406265
rect 497890 406201 497906 406265
rect 497970 406201 497986 406265
rect 498050 406201 498066 406265
rect 498130 406201 498146 406265
rect 498210 406201 498226 406265
rect 498290 406201 498306 406265
rect 498370 406201 498398 406265
rect 497098 405546 498398 406201
rect 497098 405482 497126 405546
rect 497190 405482 497206 405546
rect 497270 405482 497286 405546
rect 497350 405482 497366 405546
rect 497430 405482 497446 405546
rect 497510 405482 497526 405546
rect 497590 405482 497606 405546
rect 497670 405482 497826 405546
rect 497890 405482 497906 405546
rect 497970 405482 497986 405546
rect 498050 405482 498066 405546
rect 498130 405482 498146 405546
rect 498210 405482 498226 405546
rect 498290 405482 498306 405546
rect 498370 405482 498398 405546
rect 497098 404827 498398 405482
rect 497098 404763 497126 404827
rect 497190 404763 497206 404827
rect 497270 404763 497286 404827
rect 497350 404763 497366 404827
rect 497430 404763 497446 404827
rect 497510 404763 497526 404827
rect 497590 404763 497606 404827
rect 497670 404763 497826 404827
rect 497890 404763 497906 404827
rect 497970 404763 497986 404827
rect 498050 404763 498066 404827
rect 498130 404763 498146 404827
rect 498210 404763 498226 404827
rect 498290 404763 498306 404827
rect 498370 404763 498398 404827
rect 497098 404108 498398 404763
rect 497098 404044 497126 404108
rect 497190 404044 497206 404108
rect 497270 404044 497286 404108
rect 497350 404044 497366 404108
rect 497430 404044 497446 404108
rect 497510 404044 497526 404108
rect 497590 404044 497606 404108
rect 497670 404044 497826 404108
rect 497890 404044 497906 404108
rect 497970 404044 497986 404108
rect 498050 404044 498066 404108
rect 498130 404044 498146 404108
rect 498210 404044 498226 404108
rect 498290 404044 498306 404108
rect 498370 404044 498398 404108
rect 497098 403389 498398 404044
rect 497098 403325 497126 403389
rect 497190 403325 497206 403389
rect 497270 403325 497286 403389
rect 497350 403325 497366 403389
rect 497430 403325 497446 403389
rect 497510 403325 497526 403389
rect 497590 403325 497606 403389
rect 497670 403325 497826 403389
rect 497890 403325 497906 403389
rect 497970 403325 497986 403389
rect 498050 403325 498066 403389
rect 498130 403325 498146 403389
rect 498210 403325 498226 403389
rect 498290 403325 498306 403389
rect 498370 403325 498398 403389
rect 497098 402670 498398 403325
rect 497098 402606 497126 402670
rect 497190 402606 497206 402670
rect 497270 402606 497286 402670
rect 497350 402606 497366 402670
rect 497430 402606 497446 402670
rect 497510 402606 497526 402670
rect 497590 402606 497606 402670
rect 497670 402606 497826 402670
rect 497890 402606 497906 402670
rect 497970 402606 497986 402670
rect 498050 402606 498066 402670
rect 498130 402606 498146 402670
rect 498210 402606 498226 402670
rect 498290 402606 498306 402670
rect 498370 402606 498398 402670
rect 497098 401951 498398 402606
rect 497098 401887 497126 401951
rect 497190 401887 497206 401951
rect 497270 401887 497286 401951
rect 497350 401887 497366 401951
rect 497430 401887 497446 401951
rect 497510 401887 497526 401951
rect 497590 401887 497606 401951
rect 497670 401887 497826 401951
rect 497890 401887 497906 401951
rect 497970 401887 497986 401951
rect 498050 401887 498066 401951
rect 498130 401887 498146 401951
rect 498210 401887 498226 401951
rect 498290 401887 498306 401951
rect 498370 401887 498398 401951
rect 497098 401866 498398 401887
rect 500858 405873 502158 406528
rect 500858 405809 500886 405873
rect 500950 405809 500966 405873
rect 501030 405809 501046 405873
rect 501110 405809 501126 405873
rect 501190 405809 501206 405873
rect 501270 405809 501286 405873
rect 501350 405809 501366 405873
rect 501430 405809 501586 405873
rect 501650 405809 501666 405873
rect 501730 405809 501746 405873
rect 501810 405809 501826 405873
rect 501890 405809 501906 405873
rect 501970 405809 501986 405873
rect 502050 405809 502066 405873
rect 502130 405809 502158 405873
rect 500858 405154 502158 405809
rect 566246 405476 566472 405481
rect 566246 405400 566256 405476
rect 500858 405090 500886 405154
rect 500950 405090 500966 405154
rect 501030 405090 501046 405154
rect 501110 405090 501126 405154
rect 501190 405090 501206 405154
rect 501270 405090 501286 405154
rect 501350 405090 501366 405154
rect 501430 405090 501586 405154
rect 501650 405090 501666 405154
rect 501730 405090 501746 405154
rect 501810 405090 501826 405154
rect 501890 405090 501906 405154
rect 501970 405090 501986 405154
rect 502050 405090 502066 405154
rect 502130 405090 502158 405154
rect 500858 404435 502158 405090
rect 500858 404371 500886 404435
rect 500950 404371 500966 404435
rect 501030 404371 501046 404435
rect 501110 404371 501126 404435
rect 501190 404371 501206 404435
rect 501270 404371 501286 404435
rect 501350 404371 501366 404435
rect 501430 404371 501586 404435
rect 501650 404371 501666 404435
rect 501730 404371 501746 404435
rect 501810 404371 501826 404435
rect 501890 404371 501906 404435
rect 501970 404371 501986 404435
rect 502050 404371 502066 404435
rect 502130 404371 502158 404435
rect 500858 403716 502158 404371
rect 500858 403652 500886 403716
rect 500950 403652 500966 403716
rect 501030 403652 501046 403716
rect 501110 403652 501126 403716
rect 501190 403652 501206 403716
rect 501270 403652 501286 403716
rect 501350 403652 501366 403716
rect 501430 403652 501586 403716
rect 501650 403652 501666 403716
rect 501730 403652 501746 403716
rect 501810 403652 501826 403716
rect 501890 403652 501906 403716
rect 501970 403652 501986 403716
rect 502050 403652 502066 403716
rect 502130 403652 502158 403716
rect 500858 402997 502158 403652
rect 500858 402933 500886 402997
rect 500950 402933 500966 402997
rect 501030 402933 501046 402997
rect 501110 402933 501126 402997
rect 501190 402933 501206 402997
rect 501270 402933 501286 402997
rect 501350 402933 501366 402997
rect 501430 402933 501586 402997
rect 501650 402933 501666 402997
rect 501730 402933 501746 402997
rect 501810 402933 501826 402997
rect 501890 402933 501906 402997
rect 501970 402933 501986 402997
rect 502050 402933 502066 402997
rect 502130 402933 502158 402997
rect 500858 402278 502158 402933
rect 500858 402214 500886 402278
rect 500950 402214 500966 402278
rect 501030 402214 501046 402278
rect 501110 402214 501126 402278
rect 501190 402214 501206 402278
rect 501270 402214 501286 402278
rect 501350 402214 501366 402278
rect 501430 402214 501586 402278
rect 501650 402214 501666 402278
rect 501730 402214 501746 402278
rect 501810 402214 501826 402278
rect 501890 402214 501906 402278
rect 501970 402214 501986 402278
rect 502050 402214 502066 402278
rect 502130 402214 502158 402278
rect 493338 401558 494638 401590
rect 493338 401502 493350 401558
rect 493406 401502 494638 401558
rect 493338 401478 494638 401502
rect 493338 401422 493350 401478
rect 493406 401422 494638 401478
rect 493338 400974 494638 401422
rect 494738 401560 494858 401588
rect 494738 401496 494766 401560
rect 494830 401496 494858 401560
rect 494738 401480 494770 401496
rect 494826 401480 494858 401496
rect 498218 401554 498282 401560
rect 498218 401484 498282 401490
rect 500858 401559 502158 402214
rect 542962 405288 566256 405400
rect 504805 402056 504871 402061
rect 504805 402000 504810 402056
rect 504866 402000 504871 402056
rect 504805 401995 504871 402000
rect 500858 401495 500886 401559
rect 500950 401495 500966 401559
rect 501030 401495 501046 401559
rect 501110 401495 501126 401559
rect 501190 401495 501206 401559
rect 501270 401495 501286 401559
rect 501350 401495 501366 401559
rect 501430 401495 501586 401559
rect 501650 401495 501666 401559
rect 501730 401495 501746 401559
rect 501810 401495 501826 401559
rect 501890 401495 501906 401559
rect 501970 401495 501986 401559
rect 502050 401495 502066 401559
rect 502130 401495 502158 401559
rect 494738 401416 494766 401480
rect 494830 401416 494858 401480
rect 494738 401388 494858 401416
rect 493338 400910 493366 400974
rect 493430 400910 493446 400974
rect 493510 400910 493526 400974
rect 493590 400910 493606 400974
rect 493670 400910 493686 400974
rect 493750 400910 493766 400974
rect 493830 400910 493846 400974
rect 493910 400910 494066 400974
rect 494130 400910 494146 400974
rect 494210 400910 494226 400974
rect 494290 400910 494306 400974
rect 494370 400910 494386 400974
rect 494450 400910 494466 400974
rect 494530 400910 494546 400974
rect 494610 400910 494638 400974
rect 493338 400255 494638 400910
rect 493338 400191 493366 400255
rect 493430 400191 493446 400255
rect 493510 400191 493526 400255
rect 493590 400191 493606 400255
rect 493670 400191 493686 400255
rect 493750 400191 493766 400255
rect 493830 400191 493846 400255
rect 493910 400191 494066 400255
rect 494130 400191 494146 400255
rect 494210 400191 494226 400255
rect 494290 400191 494306 400255
rect 494370 400191 494386 400255
rect 494450 400191 494466 400255
rect 494530 400191 494546 400255
rect 494610 400191 494638 400255
rect 493338 399536 494638 400191
rect 498220 399945 498280 401484
rect 500858 401474 502158 401495
rect 504808 401422 504868 401995
rect 504806 401416 504870 401422
rect 504806 401346 504870 401352
rect 498583 400400 498649 400405
rect 498583 400344 498588 400400
rect 498644 400344 498649 400400
rect 498583 400339 498649 400344
rect 498217 399940 498283 399945
rect 498217 399884 498222 399940
rect 498278 399884 498283 399940
rect 498217 399879 498283 399884
rect 493338 399472 493366 399536
rect 493430 399472 493446 399536
rect 493510 399472 493526 399536
rect 493590 399472 493606 399536
rect 493670 399472 493686 399536
rect 493750 399472 493766 399536
rect 493830 399472 493846 399536
rect 493910 399472 494066 399536
rect 494130 399472 494146 399536
rect 494210 399472 494226 399536
rect 494290 399472 494306 399536
rect 494370 399472 494386 399536
rect 494450 399472 494466 399536
rect 494530 399472 494546 399536
rect 494610 399472 494638 399536
rect 493338 398817 494638 399472
rect 493338 398753 493366 398817
rect 493430 398753 493446 398817
rect 493510 398753 493526 398817
rect 493590 398753 493606 398817
rect 493670 398753 493686 398817
rect 493750 398753 493766 398817
rect 493830 398753 493846 398817
rect 493910 398753 494066 398817
rect 494130 398753 494146 398817
rect 494210 398753 494226 398817
rect 494290 398753 494306 398817
rect 494370 398753 494386 398817
rect 494450 398753 494466 398817
rect 494530 398753 494546 398817
rect 494610 398753 494638 398817
rect 493338 398098 494638 398753
rect 493338 398034 493366 398098
rect 493430 398034 493446 398098
rect 493510 398034 493526 398098
rect 493590 398034 493606 398098
rect 493670 398034 493686 398098
rect 493750 398034 493766 398098
rect 493830 398034 493846 398098
rect 493910 398034 494066 398098
rect 494130 398034 494146 398098
rect 494210 398034 494226 398098
rect 494290 398034 494306 398098
rect 494370 398034 494386 398098
rect 494450 398034 494466 398098
rect 494530 398034 494546 398098
rect 494610 398034 494638 398098
rect 493338 397379 494638 398034
rect 493338 397315 493366 397379
rect 493430 397315 493446 397379
rect 493510 397315 493526 397379
rect 493590 397315 493606 397379
rect 493670 397315 493686 397379
rect 493750 397315 493766 397379
rect 493830 397315 493846 397379
rect 493910 397315 494066 397379
rect 494130 397315 494146 397379
rect 494210 397315 494226 397379
rect 494290 397315 494306 397379
rect 494370 397315 494386 397379
rect 494450 397315 494466 397379
rect 494530 397315 494546 397379
rect 494610 397315 494638 397379
rect 493338 396660 494638 397315
rect 494926 397282 494986 397366
rect 494924 397277 494988 397282
rect 494923 397276 494989 397277
rect 494923 397212 494924 397276
rect 494988 397212 494989 397276
rect 494923 397211 494989 397212
rect 494924 397206 494988 397211
rect 493338 396596 493366 396660
rect 493430 396596 493446 396660
rect 493510 396596 493526 396660
rect 493590 396596 493606 396660
rect 493670 396596 493686 396660
rect 493750 396596 493766 396660
rect 493830 396596 493846 396660
rect 493910 396596 494066 396660
rect 494130 396596 494146 396660
rect 494210 396596 494226 396660
rect 494290 396596 494306 396660
rect 494370 396596 494386 396660
rect 494450 396596 494466 396660
rect 494530 396596 494546 396660
rect 494610 396596 494638 396660
rect 493338 395941 494638 396596
rect 493338 395877 493366 395941
rect 493430 395877 493446 395941
rect 493510 395877 493526 395941
rect 493590 395877 493606 395941
rect 493670 395877 493686 395941
rect 493750 395877 493766 395941
rect 493830 395877 493846 395941
rect 493910 395877 494066 395941
rect 494130 395877 494146 395941
rect 494210 395877 494226 395941
rect 494290 395877 494306 395941
rect 494370 395877 494386 395941
rect 494450 395877 494466 395941
rect 494530 395877 494546 395941
rect 494610 395877 494638 395941
rect 493338 395222 494638 395877
rect 493338 395158 493366 395222
rect 493430 395158 493446 395222
rect 493510 395158 493526 395222
rect 493590 395158 493606 395222
rect 493670 395158 493686 395222
rect 493750 395158 493766 395222
rect 493830 395158 493846 395222
rect 493910 395158 494066 395222
rect 494130 395158 494146 395222
rect 494210 395158 494226 395222
rect 494290 395158 494306 395222
rect 494370 395158 494386 395222
rect 494450 395158 494466 395222
rect 494530 395158 494546 395222
rect 494610 395158 494638 395222
rect 493338 394503 494638 395158
rect 493338 394439 493366 394503
rect 493430 394439 493446 394503
rect 493510 394439 493526 394503
rect 493590 394439 493606 394503
rect 493670 394439 493686 394503
rect 493750 394439 493766 394503
rect 493830 394439 493846 394503
rect 493910 394439 494066 394503
rect 494130 394439 494146 394503
rect 494210 394439 494226 394503
rect 494290 394439 494306 394503
rect 494370 394439 494386 394503
rect 494450 394439 494466 394503
rect 494530 394439 494546 394503
rect 494610 394439 494638 394503
rect 493338 394418 494638 394439
rect 498586 391205 498646 400339
rect 500858 399794 502158 399826
rect 500858 399738 500870 399794
rect 500926 399738 502158 399794
rect 500858 399714 502158 399738
rect 500858 399658 500870 399714
rect 500926 399658 502158 399714
rect 500858 399210 502158 399658
rect 502258 399796 502378 399824
rect 502258 399732 502286 399796
rect 502350 399732 502378 399796
rect 502258 399716 502290 399732
rect 502346 399716 502378 399732
rect 502258 399652 502286 399716
rect 502350 399652 502378 399716
rect 502258 399624 502378 399652
rect 502366 399485 502430 399490
rect 502365 399484 502431 399485
rect 502365 399420 502366 399484
rect 502430 399420 502431 399484
rect 502365 399419 502431 399420
rect 502366 399414 502430 399419
rect 502368 399330 502428 399414
rect 500858 399146 500886 399210
rect 500950 399146 500966 399210
rect 501030 399146 501046 399210
rect 501110 399146 501126 399210
rect 501190 399146 501206 399210
rect 501270 399146 501286 399210
rect 501350 399146 501366 399210
rect 501430 399146 501586 399210
rect 501650 399146 501666 399210
rect 501730 399146 501746 399210
rect 501810 399146 501826 399210
rect 501890 399146 501906 399210
rect 501970 399146 501986 399210
rect 502050 399146 502066 399210
rect 502130 399146 502158 399210
rect 500858 398491 502158 399146
rect 500858 398427 500886 398491
rect 500950 398427 500966 398491
rect 501030 398427 501046 398491
rect 501110 398427 501126 398491
rect 501190 398427 501206 398491
rect 501270 398427 501286 398491
rect 501350 398427 501366 398491
rect 501430 398427 501586 398491
rect 501650 398427 501666 398491
rect 501730 398427 501746 398491
rect 501810 398427 501826 398491
rect 501890 398427 501906 398491
rect 501970 398427 501986 398491
rect 502050 398427 502066 398491
rect 502130 398427 502158 398491
rect 500858 397772 502158 398427
rect 500858 397708 500886 397772
rect 500950 397708 500966 397772
rect 501030 397708 501046 397772
rect 501110 397708 501126 397772
rect 501190 397708 501206 397772
rect 501270 397708 501286 397772
rect 501350 397708 501366 397772
rect 501430 397708 501586 397772
rect 501650 397708 501666 397772
rect 501730 397708 501746 397772
rect 501810 397708 501826 397772
rect 501890 397708 501906 397772
rect 501970 397708 501986 397772
rect 502050 397708 502066 397772
rect 502130 397708 502158 397772
rect 500858 397053 502158 397708
rect 500858 396989 500886 397053
rect 500950 396989 500966 397053
rect 501030 396989 501046 397053
rect 501110 396989 501126 397053
rect 501190 396989 501206 397053
rect 501270 396989 501286 397053
rect 501350 396989 501366 397053
rect 501430 396989 501586 397053
rect 501650 396989 501666 397053
rect 501730 396989 501746 397053
rect 501810 396989 501826 397053
rect 501890 396989 501906 397053
rect 501970 396989 501986 397053
rect 502050 396989 502066 397053
rect 502130 396989 502158 397053
rect 500858 396334 502158 396989
rect 500858 396270 500886 396334
rect 500950 396270 500966 396334
rect 501030 396270 501046 396334
rect 501110 396270 501126 396334
rect 501190 396270 501206 396334
rect 501270 396270 501286 396334
rect 501350 396270 501366 396334
rect 501430 396270 501586 396334
rect 501650 396270 501666 396334
rect 501730 396270 501746 396334
rect 501810 396270 501826 396334
rect 501890 396270 501906 396334
rect 501970 396270 501986 396334
rect 502050 396270 502066 396334
rect 502130 396270 502158 396334
rect 500858 395615 502158 396270
rect 500858 395551 500886 395615
rect 500950 395551 500966 395615
rect 501030 395551 501046 395615
rect 501110 395551 501126 395615
rect 501190 395551 501206 395615
rect 501270 395551 501286 395615
rect 501350 395551 501366 395615
rect 501430 395551 501586 395615
rect 501650 395551 501666 395615
rect 501730 395551 501746 395615
rect 501810 395551 501826 395615
rect 501890 395551 501906 395615
rect 501970 395551 501986 395615
rect 502050 395551 502066 395615
rect 502130 395551 502158 395615
rect 500858 394896 502158 395551
rect 500858 394832 500886 394896
rect 500950 394832 500966 394896
rect 501030 394832 501046 394896
rect 501110 394832 501126 394896
rect 501190 394832 501206 394896
rect 501270 394832 501286 394896
rect 501350 394832 501366 394896
rect 501430 394832 501586 394896
rect 501650 394832 501666 394896
rect 501730 394832 501746 394896
rect 501810 394832 501826 394896
rect 501890 394832 501906 394896
rect 501970 394832 501986 394896
rect 502050 394832 502066 394896
rect 502130 394832 502158 394896
rect 500858 394177 502158 394832
rect 500858 394113 500886 394177
rect 500950 394113 500966 394177
rect 501030 394113 501046 394177
rect 501110 394113 501126 394177
rect 501190 394113 501206 394177
rect 501270 394113 501286 394177
rect 501350 394113 501366 394177
rect 501430 394113 501586 394177
rect 501650 394113 501666 394177
rect 501730 394113 501746 394177
rect 501810 394113 501826 394177
rect 501890 394113 501906 394177
rect 501970 394113 501986 394177
rect 502050 394113 502066 394177
rect 502130 394113 502158 394177
rect 500858 393458 502158 394113
rect 500858 393394 500886 393458
rect 500950 393394 500966 393458
rect 501030 393394 501046 393458
rect 501110 393394 501126 393458
rect 501190 393394 501206 393458
rect 501270 393394 501286 393458
rect 501350 393394 501366 393458
rect 501430 393394 501586 393458
rect 501650 393394 501666 393458
rect 501730 393394 501746 393458
rect 501810 393394 501826 393458
rect 501890 393394 501906 393458
rect 501970 393394 501986 393458
rect 502050 393394 502066 393458
rect 502130 393394 502158 393458
rect 500660 392769 500720 392812
rect 500657 392764 500723 392769
rect 500657 392722 500662 392764
rect 500718 392722 500723 392764
rect 500657 392703 500658 392722
rect 500722 392703 500723 392722
rect 500858 392739 502158 393394
rect 500658 392652 500722 392658
rect 500858 392675 500886 392739
rect 500950 392675 500966 392739
rect 501030 392675 501046 392739
rect 501110 392675 501126 392739
rect 501190 392675 501206 392739
rect 501270 392675 501286 392739
rect 501350 392675 501366 392739
rect 501430 392675 501586 392739
rect 501650 392675 501666 392739
rect 501730 392675 501746 392739
rect 501810 392675 501826 392739
rect 501890 392675 501906 392739
rect 501970 392675 501986 392739
rect 502050 392675 502066 392739
rect 502130 392675 502158 392739
rect 500858 392654 502158 392675
rect 498583 391200 498649 391205
rect 498583 391144 498588 391200
rect 498644 391144 498649 391200
rect 498583 391139 498649 391144
rect 542962 389490 543074 405288
rect 566246 405258 566256 405288
rect 566462 405400 566472 405476
rect 580064 405402 580192 405407
rect 580064 405400 580074 405402
rect 566462 405292 580074 405400
rect 580182 405400 580192 405402
rect 580182 405292 583872 405400
rect 566462 405288 583872 405292
rect 566462 405258 566472 405288
rect 580064 405287 580192 405288
rect 566246 405253 566472 405258
rect 559726 403368 559936 403373
rect 559726 403192 559736 403368
rect 559926 403192 559936 403368
rect 559726 403187 559936 403192
rect 573528 403312 573898 403317
rect 573528 402980 573538 403312
rect 573888 402980 573898 403312
rect 573528 402975 573898 402980
rect 541910 389470 543074 389490
rect 541910 389388 541952 389470
rect 542058 389388 543074 389470
rect 541910 389378 543074 389388
rect 508378 388720 509678 388752
rect 508378 388664 508390 388720
rect 508446 388664 509678 388720
rect 508378 388640 509678 388664
rect 508378 388584 508390 388640
rect 508446 388584 509678 388640
rect 508378 388136 509678 388584
rect 509778 388722 509898 388750
rect 509778 388658 509806 388722
rect 509870 388658 509898 388722
rect 509778 388642 509810 388658
rect 509866 388642 509898 388658
rect 509778 388578 509806 388642
rect 509870 388578 509898 388642
rect 509778 388550 509898 388578
rect 508378 388072 508406 388136
rect 508470 388072 508486 388136
rect 508550 388072 508566 388136
rect 508630 388072 508646 388136
rect 508710 388072 508726 388136
rect 508790 388072 508806 388136
rect 508870 388072 508886 388136
rect 508950 388072 509106 388136
rect 509170 388072 509186 388136
rect 509250 388072 509266 388136
rect 509330 388072 509346 388136
rect 509410 388072 509426 388136
rect 509490 388072 509506 388136
rect 509570 388072 509586 388136
rect 509650 388072 509678 388136
rect 508378 387417 509678 388072
rect 508378 387353 508406 387417
rect 508470 387353 508486 387417
rect 508550 387353 508566 387417
rect 508630 387353 508646 387417
rect 508710 387353 508726 387417
rect 508790 387353 508806 387417
rect 508870 387353 508886 387417
rect 508950 387353 509106 387417
rect 509170 387353 509186 387417
rect 509250 387353 509266 387417
rect 509330 387353 509346 387417
rect 509410 387353 509426 387417
rect 509490 387353 509506 387417
rect 509570 387353 509586 387417
rect 509650 387353 509678 387417
rect 508378 386698 509678 387353
rect 508378 386634 508406 386698
rect 508470 386634 508486 386698
rect 508550 386634 508566 386698
rect 508630 386634 508646 386698
rect 508710 386634 508726 386698
rect 508790 386634 508806 386698
rect 508870 386634 508886 386698
rect 508950 386634 509106 386698
rect 509170 386634 509186 386698
rect 509250 386634 509266 386698
rect 509330 386634 509346 386698
rect 509410 386634 509426 386698
rect 509490 386634 509506 386698
rect 509570 386634 509586 386698
rect 509650 386634 509678 386698
rect 508378 385979 509678 386634
rect 508378 385915 508406 385979
rect 508470 385915 508486 385979
rect 508550 385915 508566 385979
rect 508630 385915 508646 385979
rect 508710 385915 508726 385979
rect 508790 385915 508806 385979
rect 508870 385915 508886 385979
rect 508950 385915 509106 385979
rect 509170 385915 509186 385979
rect 509250 385915 509266 385979
rect 509330 385915 509346 385979
rect 509410 385915 509426 385979
rect 509490 385915 509506 385979
rect 509570 385915 509586 385979
rect 509650 385915 509678 385979
rect 505049 385496 505115 385501
rect 505049 385440 505054 385496
rect 505110 385440 505115 385496
rect 505049 385435 505115 385440
rect 505052 385276 505112 385435
rect 505050 385270 505114 385276
rect 505050 385200 505114 385206
rect 508378 385260 509678 385915
rect 516273 385496 516339 385501
rect 516273 385440 516278 385496
rect 516334 385440 516339 385496
rect 516273 385435 516339 385440
rect 516276 385276 516336 385435
rect 508378 385196 508406 385260
rect 508470 385196 508486 385260
rect 508550 385196 508566 385260
rect 508630 385196 508646 385260
rect 508710 385196 508726 385260
rect 508790 385196 508806 385260
rect 508870 385196 508886 385260
rect 508950 385196 509106 385260
rect 509170 385196 509186 385260
rect 509250 385196 509266 385260
rect 509330 385196 509346 385260
rect 509410 385196 509426 385260
rect 509490 385196 509506 385260
rect 509570 385196 509586 385260
rect 509650 385196 509678 385260
rect 516274 385270 516338 385276
rect 516274 385200 516338 385206
rect 504618 384996 505918 385028
rect 504618 384940 504630 384996
rect 504686 384940 505918 384996
rect 504618 384916 505918 384940
rect 504618 384860 504630 384916
rect 504686 384860 505918 384916
rect 504618 384412 505918 384860
rect 506018 384998 506138 385026
rect 506018 384934 506046 384998
rect 506110 384934 506138 384998
rect 506018 384918 506050 384934
rect 506106 384918 506138 384934
rect 506018 384854 506046 384918
rect 506110 384854 506138 384918
rect 506018 384826 506138 384854
rect 504618 384348 504646 384412
rect 504710 384348 504726 384412
rect 504790 384348 504806 384412
rect 504870 384348 504886 384412
rect 504950 384348 504966 384412
rect 505030 384348 505046 384412
rect 505110 384348 505126 384412
rect 505190 384348 505346 384412
rect 505410 384348 505426 384412
rect 505490 384348 505506 384412
rect 505570 384348 505586 384412
rect 505650 384348 505666 384412
rect 505730 384348 505746 384412
rect 505810 384348 505826 384412
rect 505890 384348 505918 384412
rect 504618 383693 505918 384348
rect 504618 383629 504646 383693
rect 504710 383629 504726 383693
rect 504790 383629 504806 383693
rect 504870 383629 504886 383693
rect 504950 383629 504966 383693
rect 505030 383629 505046 383693
rect 505110 383629 505126 383693
rect 505190 383629 505346 383693
rect 505410 383629 505426 383693
rect 505490 383629 505506 383693
rect 505570 383629 505586 383693
rect 505650 383629 505666 383693
rect 505730 383629 505746 383693
rect 505810 383629 505826 383693
rect 505890 383629 505918 383693
rect 504618 382974 505918 383629
rect 504618 382910 504646 382974
rect 504710 382910 504726 382974
rect 504790 382910 504806 382974
rect 504870 382910 504886 382974
rect 504950 382910 504966 382974
rect 505030 382910 505046 382974
rect 505110 382910 505126 382974
rect 505190 382910 505346 382974
rect 505410 382910 505426 382974
rect 505490 382910 505506 382974
rect 505570 382910 505586 382974
rect 505650 382910 505666 382974
rect 505730 382910 505746 382974
rect 505810 382910 505826 382974
rect 505890 382910 505918 382974
rect 504618 382255 505918 382910
rect 504618 382191 504646 382255
rect 504710 382191 504726 382255
rect 504790 382191 504806 382255
rect 504870 382191 504886 382255
rect 504950 382191 504966 382255
rect 505030 382191 505046 382255
rect 505110 382191 505126 382255
rect 505190 382191 505346 382255
rect 505410 382191 505426 382255
rect 505490 382191 505506 382255
rect 505570 382191 505586 382255
rect 505650 382191 505666 382255
rect 505730 382191 505746 382255
rect 505810 382191 505826 382255
rect 505890 382191 505918 382255
rect 504442 381550 504502 381634
rect 504440 381545 504504 381550
rect 504439 381544 504505 381545
rect 504439 381480 504440 381544
rect 504504 381480 504505 381544
rect 504439 381479 504505 381480
rect 504618 381536 505918 382191
rect 508378 384541 509678 385196
rect 508378 384477 508406 384541
rect 508470 384477 508486 384541
rect 508550 384477 508566 384541
rect 508630 384477 508646 384541
rect 508710 384477 508726 384541
rect 508790 384477 508806 384541
rect 508870 384477 508886 384541
rect 508950 384477 509106 384541
rect 509170 384477 509186 384541
rect 509250 384477 509266 384541
rect 509330 384477 509346 384541
rect 509410 384477 509426 384541
rect 509490 384477 509506 384541
rect 509570 384477 509586 384541
rect 509650 384477 509678 384541
rect 508378 383822 509678 384477
rect 508378 383758 508406 383822
rect 508470 383758 508486 383822
rect 508550 383758 508566 383822
rect 508630 383758 508646 383822
rect 508710 383758 508726 383822
rect 508790 383758 508806 383822
rect 508870 383758 508886 383822
rect 508950 383758 509106 383822
rect 509170 383758 509186 383822
rect 509250 383758 509266 383822
rect 509330 383758 509346 383822
rect 509410 383758 509426 383822
rect 509490 383758 509506 383822
rect 509570 383758 509586 383822
rect 509650 383758 509678 383822
rect 508378 383103 509678 383758
rect 508378 383039 508406 383103
rect 508470 383039 508486 383103
rect 508550 383039 508566 383103
rect 508630 383039 508646 383103
rect 508710 383039 508726 383103
rect 508790 383039 508806 383103
rect 508870 383039 508886 383103
rect 508950 383039 509106 383103
rect 509170 383039 509186 383103
rect 509250 383039 509266 383103
rect 509330 383039 509346 383103
rect 509410 383039 509426 383103
rect 509490 383039 509506 383103
rect 509570 383039 509586 383103
rect 509650 383039 509678 383103
rect 508378 382384 509678 383039
rect 508378 382320 508406 382384
rect 508470 382320 508486 382384
rect 508550 382320 508566 382384
rect 508630 382320 508646 382384
rect 508710 382320 508726 382384
rect 508790 382320 508806 382384
rect 508870 382320 508886 382384
rect 508950 382320 509106 382384
rect 509170 382320 509186 382384
rect 509250 382320 509266 382384
rect 509330 382320 509346 382384
rect 509410 382320 509426 382384
rect 509490 382320 509506 382384
rect 509570 382320 509586 382384
rect 509650 382320 509678 382384
rect 508222 381682 508286 381688
rect 508222 381612 508286 381618
rect 508378 381665 509678 382320
rect 508224 381545 508284 381612
rect 508378 381601 508406 381665
rect 508470 381601 508486 381665
rect 508550 381601 508566 381665
rect 508630 381601 508646 381665
rect 508710 381601 508726 381665
rect 508790 381601 508806 381665
rect 508870 381601 508886 381665
rect 508950 381601 509106 381665
rect 509170 381601 509186 381665
rect 509250 381601 509266 381665
rect 509330 381601 509346 381665
rect 509410 381601 509426 381665
rect 509490 381601 509506 381665
rect 509570 381601 509586 381665
rect 509650 381601 509678 381665
rect 512138 384996 513438 385028
rect 512138 384940 512150 384996
rect 512206 384940 513438 384996
rect 512138 384916 513438 384940
rect 512138 384860 512150 384916
rect 512206 384860 513438 384916
rect 512138 384412 513438 384860
rect 513538 384998 513658 385026
rect 513538 384934 513566 384998
rect 513630 384934 513658 384998
rect 513538 384918 513570 384934
rect 513626 384918 513658 384934
rect 513538 384854 513566 384918
rect 513630 384854 513658 384918
rect 513538 384826 513658 384854
rect 515898 384996 517198 385028
rect 515898 384940 515910 384996
rect 515966 384940 517198 384996
rect 515898 384916 517198 384940
rect 515898 384860 515910 384916
rect 515966 384860 517198 384916
rect 512138 384348 512166 384412
rect 512230 384348 512246 384412
rect 512310 384348 512326 384412
rect 512390 384348 512406 384412
rect 512470 384348 512486 384412
rect 512550 384348 512566 384412
rect 512630 384348 512646 384412
rect 512710 384348 512866 384412
rect 512930 384348 512946 384412
rect 513010 384348 513026 384412
rect 513090 384348 513106 384412
rect 513170 384348 513186 384412
rect 513250 384348 513266 384412
rect 513330 384348 513346 384412
rect 513410 384348 513438 384412
rect 512138 383693 513438 384348
rect 512138 383629 512166 383693
rect 512230 383629 512246 383693
rect 512310 383629 512326 383693
rect 512390 383629 512406 383693
rect 512470 383629 512486 383693
rect 512550 383629 512566 383693
rect 512630 383629 512646 383693
rect 512710 383629 512866 383693
rect 512930 383629 512946 383693
rect 513010 383629 513026 383693
rect 513090 383629 513106 383693
rect 513170 383629 513186 383693
rect 513250 383629 513266 383693
rect 513330 383629 513346 383693
rect 513410 383629 513438 383693
rect 512138 382974 513438 383629
rect 512138 382910 512166 382974
rect 512230 382910 512246 382974
rect 512310 382910 512326 382974
rect 512390 382910 512406 382974
rect 512470 382910 512486 382974
rect 512550 382910 512566 382974
rect 512630 382910 512646 382974
rect 512710 382910 512866 382974
rect 512930 382910 512946 382974
rect 513010 382910 513026 382974
rect 513090 382910 513106 382974
rect 513170 382910 513186 382974
rect 513250 382910 513266 382974
rect 513330 382910 513346 382974
rect 513410 382910 513438 382974
rect 512138 382255 513438 382910
rect 512138 382191 512166 382255
rect 512230 382191 512246 382255
rect 512310 382191 512326 382255
rect 512390 382191 512406 382255
rect 512470 382191 512486 382255
rect 512550 382191 512566 382255
rect 512630 382191 512646 382255
rect 512710 382191 512866 382255
rect 512930 382191 512946 382255
rect 513010 382191 513026 382255
rect 513090 382191 513106 382255
rect 513170 382191 513186 382255
rect 513250 382191 513266 382255
rect 513330 382191 513346 382255
rect 513410 382191 513438 382255
rect 508378 381580 509678 381601
rect 511884 381550 511944 381634
rect 511882 381545 511946 381550
rect 504440 381474 504504 381479
rect 504618 381472 504646 381536
rect 504710 381472 504726 381536
rect 504790 381472 504806 381536
rect 504870 381472 504886 381536
rect 504950 381472 504966 381536
rect 505030 381472 505046 381536
rect 505110 381472 505126 381536
rect 505190 381472 505346 381536
rect 505410 381472 505426 381536
rect 505490 381472 505506 381536
rect 505570 381472 505586 381536
rect 505650 381472 505666 381536
rect 505730 381472 505746 381536
rect 505810 381472 505826 381536
rect 505890 381472 505918 381536
rect 508221 381540 508287 381545
rect 508221 381484 508226 381540
rect 508282 381484 508287 381540
rect 508221 381479 508287 381484
rect 511881 381544 511947 381545
rect 511881 381480 511882 381544
rect 511946 381480 511947 381544
rect 511881 381479 511947 381480
rect 512138 381536 513438 382191
rect 515898 384412 517198 384860
rect 517298 384998 517418 385026
rect 517298 384934 517326 384998
rect 517390 384934 517418 384998
rect 517298 384918 517330 384934
rect 517386 384918 517418 384934
rect 517298 384854 517326 384918
rect 517390 384854 517418 384918
rect 517298 384826 517418 384854
rect 515898 384348 515926 384412
rect 515990 384348 516006 384412
rect 516070 384348 516086 384412
rect 516150 384348 516166 384412
rect 516230 384348 516246 384412
rect 516310 384348 516326 384412
rect 516390 384348 516406 384412
rect 516470 384348 516626 384412
rect 516690 384348 516706 384412
rect 516770 384348 516786 384412
rect 516850 384348 516866 384412
rect 516930 384348 516946 384412
rect 517010 384348 517026 384412
rect 517090 384348 517106 384412
rect 517170 384348 517198 384412
rect 515898 383693 517198 384348
rect 515898 383629 515926 383693
rect 515990 383629 516006 383693
rect 516070 383629 516086 383693
rect 516150 383629 516166 383693
rect 516230 383629 516246 383693
rect 516310 383629 516326 383693
rect 516390 383629 516406 383693
rect 516470 383629 516626 383693
rect 516690 383629 516706 383693
rect 516770 383629 516786 383693
rect 516850 383629 516866 383693
rect 516930 383629 516946 383693
rect 517010 383629 517026 383693
rect 517090 383629 517106 383693
rect 517170 383629 517198 383693
rect 515898 382974 517198 383629
rect 515898 382910 515926 382974
rect 515990 382910 516006 382974
rect 516070 382910 516086 382974
rect 516150 382910 516166 382974
rect 516230 382910 516246 382974
rect 516310 382910 516326 382974
rect 516390 382910 516406 382974
rect 516470 382910 516626 382974
rect 516690 382910 516706 382974
rect 516770 382910 516786 382974
rect 516850 382910 516866 382974
rect 516930 382910 516946 382974
rect 517010 382910 517026 382974
rect 517090 382910 517106 382974
rect 517170 382910 517198 382974
rect 515898 382255 517198 382910
rect 515898 382191 515926 382255
rect 515990 382191 516006 382255
rect 516070 382191 516086 382255
rect 516150 382191 516166 382255
rect 516230 382191 516246 382255
rect 516310 382191 516326 382255
rect 516390 382191 516406 382255
rect 516470 382191 516626 382255
rect 516690 382191 516706 382255
rect 516770 382191 516786 382255
rect 516850 382191 516866 382255
rect 516930 382191 516946 382255
rect 517010 382191 517026 382255
rect 517090 382191 517106 382255
rect 517170 382191 517198 382255
rect 515666 381550 515726 381634
rect 515664 381545 515728 381550
rect 504618 380817 505918 381472
rect 508224 380860 508284 381479
rect 511882 381474 511946 381479
rect 512138 381472 512166 381536
rect 512230 381472 512246 381536
rect 512310 381472 512326 381536
rect 512390 381472 512406 381536
rect 512470 381472 512486 381536
rect 512550 381472 512566 381536
rect 512630 381472 512646 381536
rect 512710 381472 512866 381536
rect 512930 381472 512946 381536
rect 513010 381472 513026 381536
rect 513090 381472 513106 381536
rect 513170 381472 513186 381536
rect 513250 381472 513266 381536
rect 513330 381472 513346 381536
rect 513410 381472 513438 381536
rect 515663 381544 515729 381545
rect 515663 381480 515664 381544
rect 515728 381480 515729 381544
rect 515663 381479 515729 381480
rect 515898 381536 517198 382191
rect 515664 381474 515728 381479
rect 508378 381272 509678 381304
rect 508378 381216 508390 381272
rect 508446 381216 509678 381272
rect 508378 381192 509678 381216
rect 508378 381136 508390 381192
rect 508446 381136 509678 381192
rect 504618 380753 504646 380817
rect 504710 380753 504726 380817
rect 504790 380753 504806 380817
rect 504870 380753 504886 380817
rect 504950 380753 504966 380817
rect 505030 380753 505046 380817
rect 505110 380753 505126 380817
rect 505190 380753 505346 380817
rect 505410 380753 505426 380817
rect 505490 380753 505506 380817
rect 505570 380753 505586 380817
rect 505650 380753 505666 380817
rect 505730 380753 505746 380817
rect 505810 380753 505826 380817
rect 505890 380753 505918 380817
rect 508222 380854 508286 380860
rect 508222 380784 508286 380790
rect 504618 380098 505918 380753
rect 504618 380034 504646 380098
rect 504710 380034 504726 380098
rect 504790 380034 504806 380098
rect 504870 380034 504886 380098
rect 504950 380034 504966 380098
rect 505030 380034 505046 380098
rect 505110 380034 505126 380098
rect 505190 380034 505346 380098
rect 505410 380034 505426 380098
rect 505490 380034 505506 380098
rect 505570 380034 505586 380098
rect 505650 380034 505666 380098
rect 505730 380034 505746 380098
rect 505810 380034 505826 380098
rect 505890 380034 505918 380098
rect 504618 379379 505918 380034
rect 504618 379315 504646 379379
rect 504710 379315 504726 379379
rect 504790 379315 504806 379379
rect 504870 379315 504886 379379
rect 504950 379315 504966 379379
rect 505030 379315 505046 379379
rect 505110 379315 505126 379379
rect 505190 379315 505346 379379
rect 505410 379315 505426 379379
rect 505490 379315 505506 379379
rect 505570 379315 505586 379379
rect 505650 379315 505666 379379
rect 505730 379315 505746 379379
rect 505810 379315 505826 379379
rect 505890 379315 505918 379379
rect 504618 378660 505918 379315
rect 504618 378596 504646 378660
rect 504710 378596 504726 378660
rect 504790 378596 504806 378660
rect 504870 378596 504886 378660
rect 504950 378596 504966 378660
rect 505030 378596 505046 378660
rect 505110 378596 505126 378660
rect 505190 378596 505346 378660
rect 505410 378596 505426 378660
rect 505490 378596 505506 378660
rect 505570 378596 505586 378660
rect 505650 378596 505666 378660
rect 505730 378596 505746 378660
rect 505810 378596 505826 378660
rect 505890 378596 505918 378660
rect 504618 377941 505918 378596
rect 504618 377877 504646 377941
rect 504710 377877 504726 377941
rect 504790 377877 504806 377941
rect 504870 377877 504886 377941
rect 504950 377877 504966 377941
rect 505030 377877 505046 377941
rect 505110 377877 505126 377941
rect 505190 377877 505346 377941
rect 505410 377877 505426 377941
rect 505490 377877 505506 377941
rect 505570 377877 505586 377941
rect 505650 377877 505666 377941
rect 505730 377877 505746 377941
rect 505810 377877 505826 377941
rect 505890 377877 505918 377941
rect 504618 377856 505918 377877
rect 508378 380688 509678 381136
rect 509778 381274 509898 381302
rect 509778 381210 509806 381274
rect 509870 381210 509898 381274
rect 509778 381194 509810 381210
rect 509866 381194 509898 381210
rect 509778 381130 509806 381194
rect 509870 381130 509898 381194
rect 509778 381102 509898 381130
rect 508378 380624 508406 380688
rect 508470 380624 508486 380688
rect 508550 380624 508566 380688
rect 508630 380624 508646 380688
rect 508710 380624 508726 380688
rect 508790 380624 508806 380688
rect 508870 380624 508886 380688
rect 508950 380624 509106 380688
rect 509170 380624 509186 380688
rect 509250 380624 509266 380688
rect 509330 380624 509346 380688
rect 509410 380624 509426 380688
rect 509490 380624 509506 380688
rect 509570 380624 509586 380688
rect 509650 380624 509678 380688
rect 508378 379969 509678 380624
rect 508378 379905 508406 379969
rect 508470 379905 508486 379969
rect 508550 379905 508566 379969
rect 508630 379905 508646 379969
rect 508710 379905 508726 379969
rect 508790 379905 508806 379969
rect 508870 379905 508886 379969
rect 508950 379905 509106 379969
rect 509170 379905 509186 379969
rect 509250 379905 509266 379969
rect 509330 379905 509346 379969
rect 509410 379905 509426 379969
rect 509490 379905 509506 379969
rect 509570 379905 509586 379969
rect 509650 379905 509678 379969
rect 508378 379250 509678 379905
rect 508378 379186 508406 379250
rect 508470 379186 508486 379250
rect 508550 379186 508566 379250
rect 508630 379186 508646 379250
rect 508710 379186 508726 379250
rect 508790 379186 508806 379250
rect 508870 379186 508886 379250
rect 508950 379186 509106 379250
rect 509170 379186 509186 379250
rect 509250 379186 509266 379250
rect 509330 379186 509346 379250
rect 509410 379186 509426 379250
rect 509490 379186 509506 379250
rect 509570 379186 509586 379250
rect 509650 379186 509678 379250
rect 508378 378531 509678 379186
rect 508378 378467 508406 378531
rect 508470 378467 508486 378531
rect 508550 378467 508566 378531
rect 508630 378467 508646 378531
rect 508710 378467 508726 378531
rect 508790 378467 508806 378531
rect 508870 378467 508886 378531
rect 508950 378467 509106 378531
rect 509170 378467 509186 378531
rect 509250 378467 509266 378531
rect 509330 378467 509346 378531
rect 509410 378467 509426 378531
rect 509490 378467 509506 378531
rect 509570 378467 509586 378531
rect 509650 378467 509678 378531
rect 508378 377812 509678 378467
rect 512138 380817 513438 381472
rect 512138 380753 512166 380817
rect 512230 380753 512246 380817
rect 512310 380753 512326 380817
rect 512390 380753 512406 380817
rect 512470 380753 512486 380817
rect 512550 380753 512566 380817
rect 512630 380753 512646 380817
rect 512710 380753 512866 380817
rect 512930 380753 512946 380817
rect 513010 380753 513026 380817
rect 513090 380753 513106 380817
rect 513170 380753 513186 380817
rect 513250 380753 513266 380817
rect 513330 380753 513346 380817
rect 513410 380753 513438 380817
rect 512138 380098 513438 380753
rect 512138 380034 512166 380098
rect 512230 380034 512246 380098
rect 512310 380034 512326 380098
rect 512390 380034 512406 380098
rect 512470 380034 512486 380098
rect 512550 380034 512566 380098
rect 512630 380034 512646 380098
rect 512710 380034 512866 380098
rect 512930 380034 512946 380098
rect 513010 380034 513026 380098
rect 513090 380034 513106 380098
rect 513170 380034 513186 380098
rect 513250 380034 513266 380098
rect 513330 380034 513346 380098
rect 513410 380034 513438 380098
rect 512138 379379 513438 380034
rect 512138 379315 512166 379379
rect 512230 379315 512246 379379
rect 512310 379315 512326 379379
rect 512390 379315 512406 379379
rect 512470 379315 512486 379379
rect 512550 379315 512566 379379
rect 512630 379315 512646 379379
rect 512710 379315 512866 379379
rect 512930 379315 512946 379379
rect 513010 379315 513026 379379
rect 513090 379315 513106 379379
rect 513170 379315 513186 379379
rect 513250 379315 513266 379379
rect 513330 379315 513346 379379
rect 513410 379315 513438 379379
rect 512138 378660 513438 379315
rect 512138 378596 512166 378660
rect 512230 378596 512246 378660
rect 512310 378596 512326 378660
rect 512390 378596 512406 378660
rect 512470 378596 512486 378660
rect 512550 378596 512566 378660
rect 512630 378596 512646 378660
rect 512710 378596 512866 378660
rect 512930 378596 512946 378660
rect 513010 378596 513026 378660
rect 513090 378596 513106 378660
rect 513170 378596 513186 378660
rect 513250 378596 513266 378660
rect 513330 378596 513346 378660
rect 513410 378596 513438 378660
rect 512138 377941 513438 378596
rect 512138 377877 512166 377941
rect 512230 377877 512246 377941
rect 512310 377877 512326 377941
rect 512390 377877 512406 377941
rect 512470 377877 512486 377941
rect 512550 377877 512566 377941
rect 512630 377877 512646 377941
rect 512710 377877 512866 377941
rect 512930 377877 512946 377941
rect 513010 377877 513026 377941
rect 513090 377877 513106 377941
rect 513170 377877 513186 377941
rect 513250 377877 513266 377941
rect 513330 377877 513346 377941
rect 513410 377877 513438 377941
rect 512138 377856 513438 377877
rect 515898 381472 515926 381536
rect 515990 381472 516006 381536
rect 516070 381472 516086 381536
rect 516150 381472 516166 381536
rect 516230 381472 516246 381536
rect 516310 381472 516326 381536
rect 516390 381472 516406 381536
rect 516470 381472 516626 381536
rect 516690 381472 516706 381536
rect 516770 381472 516786 381536
rect 516850 381472 516866 381536
rect 516930 381472 516946 381536
rect 517010 381472 517026 381536
rect 517090 381472 517106 381536
rect 517170 381472 517198 381536
rect 515898 380817 517198 381472
rect 515898 380753 515926 380817
rect 515990 380753 516006 380817
rect 516070 380753 516086 380817
rect 516150 380753 516166 380817
rect 516230 380753 516246 380817
rect 516310 380753 516326 380817
rect 516390 380753 516406 380817
rect 516470 380753 516626 380817
rect 516690 380753 516706 380817
rect 516770 380753 516786 380817
rect 516850 380753 516866 380817
rect 516930 380753 516946 380817
rect 517010 380753 517026 380817
rect 517090 380753 517106 380817
rect 517170 380753 517198 380817
rect 515898 380098 517198 380753
rect 541937 380644 545137 380703
rect 541937 380564 541958 380644
rect 542066 380615 545137 380644
rect 542066 380564 545141 380615
rect 541937 380499 545141 380564
rect 541959 380497 545141 380499
rect 515898 380034 515926 380098
rect 515990 380034 516006 380098
rect 516070 380034 516086 380098
rect 516150 380034 516166 380098
rect 516230 380034 516246 380098
rect 516310 380034 516326 380098
rect 516390 380034 516406 380098
rect 516470 380034 516626 380098
rect 516690 380034 516706 380098
rect 516770 380034 516786 380098
rect 516850 380034 516866 380098
rect 516930 380034 516946 380098
rect 517010 380034 517026 380098
rect 517090 380034 517106 380098
rect 517170 380034 517198 380098
rect 515898 379379 517198 380034
rect 515898 379315 515926 379379
rect 515990 379315 516006 379379
rect 516070 379315 516086 379379
rect 516150 379315 516166 379379
rect 516230 379315 516246 379379
rect 516310 379315 516326 379379
rect 516390 379315 516406 379379
rect 516470 379315 516626 379379
rect 516690 379315 516706 379379
rect 516770 379315 516786 379379
rect 516850 379315 516866 379379
rect 516930 379315 516946 379379
rect 517010 379315 517026 379379
rect 517090 379315 517106 379379
rect 517170 379315 517198 379379
rect 515898 378660 517198 379315
rect 515898 378596 515926 378660
rect 515990 378596 516006 378660
rect 516070 378596 516086 378660
rect 516150 378596 516166 378660
rect 516230 378596 516246 378660
rect 516310 378596 516326 378660
rect 516390 378596 516406 378660
rect 516470 378596 516626 378660
rect 516690 378596 516706 378660
rect 516770 378596 516786 378660
rect 516850 378596 516866 378660
rect 516930 378596 516946 378660
rect 517010 378596 517026 378660
rect 517090 378596 517106 378660
rect 517170 378596 517198 378660
rect 515898 377941 517198 378596
rect 515898 377877 515926 377941
rect 515990 377877 516006 377941
rect 516070 377877 516086 377941
rect 516150 377877 516166 377941
rect 516230 377877 516246 377941
rect 516310 377877 516326 377941
rect 516390 377877 516406 377941
rect 516470 377877 516626 377941
rect 516690 377877 516706 377941
rect 516770 377877 516786 377941
rect 516850 377877 516866 377941
rect 516930 377877 516946 377941
rect 517010 377877 517026 377941
rect 517090 377877 517106 377941
rect 517170 377877 517198 377941
rect 515898 377856 517198 377877
rect 508378 377748 508406 377812
rect 508470 377748 508486 377812
rect 508550 377748 508566 377812
rect 508630 377748 508646 377812
rect 508710 377748 508726 377812
rect 508790 377748 508806 377812
rect 508870 377748 508886 377812
rect 508950 377748 509106 377812
rect 509170 377748 509186 377812
rect 509250 377748 509266 377812
rect 509330 377748 509346 377812
rect 509410 377748 509426 377812
rect 509490 377748 509506 377812
rect 509570 377748 509586 377812
rect 509650 377748 509678 377812
rect 506028 377410 506088 377494
rect 506026 377405 506090 377410
rect 506025 377404 506091 377405
rect 506025 377340 506026 377404
rect 506090 377340 506091 377404
rect 506025 377339 506091 377340
rect 506026 377334 506090 377339
rect 508378 377093 509678 377748
rect 508378 377029 508406 377093
rect 508470 377029 508486 377093
rect 508550 377029 508566 377093
rect 508630 377029 508646 377093
rect 508710 377029 508726 377093
rect 508790 377029 508806 377093
rect 508870 377029 508886 377093
rect 508950 377029 509106 377093
rect 509170 377029 509186 377093
rect 509250 377029 509266 377093
rect 509330 377029 509346 377093
rect 509410 377029 509426 377093
rect 509490 377029 509506 377093
rect 509570 377029 509586 377093
rect 509650 377029 509678 377093
rect 508378 376374 509678 377029
rect 508378 376310 508406 376374
rect 508470 376310 508486 376374
rect 508550 376310 508566 376374
rect 508630 376310 508646 376374
rect 508710 376310 508726 376374
rect 508790 376310 508806 376374
rect 508870 376310 508886 376374
rect 508950 376310 509106 376374
rect 509170 376310 509186 376374
rect 509250 376310 509266 376374
rect 509330 376310 509346 376374
rect 509410 376310 509426 376374
rect 509490 376310 509506 376374
rect 509570 376310 509586 376374
rect 509650 376310 509678 376374
rect 508378 375655 509678 376310
rect 508378 375591 508406 375655
rect 508470 375591 508486 375655
rect 508550 375591 508566 375655
rect 508630 375591 508646 375655
rect 508710 375591 508726 375655
rect 508790 375591 508806 375655
rect 508870 375591 508886 375655
rect 508950 375591 509106 375655
rect 509170 375591 509186 375655
rect 509250 375591 509266 375655
rect 509330 375591 509346 375655
rect 509410 375591 509426 375655
rect 509490 375591 509506 375655
rect 509570 375591 509586 375655
rect 509650 375591 509678 375655
rect 508378 374936 509678 375591
rect 508378 374872 508406 374936
rect 508470 374872 508486 374936
rect 508550 374872 508566 374936
rect 508630 374872 508646 374936
rect 508710 374872 508726 374936
rect 508790 374872 508806 374936
rect 508870 374872 508886 374936
rect 508950 374872 509106 374936
rect 509170 374872 509186 374936
rect 509250 374872 509266 374936
rect 509330 374872 509346 374936
rect 509410 374872 509426 374936
rect 509490 374872 509506 374936
rect 509570 374872 509586 374936
rect 509650 374872 509678 374936
rect 508378 374217 509678 374872
rect 508378 374153 508406 374217
rect 508470 374153 508486 374217
rect 508550 374153 508566 374217
rect 508630 374153 508646 374217
rect 508710 374153 508726 374217
rect 508790 374153 508806 374217
rect 508870 374153 508886 374217
rect 508950 374153 509106 374217
rect 509170 374153 509186 374217
rect 509250 374153 509266 374217
rect 509330 374153 509346 374217
rect 509410 374153 509426 374217
rect 509490 374153 509506 374217
rect 509570 374153 509586 374217
rect 509650 374153 509678 374217
rect 508378 374132 509678 374153
rect 493048 361474 493168 361498
rect 493048 361410 493076 361474
rect 493140 361410 493168 361474
rect 493048 361394 493168 361410
rect 493048 361330 493076 361394
rect 493140 361330 493168 361394
rect 493048 361314 493168 361330
rect 493048 361250 493076 361314
rect 493140 361250 493168 361314
rect 493048 361234 493168 361250
rect 493048 361170 493076 361234
rect 493140 361170 493168 361234
rect 493048 361154 493168 361170
rect 493048 361090 493076 361154
rect 493140 361090 493168 361154
rect 493048 361074 493168 361090
rect 493048 361010 493076 361074
rect 493140 361010 493168 361074
rect 493048 360994 493168 361010
rect 493048 360930 493076 360994
rect 493140 360930 493168 360994
rect 493048 360914 493168 360930
rect 493048 360850 493076 360914
rect 493140 360850 493168 360914
rect 493048 360834 493168 360850
rect 493048 360770 493076 360834
rect 493140 360770 493168 360834
rect 493048 360754 493168 360770
rect 493048 360690 493076 360754
rect 493140 360690 493168 360754
rect 493048 360674 493168 360690
rect 493048 360610 493076 360674
rect 493140 360610 493168 360674
rect 493048 360594 493168 360610
rect 493048 360530 493076 360594
rect 493140 360530 493168 360594
rect 493048 360514 493168 360530
rect 493048 360450 493076 360514
rect 493140 360450 493168 360514
rect 493048 360434 493168 360450
rect 493048 360370 493076 360434
rect 493140 360370 493168 360434
rect 493048 360354 493168 360370
rect 493048 360290 493076 360354
rect 493140 360290 493168 360354
rect 493048 360274 493168 360290
rect 493048 360210 493076 360274
rect 493140 360210 493168 360274
rect 493048 360194 493168 360210
rect 493048 360130 493076 360194
rect 493140 360130 493168 360194
rect 493048 360114 493168 360130
rect 493048 360050 493076 360114
rect 493140 360050 493168 360114
rect 493048 360034 493168 360050
rect 493048 359970 493076 360034
rect 493140 359970 493168 360034
rect 493048 359954 493168 359970
rect 493048 359890 493076 359954
rect 493140 359890 493168 359954
rect 493048 359866 493168 359890
rect 496808 361474 496928 361498
rect 496808 361410 496836 361474
rect 496900 361410 496928 361474
rect 496808 361394 496928 361410
rect 496808 361330 496836 361394
rect 496900 361330 496928 361394
rect 496808 361314 496928 361330
rect 496808 361250 496836 361314
rect 496900 361250 496928 361314
rect 496808 361234 496928 361250
rect 496808 361170 496836 361234
rect 496900 361170 496928 361234
rect 496808 361154 496928 361170
rect 496808 361090 496836 361154
rect 496900 361090 496928 361154
rect 496808 361074 496928 361090
rect 496808 361010 496836 361074
rect 496900 361010 496928 361074
rect 496808 360994 496928 361010
rect 496808 360930 496836 360994
rect 496900 360930 496928 360994
rect 496808 360914 496928 360930
rect 496808 360850 496836 360914
rect 496900 360850 496928 360914
rect 496808 360834 496928 360850
rect 496808 360770 496836 360834
rect 496900 360770 496928 360834
rect 496808 360754 496928 360770
rect 496808 360690 496836 360754
rect 496900 360690 496928 360754
rect 496808 360674 496928 360690
rect 496808 360610 496836 360674
rect 496900 360610 496928 360674
rect 496808 360594 496928 360610
rect 496808 360530 496836 360594
rect 496900 360530 496928 360594
rect 496808 360514 496928 360530
rect 496808 360450 496836 360514
rect 496900 360450 496928 360514
rect 496808 360434 496928 360450
rect 496808 360370 496836 360434
rect 496900 360370 496928 360434
rect 496808 360354 496928 360370
rect 496808 360290 496836 360354
rect 496900 360290 496928 360354
rect 496808 360274 496928 360290
rect 496808 360210 496836 360274
rect 496900 360210 496928 360274
rect 496808 360194 496928 360210
rect 496808 360130 496836 360194
rect 496900 360130 496928 360194
rect 496808 360114 496928 360130
rect 496808 360050 496836 360114
rect 496900 360050 496928 360114
rect 496808 360034 496928 360050
rect 496808 359970 496836 360034
rect 496900 359970 496928 360034
rect 496808 359954 496928 359970
rect 496808 359890 496836 359954
rect 496900 359890 496928 359954
rect 496808 359866 496928 359890
rect 500568 361474 500688 361498
rect 500568 361410 500596 361474
rect 500660 361410 500688 361474
rect 500568 361394 500688 361410
rect 500568 361330 500596 361394
rect 500660 361330 500688 361394
rect 500568 361314 500688 361330
rect 500568 361250 500596 361314
rect 500660 361250 500688 361314
rect 500568 361234 500688 361250
rect 500568 361170 500596 361234
rect 500660 361170 500688 361234
rect 500568 361154 500688 361170
rect 500568 361090 500596 361154
rect 500660 361090 500688 361154
rect 500568 361074 500688 361090
rect 500568 361010 500596 361074
rect 500660 361010 500688 361074
rect 500568 360994 500688 361010
rect 500568 360930 500596 360994
rect 500660 360930 500688 360994
rect 500568 360914 500688 360930
rect 500568 360850 500596 360914
rect 500660 360850 500688 360914
rect 500568 360834 500688 360850
rect 500568 360770 500596 360834
rect 500660 360770 500688 360834
rect 500568 360754 500688 360770
rect 500568 360690 500596 360754
rect 500660 360690 500688 360754
rect 500568 360674 500688 360690
rect 500568 360610 500596 360674
rect 500660 360610 500688 360674
rect 500568 360594 500688 360610
rect 500568 360530 500596 360594
rect 500660 360530 500688 360594
rect 500568 360514 500688 360530
rect 500568 360450 500596 360514
rect 500660 360450 500688 360514
rect 500568 360434 500688 360450
rect 500568 360370 500596 360434
rect 500660 360370 500688 360434
rect 500568 360354 500688 360370
rect 500568 360290 500596 360354
rect 500660 360290 500688 360354
rect 500568 360274 500688 360290
rect 500568 360210 500596 360274
rect 500660 360210 500688 360274
rect 500568 360194 500688 360210
rect 500568 360130 500596 360194
rect 500660 360130 500688 360194
rect 500568 360114 500688 360130
rect 500568 360050 500596 360114
rect 500660 360050 500688 360114
rect 500568 360034 500688 360050
rect 500568 359970 500596 360034
rect 500660 359970 500688 360034
rect 500568 359954 500688 359970
rect 500568 359890 500596 359954
rect 500660 359890 500688 359954
rect 500568 359866 500688 359890
rect 504328 361474 504448 361498
rect 504328 361410 504356 361474
rect 504420 361410 504448 361474
rect 504328 361394 504448 361410
rect 504328 361330 504356 361394
rect 504420 361330 504448 361394
rect 504328 361314 504448 361330
rect 504328 361250 504356 361314
rect 504420 361250 504448 361314
rect 504328 361234 504448 361250
rect 504328 361170 504356 361234
rect 504420 361170 504448 361234
rect 504328 361154 504448 361170
rect 504328 361090 504356 361154
rect 504420 361090 504448 361154
rect 504328 361074 504448 361090
rect 504328 361010 504356 361074
rect 504420 361010 504448 361074
rect 504328 360994 504448 361010
rect 504328 360930 504356 360994
rect 504420 360930 504448 360994
rect 504328 360914 504448 360930
rect 504328 360850 504356 360914
rect 504420 360850 504448 360914
rect 504328 360834 504448 360850
rect 504328 360770 504356 360834
rect 504420 360770 504448 360834
rect 504328 360754 504448 360770
rect 504328 360690 504356 360754
rect 504420 360690 504448 360754
rect 504328 360674 504448 360690
rect 504328 360610 504356 360674
rect 504420 360610 504448 360674
rect 504328 360594 504448 360610
rect 504328 360530 504356 360594
rect 504420 360530 504448 360594
rect 504328 360514 504448 360530
rect 504328 360450 504356 360514
rect 504420 360450 504448 360514
rect 504328 360434 504448 360450
rect 504328 360370 504356 360434
rect 504420 360370 504448 360434
rect 504328 360354 504448 360370
rect 504328 360290 504356 360354
rect 504420 360290 504448 360354
rect 504328 360274 504448 360290
rect 504328 360210 504356 360274
rect 504420 360210 504448 360274
rect 504328 360194 504448 360210
rect 504328 360130 504356 360194
rect 504420 360130 504448 360194
rect 504328 360114 504448 360130
rect 504328 360050 504356 360114
rect 504420 360050 504448 360114
rect 504328 360034 504448 360050
rect 504328 359970 504356 360034
rect 504420 359970 504448 360034
rect 504328 359954 504448 359970
rect 504328 359890 504356 359954
rect 504420 359890 504448 359954
rect 504328 359866 504448 359890
rect 508088 361474 508208 361498
rect 508088 361410 508116 361474
rect 508180 361410 508208 361474
rect 508088 361394 508208 361410
rect 508088 361330 508116 361394
rect 508180 361330 508208 361394
rect 508088 361314 508208 361330
rect 508088 361250 508116 361314
rect 508180 361250 508208 361314
rect 508088 361234 508208 361250
rect 508088 361170 508116 361234
rect 508180 361170 508208 361234
rect 508088 361154 508208 361170
rect 508088 361090 508116 361154
rect 508180 361090 508208 361154
rect 508088 361074 508208 361090
rect 508088 361010 508116 361074
rect 508180 361010 508208 361074
rect 508088 360994 508208 361010
rect 508088 360930 508116 360994
rect 508180 360930 508208 360994
rect 508088 360914 508208 360930
rect 508088 360850 508116 360914
rect 508180 360850 508208 360914
rect 508088 360834 508208 360850
rect 508088 360770 508116 360834
rect 508180 360770 508208 360834
rect 508088 360754 508208 360770
rect 508088 360690 508116 360754
rect 508180 360690 508208 360754
rect 508088 360674 508208 360690
rect 508088 360610 508116 360674
rect 508180 360610 508208 360674
rect 508088 360594 508208 360610
rect 508088 360530 508116 360594
rect 508180 360530 508208 360594
rect 508088 360514 508208 360530
rect 508088 360450 508116 360514
rect 508180 360450 508208 360514
rect 508088 360434 508208 360450
rect 508088 360370 508116 360434
rect 508180 360370 508208 360434
rect 508088 360354 508208 360370
rect 508088 360290 508116 360354
rect 508180 360290 508208 360354
rect 508088 360274 508208 360290
rect 508088 360210 508116 360274
rect 508180 360210 508208 360274
rect 508088 360194 508208 360210
rect 508088 360130 508116 360194
rect 508180 360130 508208 360194
rect 508088 360114 508208 360130
rect 508088 360050 508116 360114
rect 508180 360050 508208 360114
rect 508088 360034 508208 360050
rect 508088 359970 508116 360034
rect 508180 359970 508208 360034
rect 508088 359954 508208 359970
rect 508088 359890 508116 359954
rect 508180 359890 508208 359954
rect 508088 359866 508208 359890
rect 511848 361474 511968 361498
rect 511848 361410 511876 361474
rect 511940 361410 511968 361474
rect 511848 361394 511968 361410
rect 511848 361330 511876 361394
rect 511940 361330 511968 361394
rect 511848 361314 511968 361330
rect 511848 361250 511876 361314
rect 511940 361250 511968 361314
rect 511848 361234 511968 361250
rect 511848 361170 511876 361234
rect 511940 361170 511968 361234
rect 511848 361154 511968 361170
rect 511848 361090 511876 361154
rect 511940 361090 511968 361154
rect 511848 361074 511968 361090
rect 511848 361010 511876 361074
rect 511940 361010 511968 361074
rect 511848 360994 511968 361010
rect 511848 360930 511876 360994
rect 511940 360930 511968 360994
rect 511848 360914 511968 360930
rect 511848 360850 511876 360914
rect 511940 360850 511968 360914
rect 511848 360834 511968 360850
rect 511848 360770 511876 360834
rect 511940 360770 511968 360834
rect 511848 360754 511968 360770
rect 511848 360690 511876 360754
rect 511940 360690 511968 360754
rect 511848 360674 511968 360690
rect 511848 360610 511876 360674
rect 511940 360610 511968 360674
rect 511848 360594 511968 360610
rect 511848 360530 511876 360594
rect 511940 360530 511968 360594
rect 511848 360514 511968 360530
rect 511848 360450 511876 360514
rect 511940 360450 511968 360514
rect 511848 360434 511968 360450
rect 511848 360370 511876 360434
rect 511940 360370 511968 360434
rect 511848 360354 511968 360370
rect 511848 360290 511876 360354
rect 511940 360290 511968 360354
rect 511848 360274 511968 360290
rect 511848 360210 511876 360274
rect 511940 360210 511968 360274
rect 511848 360194 511968 360210
rect 511848 360130 511876 360194
rect 511940 360130 511968 360194
rect 511848 360114 511968 360130
rect 511848 360050 511876 360114
rect 511940 360050 511968 360114
rect 511848 360034 511968 360050
rect 511848 359970 511876 360034
rect 511940 359970 511968 360034
rect 511848 359954 511968 359970
rect 511848 359890 511876 359954
rect 511940 359890 511968 359954
rect 511848 359866 511968 359890
rect 515608 361474 515728 361498
rect 515608 361410 515636 361474
rect 515700 361410 515728 361474
rect 515608 361394 515728 361410
rect 515608 361330 515636 361394
rect 515700 361330 515728 361394
rect 515608 361314 515728 361330
rect 515608 361250 515636 361314
rect 515700 361250 515728 361314
rect 515608 361234 515728 361250
rect 515608 361170 515636 361234
rect 515700 361170 515728 361234
rect 515608 361154 515728 361170
rect 515608 361090 515636 361154
rect 515700 361090 515728 361154
rect 515608 361074 515728 361090
rect 515608 361010 515636 361074
rect 515700 361010 515728 361074
rect 515608 360994 515728 361010
rect 515608 360930 515636 360994
rect 515700 360930 515728 360994
rect 515608 360914 515728 360930
rect 515608 360850 515636 360914
rect 515700 360850 515728 360914
rect 515608 360834 515728 360850
rect 515608 360770 515636 360834
rect 515700 360770 515728 360834
rect 515608 360754 515728 360770
rect 515608 360690 515636 360754
rect 515700 360690 515728 360754
rect 515608 360674 515728 360690
rect 515608 360610 515636 360674
rect 515700 360610 515728 360674
rect 515608 360594 515728 360610
rect 515608 360530 515636 360594
rect 515700 360530 515728 360594
rect 515608 360514 515728 360530
rect 515608 360450 515636 360514
rect 515700 360450 515728 360514
rect 515608 360434 515728 360450
rect 515608 360370 515636 360434
rect 515700 360370 515728 360434
rect 515608 360354 515728 360370
rect 515608 360290 515636 360354
rect 515700 360290 515728 360354
rect 515608 360274 515728 360290
rect 515608 360210 515636 360274
rect 515700 360210 515728 360274
rect 515608 360194 515728 360210
rect 515608 360130 515636 360194
rect 515700 360130 515728 360194
rect 515608 360114 515728 360130
rect 515608 360050 515636 360114
rect 515700 360050 515728 360114
rect 515608 360034 515728 360050
rect 515608 359970 515636 360034
rect 515700 359970 515728 360034
rect 515608 359954 515728 359970
rect 515608 359890 515636 359954
rect 515700 359890 515728 359954
rect 515608 359866 515728 359890
rect 519368 361474 519488 361498
rect 519368 361410 519396 361474
rect 519460 361410 519488 361474
rect 519368 361394 519488 361410
rect 519368 361330 519396 361394
rect 519460 361330 519488 361394
rect 519368 361314 519488 361330
rect 519368 361250 519396 361314
rect 519460 361250 519488 361314
rect 519368 361234 519488 361250
rect 519368 361170 519396 361234
rect 519460 361170 519488 361234
rect 519368 361154 519488 361170
rect 519368 361090 519396 361154
rect 519460 361090 519488 361154
rect 519368 361074 519488 361090
rect 519368 361010 519396 361074
rect 519460 361010 519488 361074
rect 519368 360994 519488 361010
rect 519368 360930 519396 360994
rect 519460 360930 519488 360994
rect 519368 360914 519488 360930
rect 519368 360850 519396 360914
rect 519460 360850 519488 360914
rect 519368 360834 519488 360850
rect 519368 360770 519396 360834
rect 519460 360770 519488 360834
rect 519368 360754 519488 360770
rect 519368 360690 519396 360754
rect 519460 360690 519488 360754
rect 519368 360674 519488 360690
rect 519368 360610 519396 360674
rect 519460 360610 519488 360674
rect 519368 360594 519488 360610
rect 519368 360530 519396 360594
rect 519460 360530 519488 360594
rect 519368 360514 519488 360530
rect 519368 360450 519396 360514
rect 519460 360450 519488 360514
rect 519368 360434 519488 360450
rect 519368 360370 519396 360434
rect 519460 360370 519488 360434
rect 519368 360354 519488 360370
rect 519368 360290 519396 360354
rect 519460 360290 519488 360354
rect 519368 360274 519488 360290
rect 519368 360210 519396 360274
rect 519460 360210 519488 360274
rect 519368 360194 519488 360210
rect 519368 360130 519396 360194
rect 519460 360130 519488 360194
rect 519368 360114 519488 360130
rect 519368 360050 519396 360114
rect 519460 360050 519488 360114
rect 519368 360034 519488 360050
rect 519368 359970 519396 360034
rect 519460 359970 519488 360034
rect 519368 359954 519488 359970
rect 519368 359890 519396 359954
rect 519460 359890 519488 359954
rect 519368 359866 519488 359890
rect 523128 361474 523248 361498
rect 523128 361410 523156 361474
rect 523220 361410 523248 361474
rect 523128 361394 523248 361410
rect 523128 361330 523156 361394
rect 523220 361330 523248 361394
rect 523128 361314 523248 361330
rect 523128 361250 523156 361314
rect 523220 361250 523248 361314
rect 523128 361234 523248 361250
rect 523128 361170 523156 361234
rect 523220 361170 523248 361234
rect 523128 361154 523248 361170
rect 523128 361090 523156 361154
rect 523220 361090 523248 361154
rect 523128 361074 523248 361090
rect 523128 361010 523156 361074
rect 523220 361010 523248 361074
rect 523128 360994 523248 361010
rect 523128 360930 523156 360994
rect 523220 360930 523248 360994
rect 523128 360914 523248 360930
rect 523128 360850 523156 360914
rect 523220 360850 523248 360914
rect 523128 360834 523248 360850
rect 523128 360770 523156 360834
rect 523220 360770 523248 360834
rect 523128 360754 523248 360770
rect 523128 360690 523156 360754
rect 523220 360690 523248 360754
rect 523128 360674 523248 360690
rect 523128 360610 523156 360674
rect 523220 360610 523248 360674
rect 523128 360594 523248 360610
rect 523128 360530 523156 360594
rect 523220 360530 523248 360594
rect 523128 360514 523248 360530
rect 523128 360450 523156 360514
rect 523220 360450 523248 360514
rect 523128 360434 523248 360450
rect 523128 360370 523156 360434
rect 523220 360370 523248 360434
rect 523128 360354 523248 360370
rect 523128 360290 523156 360354
rect 523220 360290 523248 360354
rect 523128 360274 523248 360290
rect 523128 360210 523156 360274
rect 523220 360210 523248 360274
rect 523128 360194 523248 360210
rect 523128 360130 523156 360194
rect 523220 360130 523248 360194
rect 523128 360114 523248 360130
rect 523128 360050 523156 360114
rect 523220 360050 523248 360114
rect 523128 360034 523248 360050
rect 523128 359970 523156 360034
rect 523220 359970 523248 360034
rect 523128 359954 523248 359970
rect 523128 359890 523156 359954
rect 523220 359890 523248 359954
rect 523128 359866 523248 359890
rect 526888 361474 527008 361498
rect 526888 361410 526916 361474
rect 526980 361410 527008 361474
rect 526888 361394 527008 361410
rect 526888 361330 526916 361394
rect 526980 361330 527008 361394
rect 526888 361314 527008 361330
rect 526888 361250 526916 361314
rect 526980 361250 527008 361314
rect 526888 361234 527008 361250
rect 526888 361170 526916 361234
rect 526980 361170 527008 361234
rect 526888 361154 527008 361170
rect 526888 361090 526916 361154
rect 526980 361090 527008 361154
rect 526888 361074 527008 361090
rect 526888 361010 526916 361074
rect 526980 361010 527008 361074
rect 526888 360994 527008 361010
rect 526888 360930 526916 360994
rect 526980 360930 527008 360994
rect 526888 360914 527008 360930
rect 526888 360850 526916 360914
rect 526980 360850 527008 360914
rect 526888 360834 527008 360850
rect 526888 360770 526916 360834
rect 526980 360770 527008 360834
rect 526888 360754 527008 360770
rect 526888 360690 526916 360754
rect 526980 360690 527008 360754
rect 526888 360674 527008 360690
rect 526888 360610 526916 360674
rect 526980 360610 527008 360674
rect 526888 360594 527008 360610
rect 526888 360530 526916 360594
rect 526980 360530 527008 360594
rect 526888 360514 527008 360530
rect 526888 360450 526916 360514
rect 526980 360450 527008 360514
rect 526888 360434 527008 360450
rect 526888 360370 526916 360434
rect 526980 360370 527008 360434
rect 526888 360354 527008 360370
rect 526888 360290 526916 360354
rect 526980 360290 527008 360354
rect 526888 360274 527008 360290
rect 526888 360210 526916 360274
rect 526980 360210 527008 360274
rect 526888 360194 527008 360210
rect 526888 360130 526916 360194
rect 526980 360130 527008 360194
rect 526888 360114 527008 360130
rect 526888 360050 526916 360114
rect 526980 360050 527008 360114
rect 526888 360034 527008 360050
rect 526888 359970 526916 360034
rect 526980 359970 527008 360034
rect 526888 359954 527008 359970
rect 526888 359890 526916 359954
rect 526980 359890 527008 359954
rect 526888 359866 527008 359890
rect 530648 361474 530768 361498
rect 530648 361410 530676 361474
rect 530740 361410 530768 361474
rect 530648 361394 530768 361410
rect 530648 361330 530676 361394
rect 530740 361330 530768 361394
rect 530648 361314 530768 361330
rect 530648 361250 530676 361314
rect 530740 361250 530768 361314
rect 530648 361234 530768 361250
rect 530648 361170 530676 361234
rect 530740 361170 530768 361234
rect 530648 361154 530768 361170
rect 530648 361090 530676 361154
rect 530740 361090 530768 361154
rect 530648 361074 530768 361090
rect 530648 361010 530676 361074
rect 530740 361010 530768 361074
rect 530648 360994 530768 361010
rect 530648 360930 530676 360994
rect 530740 360930 530768 360994
rect 530648 360914 530768 360930
rect 530648 360850 530676 360914
rect 530740 360850 530768 360914
rect 530648 360834 530768 360850
rect 530648 360770 530676 360834
rect 530740 360770 530768 360834
rect 530648 360754 530768 360770
rect 530648 360690 530676 360754
rect 530740 360690 530768 360754
rect 530648 360674 530768 360690
rect 530648 360610 530676 360674
rect 530740 360610 530768 360674
rect 530648 360594 530768 360610
rect 530648 360530 530676 360594
rect 530740 360530 530768 360594
rect 530648 360514 530768 360530
rect 530648 360450 530676 360514
rect 530740 360450 530768 360514
rect 530648 360434 530768 360450
rect 530648 360370 530676 360434
rect 530740 360370 530768 360434
rect 530648 360354 530768 360370
rect 530648 360290 530676 360354
rect 530740 360290 530768 360354
rect 530648 360274 530768 360290
rect 530648 360210 530676 360274
rect 530740 360210 530768 360274
rect 530648 360194 530768 360210
rect 530648 360130 530676 360194
rect 530740 360130 530768 360194
rect 530648 360114 530768 360130
rect 530648 360050 530676 360114
rect 530740 360050 530768 360114
rect 530648 360034 530768 360050
rect 530648 359970 530676 360034
rect 530740 359970 530768 360034
rect 530648 359954 530768 359970
rect 530648 359890 530676 359954
rect 530740 359890 530768 359954
rect 530648 359866 530768 359890
rect 534408 361474 534528 361498
rect 534408 361410 534436 361474
rect 534500 361410 534528 361474
rect 534408 361394 534528 361410
rect 534408 361330 534436 361394
rect 534500 361330 534528 361394
rect 534408 361314 534528 361330
rect 534408 361250 534436 361314
rect 534500 361250 534528 361314
rect 534408 361234 534528 361250
rect 534408 361170 534436 361234
rect 534500 361170 534528 361234
rect 534408 361154 534528 361170
rect 534408 361090 534436 361154
rect 534500 361090 534528 361154
rect 534408 361074 534528 361090
rect 534408 361010 534436 361074
rect 534500 361010 534528 361074
rect 534408 360994 534528 361010
rect 534408 360930 534436 360994
rect 534500 360930 534528 360994
rect 534408 360914 534528 360930
rect 534408 360850 534436 360914
rect 534500 360850 534528 360914
rect 534408 360834 534528 360850
rect 534408 360770 534436 360834
rect 534500 360770 534528 360834
rect 534408 360754 534528 360770
rect 534408 360690 534436 360754
rect 534500 360690 534528 360754
rect 534408 360674 534528 360690
rect 534408 360610 534436 360674
rect 534500 360610 534528 360674
rect 534408 360594 534528 360610
rect 534408 360530 534436 360594
rect 534500 360530 534528 360594
rect 534408 360514 534528 360530
rect 534408 360450 534436 360514
rect 534500 360450 534528 360514
rect 534408 360434 534528 360450
rect 534408 360370 534436 360434
rect 534500 360370 534528 360434
rect 534408 360354 534528 360370
rect 534408 360290 534436 360354
rect 534500 360290 534528 360354
rect 534408 360274 534528 360290
rect 534408 360210 534436 360274
rect 534500 360210 534528 360274
rect 534408 360194 534528 360210
rect 534408 360130 534436 360194
rect 534500 360130 534528 360194
rect 534408 360114 534528 360130
rect 534408 360050 534436 360114
rect 534500 360050 534528 360114
rect 534408 360034 534528 360050
rect 534408 359970 534436 360034
rect 534500 359970 534528 360034
rect 534408 359954 534528 359970
rect 534408 359890 534436 359954
rect 534500 359890 534528 359954
rect 534408 359866 534528 359890
rect 545023 359903 545141 380497
rect 566264 359978 566510 359983
rect 566264 359903 566274 359978
rect 545023 359786 566274 359903
rect 566500 359903 566510 359978
rect 580242 359906 580368 359911
rect 580242 359903 580252 359906
rect 566500 359786 580252 359903
rect 580358 359903 580368 359906
rect 580358 359786 580941 359903
rect 545023 359785 580941 359786
rect 566264 359781 566510 359785
rect 580242 359781 580368 359785
rect 491168 359026 491288 359050
rect 491168 358962 491196 359026
rect 491260 358962 491288 359026
rect 491168 358946 491288 358962
rect 491168 358882 491196 358946
rect 491260 358882 491288 358946
rect 491168 358866 491288 358882
rect 491168 358802 491196 358866
rect 491260 358802 491288 358866
rect 491168 358786 491288 358802
rect 491168 358722 491196 358786
rect 491260 358722 491288 358786
rect 491168 358706 491288 358722
rect 491168 358642 491196 358706
rect 491260 358642 491288 358706
rect 491168 358626 491288 358642
rect 491168 358562 491196 358626
rect 491260 358562 491288 358626
rect 491168 358546 491288 358562
rect 491168 358482 491196 358546
rect 491260 358482 491288 358546
rect 491168 358466 491288 358482
rect 491168 358402 491196 358466
rect 491260 358402 491288 358466
rect 491168 358386 491288 358402
rect 491168 358322 491196 358386
rect 491260 358322 491288 358386
rect 491168 358306 491288 358322
rect 491168 358242 491196 358306
rect 491260 358242 491288 358306
rect 491168 358226 491288 358242
rect 491168 358162 491196 358226
rect 491260 358162 491288 358226
rect 491168 358146 491288 358162
rect 491168 358082 491196 358146
rect 491260 358082 491288 358146
rect 491168 358066 491288 358082
rect 491168 358002 491196 358066
rect 491260 358002 491288 358066
rect 491168 357986 491288 358002
rect 491168 357922 491196 357986
rect 491260 357922 491288 357986
rect 491168 357906 491288 357922
rect 491168 357842 491196 357906
rect 491260 357842 491288 357906
rect 491168 357826 491288 357842
rect 491168 357762 491196 357826
rect 491260 357762 491288 357826
rect 491168 357746 491288 357762
rect 491168 357682 491196 357746
rect 491260 357682 491288 357746
rect 491168 357666 491288 357682
rect 491168 357602 491196 357666
rect 491260 357602 491288 357666
rect 491168 357586 491288 357602
rect 491168 357522 491196 357586
rect 491260 357522 491288 357586
rect 491168 357506 491288 357522
rect 491168 357442 491196 357506
rect 491260 357442 491288 357506
rect 491168 357418 491288 357442
rect 494928 359026 495048 359050
rect 494928 358962 494956 359026
rect 495020 358962 495048 359026
rect 494928 358946 495048 358962
rect 494928 358882 494956 358946
rect 495020 358882 495048 358946
rect 494928 358866 495048 358882
rect 494928 358802 494956 358866
rect 495020 358802 495048 358866
rect 494928 358786 495048 358802
rect 494928 358722 494956 358786
rect 495020 358722 495048 358786
rect 494928 358706 495048 358722
rect 494928 358642 494956 358706
rect 495020 358642 495048 358706
rect 494928 358626 495048 358642
rect 494928 358562 494956 358626
rect 495020 358562 495048 358626
rect 494928 358546 495048 358562
rect 494928 358482 494956 358546
rect 495020 358482 495048 358546
rect 494928 358466 495048 358482
rect 494928 358402 494956 358466
rect 495020 358402 495048 358466
rect 494928 358386 495048 358402
rect 494928 358322 494956 358386
rect 495020 358322 495048 358386
rect 494928 358306 495048 358322
rect 494928 358242 494956 358306
rect 495020 358242 495048 358306
rect 494928 358226 495048 358242
rect 494928 358162 494956 358226
rect 495020 358162 495048 358226
rect 494928 358146 495048 358162
rect 494928 358082 494956 358146
rect 495020 358082 495048 358146
rect 494928 358066 495048 358082
rect 494928 358002 494956 358066
rect 495020 358002 495048 358066
rect 494928 357986 495048 358002
rect 494928 357922 494956 357986
rect 495020 357922 495048 357986
rect 494928 357906 495048 357922
rect 494928 357842 494956 357906
rect 495020 357842 495048 357906
rect 494928 357826 495048 357842
rect 494928 357762 494956 357826
rect 495020 357762 495048 357826
rect 494928 357746 495048 357762
rect 494928 357682 494956 357746
rect 495020 357682 495048 357746
rect 494928 357666 495048 357682
rect 494928 357602 494956 357666
rect 495020 357602 495048 357666
rect 494928 357586 495048 357602
rect 494928 357522 494956 357586
rect 495020 357522 495048 357586
rect 494928 357506 495048 357522
rect 494928 357442 494956 357506
rect 495020 357442 495048 357506
rect 494928 357418 495048 357442
rect 498688 359026 498808 359050
rect 498688 358962 498716 359026
rect 498780 358962 498808 359026
rect 498688 358946 498808 358962
rect 498688 358882 498716 358946
rect 498780 358882 498808 358946
rect 498688 358866 498808 358882
rect 498688 358802 498716 358866
rect 498780 358802 498808 358866
rect 498688 358786 498808 358802
rect 498688 358722 498716 358786
rect 498780 358722 498808 358786
rect 498688 358706 498808 358722
rect 498688 358642 498716 358706
rect 498780 358642 498808 358706
rect 498688 358626 498808 358642
rect 498688 358562 498716 358626
rect 498780 358562 498808 358626
rect 498688 358546 498808 358562
rect 498688 358482 498716 358546
rect 498780 358482 498808 358546
rect 498688 358466 498808 358482
rect 498688 358402 498716 358466
rect 498780 358402 498808 358466
rect 498688 358386 498808 358402
rect 498688 358322 498716 358386
rect 498780 358322 498808 358386
rect 498688 358306 498808 358322
rect 498688 358242 498716 358306
rect 498780 358242 498808 358306
rect 498688 358226 498808 358242
rect 498688 358162 498716 358226
rect 498780 358162 498808 358226
rect 498688 358146 498808 358162
rect 498688 358082 498716 358146
rect 498780 358082 498808 358146
rect 498688 358066 498808 358082
rect 498688 358002 498716 358066
rect 498780 358002 498808 358066
rect 498688 357986 498808 358002
rect 498688 357922 498716 357986
rect 498780 357922 498808 357986
rect 498688 357906 498808 357922
rect 498688 357842 498716 357906
rect 498780 357842 498808 357906
rect 498688 357826 498808 357842
rect 498688 357762 498716 357826
rect 498780 357762 498808 357826
rect 498688 357746 498808 357762
rect 498688 357682 498716 357746
rect 498780 357682 498808 357746
rect 498688 357666 498808 357682
rect 498688 357602 498716 357666
rect 498780 357602 498808 357666
rect 498688 357586 498808 357602
rect 498688 357522 498716 357586
rect 498780 357522 498808 357586
rect 498688 357506 498808 357522
rect 498688 357442 498716 357506
rect 498780 357442 498808 357506
rect 498688 357418 498808 357442
rect 502448 359026 502568 359050
rect 502448 358962 502476 359026
rect 502540 358962 502568 359026
rect 502448 358946 502568 358962
rect 502448 358882 502476 358946
rect 502540 358882 502568 358946
rect 502448 358866 502568 358882
rect 502448 358802 502476 358866
rect 502540 358802 502568 358866
rect 502448 358786 502568 358802
rect 502448 358722 502476 358786
rect 502540 358722 502568 358786
rect 502448 358706 502568 358722
rect 502448 358642 502476 358706
rect 502540 358642 502568 358706
rect 502448 358626 502568 358642
rect 502448 358562 502476 358626
rect 502540 358562 502568 358626
rect 502448 358546 502568 358562
rect 502448 358482 502476 358546
rect 502540 358482 502568 358546
rect 502448 358466 502568 358482
rect 502448 358402 502476 358466
rect 502540 358402 502568 358466
rect 502448 358386 502568 358402
rect 502448 358322 502476 358386
rect 502540 358322 502568 358386
rect 502448 358306 502568 358322
rect 502448 358242 502476 358306
rect 502540 358242 502568 358306
rect 502448 358226 502568 358242
rect 502448 358162 502476 358226
rect 502540 358162 502568 358226
rect 502448 358146 502568 358162
rect 502448 358082 502476 358146
rect 502540 358082 502568 358146
rect 502448 358066 502568 358082
rect 502448 358002 502476 358066
rect 502540 358002 502568 358066
rect 502448 357986 502568 358002
rect 502448 357922 502476 357986
rect 502540 357922 502568 357986
rect 502448 357906 502568 357922
rect 502448 357842 502476 357906
rect 502540 357842 502568 357906
rect 502448 357826 502568 357842
rect 502448 357762 502476 357826
rect 502540 357762 502568 357826
rect 502448 357746 502568 357762
rect 502448 357682 502476 357746
rect 502540 357682 502568 357746
rect 502448 357666 502568 357682
rect 502448 357602 502476 357666
rect 502540 357602 502568 357666
rect 502448 357586 502568 357602
rect 502448 357522 502476 357586
rect 502540 357522 502568 357586
rect 502448 357506 502568 357522
rect 502448 357442 502476 357506
rect 502540 357442 502568 357506
rect 502448 357418 502568 357442
rect 506208 359026 506328 359050
rect 506208 358962 506236 359026
rect 506300 358962 506328 359026
rect 506208 358946 506328 358962
rect 506208 358882 506236 358946
rect 506300 358882 506328 358946
rect 506208 358866 506328 358882
rect 506208 358802 506236 358866
rect 506300 358802 506328 358866
rect 506208 358786 506328 358802
rect 506208 358722 506236 358786
rect 506300 358722 506328 358786
rect 506208 358706 506328 358722
rect 506208 358642 506236 358706
rect 506300 358642 506328 358706
rect 506208 358626 506328 358642
rect 506208 358562 506236 358626
rect 506300 358562 506328 358626
rect 506208 358546 506328 358562
rect 506208 358482 506236 358546
rect 506300 358482 506328 358546
rect 506208 358466 506328 358482
rect 506208 358402 506236 358466
rect 506300 358402 506328 358466
rect 506208 358386 506328 358402
rect 506208 358322 506236 358386
rect 506300 358322 506328 358386
rect 506208 358306 506328 358322
rect 506208 358242 506236 358306
rect 506300 358242 506328 358306
rect 506208 358226 506328 358242
rect 506208 358162 506236 358226
rect 506300 358162 506328 358226
rect 506208 358146 506328 358162
rect 506208 358082 506236 358146
rect 506300 358082 506328 358146
rect 506208 358066 506328 358082
rect 506208 358002 506236 358066
rect 506300 358002 506328 358066
rect 506208 357986 506328 358002
rect 506208 357922 506236 357986
rect 506300 357922 506328 357986
rect 506208 357906 506328 357922
rect 506208 357842 506236 357906
rect 506300 357842 506328 357906
rect 506208 357826 506328 357842
rect 506208 357762 506236 357826
rect 506300 357762 506328 357826
rect 506208 357746 506328 357762
rect 506208 357682 506236 357746
rect 506300 357682 506328 357746
rect 506208 357666 506328 357682
rect 506208 357602 506236 357666
rect 506300 357602 506328 357666
rect 506208 357586 506328 357602
rect 506208 357522 506236 357586
rect 506300 357522 506328 357586
rect 506208 357506 506328 357522
rect 506208 357442 506236 357506
rect 506300 357442 506328 357506
rect 506208 357418 506328 357442
rect 509968 359026 510088 359050
rect 509968 358962 509996 359026
rect 510060 358962 510088 359026
rect 509968 358946 510088 358962
rect 509968 358882 509996 358946
rect 510060 358882 510088 358946
rect 509968 358866 510088 358882
rect 509968 358802 509996 358866
rect 510060 358802 510088 358866
rect 509968 358786 510088 358802
rect 509968 358722 509996 358786
rect 510060 358722 510088 358786
rect 509968 358706 510088 358722
rect 509968 358642 509996 358706
rect 510060 358642 510088 358706
rect 509968 358626 510088 358642
rect 509968 358562 509996 358626
rect 510060 358562 510088 358626
rect 509968 358546 510088 358562
rect 509968 358482 509996 358546
rect 510060 358482 510088 358546
rect 509968 358466 510088 358482
rect 509968 358402 509996 358466
rect 510060 358402 510088 358466
rect 509968 358386 510088 358402
rect 509968 358322 509996 358386
rect 510060 358322 510088 358386
rect 509968 358306 510088 358322
rect 509968 358242 509996 358306
rect 510060 358242 510088 358306
rect 509968 358226 510088 358242
rect 509968 358162 509996 358226
rect 510060 358162 510088 358226
rect 509968 358146 510088 358162
rect 509968 358082 509996 358146
rect 510060 358082 510088 358146
rect 509968 358066 510088 358082
rect 509968 358002 509996 358066
rect 510060 358002 510088 358066
rect 509968 357986 510088 358002
rect 509968 357922 509996 357986
rect 510060 357922 510088 357986
rect 509968 357906 510088 357922
rect 509968 357842 509996 357906
rect 510060 357842 510088 357906
rect 509968 357826 510088 357842
rect 509968 357762 509996 357826
rect 510060 357762 510088 357826
rect 509968 357746 510088 357762
rect 509968 357682 509996 357746
rect 510060 357682 510088 357746
rect 509968 357666 510088 357682
rect 509968 357602 509996 357666
rect 510060 357602 510088 357666
rect 509968 357586 510088 357602
rect 509968 357522 509996 357586
rect 510060 357522 510088 357586
rect 509968 357506 510088 357522
rect 509968 357442 509996 357506
rect 510060 357442 510088 357506
rect 509968 357418 510088 357442
rect 513728 359026 513848 359050
rect 513728 358962 513756 359026
rect 513820 358962 513848 359026
rect 513728 358946 513848 358962
rect 513728 358882 513756 358946
rect 513820 358882 513848 358946
rect 513728 358866 513848 358882
rect 513728 358802 513756 358866
rect 513820 358802 513848 358866
rect 513728 358786 513848 358802
rect 513728 358722 513756 358786
rect 513820 358722 513848 358786
rect 513728 358706 513848 358722
rect 513728 358642 513756 358706
rect 513820 358642 513848 358706
rect 513728 358626 513848 358642
rect 513728 358562 513756 358626
rect 513820 358562 513848 358626
rect 513728 358546 513848 358562
rect 513728 358482 513756 358546
rect 513820 358482 513848 358546
rect 513728 358466 513848 358482
rect 513728 358402 513756 358466
rect 513820 358402 513848 358466
rect 513728 358386 513848 358402
rect 513728 358322 513756 358386
rect 513820 358322 513848 358386
rect 513728 358306 513848 358322
rect 513728 358242 513756 358306
rect 513820 358242 513848 358306
rect 513728 358226 513848 358242
rect 513728 358162 513756 358226
rect 513820 358162 513848 358226
rect 513728 358146 513848 358162
rect 513728 358082 513756 358146
rect 513820 358082 513848 358146
rect 513728 358066 513848 358082
rect 513728 358002 513756 358066
rect 513820 358002 513848 358066
rect 513728 357986 513848 358002
rect 513728 357922 513756 357986
rect 513820 357922 513848 357986
rect 513728 357906 513848 357922
rect 513728 357842 513756 357906
rect 513820 357842 513848 357906
rect 513728 357826 513848 357842
rect 513728 357762 513756 357826
rect 513820 357762 513848 357826
rect 513728 357746 513848 357762
rect 513728 357682 513756 357746
rect 513820 357682 513848 357746
rect 513728 357666 513848 357682
rect 513728 357602 513756 357666
rect 513820 357602 513848 357666
rect 513728 357586 513848 357602
rect 513728 357522 513756 357586
rect 513820 357522 513848 357586
rect 513728 357506 513848 357522
rect 513728 357442 513756 357506
rect 513820 357442 513848 357506
rect 513728 357418 513848 357442
rect 517488 359026 517608 359050
rect 517488 358962 517516 359026
rect 517580 358962 517608 359026
rect 517488 358946 517608 358962
rect 517488 358882 517516 358946
rect 517580 358882 517608 358946
rect 517488 358866 517608 358882
rect 517488 358802 517516 358866
rect 517580 358802 517608 358866
rect 517488 358786 517608 358802
rect 517488 358722 517516 358786
rect 517580 358722 517608 358786
rect 517488 358706 517608 358722
rect 517488 358642 517516 358706
rect 517580 358642 517608 358706
rect 517488 358626 517608 358642
rect 517488 358562 517516 358626
rect 517580 358562 517608 358626
rect 517488 358546 517608 358562
rect 517488 358482 517516 358546
rect 517580 358482 517608 358546
rect 517488 358466 517608 358482
rect 517488 358402 517516 358466
rect 517580 358402 517608 358466
rect 517488 358386 517608 358402
rect 517488 358322 517516 358386
rect 517580 358322 517608 358386
rect 517488 358306 517608 358322
rect 517488 358242 517516 358306
rect 517580 358242 517608 358306
rect 517488 358226 517608 358242
rect 517488 358162 517516 358226
rect 517580 358162 517608 358226
rect 517488 358146 517608 358162
rect 517488 358082 517516 358146
rect 517580 358082 517608 358146
rect 517488 358066 517608 358082
rect 517488 358002 517516 358066
rect 517580 358002 517608 358066
rect 517488 357986 517608 358002
rect 517488 357922 517516 357986
rect 517580 357922 517608 357986
rect 517488 357906 517608 357922
rect 517488 357842 517516 357906
rect 517580 357842 517608 357906
rect 517488 357826 517608 357842
rect 517488 357762 517516 357826
rect 517580 357762 517608 357826
rect 517488 357746 517608 357762
rect 517488 357682 517516 357746
rect 517580 357682 517608 357746
rect 517488 357666 517608 357682
rect 517488 357602 517516 357666
rect 517580 357602 517608 357666
rect 517488 357586 517608 357602
rect 517488 357522 517516 357586
rect 517580 357522 517608 357586
rect 517488 357506 517608 357522
rect 517488 357442 517516 357506
rect 517580 357442 517608 357506
rect 517488 357418 517608 357442
rect 521248 359026 521368 359050
rect 521248 358962 521276 359026
rect 521340 358962 521368 359026
rect 521248 358946 521368 358962
rect 521248 358882 521276 358946
rect 521340 358882 521368 358946
rect 521248 358866 521368 358882
rect 521248 358802 521276 358866
rect 521340 358802 521368 358866
rect 521248 358786 521368 358802
rect 521248 358722 521276 358786
rect 521340 358722 521368 358786
rect 521248 358706 521368 358722
rect 521248 358642 521276 358706
rect 521340 358642 521368 358706
rect 521248 358626 521368 358642
rect 521248 358562 521276 358626
rect 521340 358562 521368 358626
rect 521248 358546 521368 358562
rect 521248 358482 521276 358546
rect 521340 358482 521368 358546
rect 521248 358466 521368 358482
rect 521248 358402 521276 358466
rect 521340 358402 521368 358466
rect 521248 358386 521368 358402
rect 521248 358322 521276 358386
rect 521340 358322 521368 358386
rect 521248 358306 521368 358322
rect 521248 358242 521276 358306
rect 521340 358242 521368 358306
rect 521248 358226 521368 358242
rect 521248 358162 521276 358226
rect 521340 358162 521368 358226
rect 521248 358146 521368 358162
rect 521248 358082 521276 358146
rect 521340 358082 521368 358146
rect 521248 358066 521368 358082
rect 521248 358002 521276 358066
rect 521340 358002 521368 358066
rect 521248 357986 521368 358002
rect 521248 357922 521276 357986
rect 521340 357922 521368 357986
rect 521248 357906 521368 357922
rect 521248 357842 521276 357906
rect 521340 357842 521368 357906
rect 521248 357826 521368 357842
rect 521248 357762 521276 357826
rect 521340 357762 521368 357826
rect 521248 357746 521368 357762
rect 521248 357682 521276 357746
rect 521340 357682 521368 357746
rect 521248 357666 521368 357682
rect 521248 357602 521276 357666
rect 521340 357602 521368 357666
rect 521248 357586 521368 357602
rect 521248 357522 521276 357586
rect 521340 357522 521368 357586
rect 521248 357506 521368 357522
rect 521248 357442 521276 357506
rect 521340 357442 521368 357506
rect 521248 357418 521368 357442
rect 525008 359026 525128 359050
rect 525008 358962 525036 359026
rect 525100 358962 525128 359026
rect 525008 358946 525128 358962
rect 525008 358882 525036 358946
rect 525100 358882 525128 358946
rect 525008 358866 525128 358882
rect 525008 358802 525036 358866
rect 525100 358802 525128 358866
rect 525008 358786 525128 358802
rect 525008 358722 525036 358786
rect 525100 358722 525128 358786
rect 525008 358706 525128 358722
rect 525008 358642 525036 358706
rect 525100 358642 525128 358706
rect 525008 358626 525128 358642
rect 525008 358562 525036 358626
rect 525100 358562 525128 358626
rect 525008 358546 525128 358562
rect 525008 358482 525036 358546
rect 525100 358482 525128 358546
rect 525008 358466 525128 358482
rect 525008 358402 525036 358466
rect 525100 358402 525128 358466
rect 525008 358386 525128 358402
rect 525008 358322 525036 358386
rect 525100 358322 525128 358386
rect 525008 358306 525128 358322
rect 525008 358242 525036 358306
rect 525100 358242 525128 358306
rect 525008 358226 525128 358242
rect 525008 358162 525036 358226
rect 525100 358162 525128 358226
rect 525008 358146 525128 358162
rect 525008 358082 525036 358146
rect 525100 358082 525128 358146
rect 525008 358066 525128 358082
rect 525008 358002 525036 358066
rect 525100 358002 525128 358066
rect 525008 357986 525128 358002
rect 525008 357922 525036 357986
rect 525100 357922 525128 357986
rect 525008 357906 525128 357922
rect 525008 357842 525036 357906
rect 525100 357842 525128 357906
rect 525008 357826 525128 357842
rect 525008 357762 525036 357826
rect 525100 357762 525128 357826
rect 525008 357746 525128 357762
rect 525008 357682 525036 357746
rect 525100 357682 525128 357746
rect 525008 357666 525128 357682
rect 525008 357602 525036 357666
rect 525100 357602 525128 357666
rect 525008 357586 525128 357602
rect 525008 357522 525036 357586
rect 525100 357522 525128 357586
rect 525008 357506 525128 357522
rect 525008 357442 525036 357506
rect 525100 357442 525128 357506
rect 525008 357418 525128 357442
rect 528768 359026 528888 359050
rect 528768 358962 528796 359026
rect 528860 358962 528888 359026
rect 528768 358946 528888 358962
rect 528768 358882 528796 358946
rect 528860 358882 528888 358946
rect 528768 358866 528888 358882
rect 528768 358802 528796 358866
rect 528860 358802 528888 358866
rect 528768 358786 528888 358802
rect 528768 358722 528796 358786
rect 528860 358722 528888 358786
rect 528768 358706 528888 358722
rect 528768 358642 528796 358706
rect 528860 358642 528888 358706
rect 528768 358626 528888 358642
rect 528768 358562 528796 358626
rect 528860 358562 528888 358626
rect 528768 358546 528888 358562
rect 528768 358482 528796 358546
rect 528860 358482 528888 358546
rect 528768 358466 528888 358482
rect 528768 358402 528796 358466
rect 528860 358402 528888 358466
rect 528768 358386 528888 358402
rect 528768 358322 528796 358386
rect 528860 358322 528888 358386
rect 528768 358306 528888 358322
rect 528768 358242 528796 358306
rect 528860 358242 528888 358306
rect 528768 358226 528888 358242
rect 528768 358162 528796 358226
rect 528860 358162 528888 358226
rect 528768 358146 528888 358162
rect 528768 358082 528796 358146
rect 528860 358082 528888 358146
rect 528768 358066 528888 358082
rect 528768 358002 528796 358066
rect 528860 358002 528888 358066
rect 528768 357986 528888 358002
rect 528768 357922 528796 357986
rect 528860 357922 528888 357986
rect 528768 357906 528888 357922
rect 528768 357842 528796 357906
rect 528860 357842 528888 357906
rect 528768 357826 528888 357842
rect 528768 357762 528796 357826
rect 528860 357762 528888 357826
rect 528768 357746 528888 357762
rect 528768 357682 528796 357746
rect 528860 357682 528888 357746
rect 528768 357666 528888 357682
rect 528768 357602 528796 357666
rect 528860 357602 528888 357666
rect 528768 357586 528888 357602
rect 528768 357522 528796 357586
rect 528860 357522 528888 357586
rect 528768 357506 528888 357522
rect 528768 357442 528796 357506
rect 528860 357442 528888 357506
rect 528768 357418 528888 357442
rect 532528 359026 532648 359050
rect 532528 358962 532556 359026
rect 532620 358962 532648 359026
rect 532528 358946 532648 358962
rect 532528 358882 532556 358946
rect 532620 358882 532648 358946
rect 532528 358866 532648 358882
rect 532528 358802 532556 358866
rect 532620 358802 532648 358866
rect 532528 358786 532648 358802
rect 532528 358722 532556 358786
rect 532620 358722 532648 358786
rect 532528 358706 532648 358722
rect 532528 358642 532556 358706
rect 532620 358642 532648 358706
rect 532528 358626 532648 358642
rect 532528 358562 532556 358626
rect 532620 358562 532648 358626
rect 532528 358546 532648 358562
rect 532528 358482 532556 358546
rect 532620 358482 532648 358546
rect 532528 358466 532648 358482
rect 532528 358402 532556 358466
rect 532620 358402 532648 358466
rect 532528 358386 532648 358402
rect 532528 358322 532556 358386
rect 532620 358322 532648 358386
rect 532528 358306 532648 358322
rect 532528 358242 532556 358306
rect 532620 358242 532648 358306
rect 532528 358226 532648 358242
rect 532528 358162 532556 358226
rect 532620 358162 532648 358226
rect 532528 358146 532648 358162
rect 532528 358082 532556 358146
rect 532620 358082 532648 358146
rect 532528 358066 532648 358082
rect 532528 358002 532556 358066
rect 532620 358002 532648 358066
rect 532528 357986 532648 358002
rect 532528 357922 532556 357986
rect 532620 357922 532648 357986
rect 532528 357906 532648 357922
rect 532528 357842 532556 357906
rect 532620 357842 532648 357906
rect 532528 357826 532648 357842
rect 532528 357762 532556 357826
rect 532620 357762 532648 357826
rect 532528 357746 532648 357762
rect 532528 357682 532556 357746
rect 532620 357682 532648 357746
rect 532528 357666 532648 357682
rect 532528 357602 532556 357666
rect 532620 357602 532648 357666
rect 532528 357586 532648 357602
rect 532528 357522 532556 357586
rect 532620 357522 532648 357586
rect 532528 357506 532648 357522
rect 532528 357442 532556 357506
rect 532620 357442 532648 357506
rect 532528 357418 532648 357442
rect 536288 359026 536408 359050
rect 536288 358962 536316 359026
rect 536380 358962 536408 359026
rect 536288 358946 536408 358962
rect 536288 358882 536316 358946
rect 536380 358882 536408 358946
rect 536288 358866 536408 358882
rect 536288 358802 536316 358866
rect 536380 358802 536408 358866
rect 580823 358984 580941 359785
rect 580823 358866 583840 358984
rect 580823 358859 580941 358866
rect 536288 358786 536408 358802
rect 536288 358722 536316 358786
rect 536380 358722 536408 358786
rect 536288 358706 536408 358722
rect 536288 358642 536316 358706
rect 536380 358642 536408 358706
rect 536288 358626 536408 358642
rect 536288 358562 536316 358626
rect 536380 358562 536408 358626
rect 536288 358546 536408 358562
rect 536288 358482 536316 358546
rect 536380 358482 536408 358546
rect 536288 358466 536408 358482
rect 536288 358402 536316 358466
rect 536380 358402 536408 358466
rect 536288 358386 536408 358402
rect 536288 358322 536316 358386
rect 536380 358322 536408 358386
rect 536288 358306 536408 358322
rect 536288 358242 536316 358306
rect 536380 358242 536408 358306
rect 536288 358226 536408 358242
rect 536288 358162 536316 358226
rect 536380 358162 536408 358226
rect 536288 358146 536408 358162
rect 536288 358082 536316 358146
rect 536380 358082 536408 358146
rect 536288 358066 536408 358082
rect 536288 358002 536316 358066
rect 536380 358002 536408 358066
rect 536288 357986 536408 358002
rect 536288 357922 536316 357986
rect 536380 357922 536408 357986
rect 536288 357906 536408 357922
rect 536288 357842 536316 357906
rect 536380 357842 536408 357906
rect 536288 357826 536408 357842
rect 559702 358052 559930 358057
rect 559702 357844 559712 358052
rect 559920 357844 559930 358052
rect 559702 357839 559930 357844
rect 573530 357920 573888 357925
rect 536288 357762 536316 357826
rect 536380 357762 536408 357826
rect 536288 357746 536408 357762
rect 536288 357682 536316 357746
rect 536380 357682 536408 357746
rect 536288 357666 536408 357682
rect 536288 357602 536316 357666
rect 536380 357602 536408 357666
rect 536288 357586 536408 357602
rect 573530 357594 573540 357920
rect 573878 357594 573888 357920
rect 573530 357589 573888 357594
rect 536288 357522 536316 357586
rect 536380 357522 536408 357586
rect 536288 357506 536408 357522
rect 536288 357442 536316 357506
rect 536380 357442 536408 357506
rect 536288 357418 536408 357442
rect 508335 356582 509603 356589
rect 508335 356446 508362 356582
rect 508652 356446 509603 356582
rect 508335 356375 509603 356446
rect 509393 313770 509603 356375
rect 566116 313804 566356 313809
rect 566116 313770 566126 313804
rect 509393 313610 566126 313770
rect 566346 313770 566356 313804
rect 580748 313770 580954 313775
rect 566346 313610 580758 313770
rect 509393 313602 580758 313610
rect 580944 313727 583738 313770
rect 580944 313602 583873 313727
rect 509393 313593 583873 313602
rect 559642 311744 559870 311749
rect 559642 311536 559652 311744
rect 559860 311536 559870 311744
rect 559642 311531 559870 311536
rect 573482 311700 573844 311705
rect 573482 311420 573492 311700
rect 573834 311420 573844 311700
rect 573482 311415 573844 311420
<< via3 >>
rect 510704 689882 515202 697378
rect 520704 689858 525202 697354
rect 567306 640080 573722 644324
rect 567306 630012 573722 634256
rect 559802 492324 560012 492536
rect 573564 491888 573874 492160
rect 491196 414026 491260 414030
rect 491196 413970 491200 414026
rect 491200 413970 491256 414026
rect 491256 413970 491260 414026
rect 491196 413966 491260 413970
rect 491196 413946 491260 413950
rect 491196 413890 491200 413946
rect 491200 413890 491256 413946
rect 491256 413890 491260 413946
rect 491196 413886 491260 413890
rect 491196 413866 491260 413870
rect 491196 413810 491200 413866
rect 491200 413810 491256 413866
rect 491256 413810 491260 413866
rect 491196 413806 491260 413810
rect 491196 413786 491260 413790
rect 491196 413730 491200 413786
rect 491200 413730 491256 413786
rect 491256 413730 491260 413786
rect 491196 413726 491260 413730
rect 491196 413706 491260 413710
rect 491196 413650 491200 413706
rect 491200 413650 491256 413706
rect 491256 413650 491260 413706
rect 491196 413646 491260 413650
rect 491196 413626 491260 413630
rect 491196 413570 491200 413626
rect 491200 413570 491256 413626
rect 491256 413570 491260 413626
rect 491196 413566 491260 413570
rect 491196 413546 491260 413550
rect 491196 413490 491200 413546
rect 491200 413490 491256 413546
rect 491256 413490 491260 413546
rect 491196 413486 491260 413490
rect 491196 413466 491260 413470
rect 491196 413410 491200 413466
rect 491200 413410 491256 413466
rect 491256 413410 491260 413466
rect 491196 413406 491260 413410
rect 491196 413386 491260 413390
rect 491196 413330 491200 413386
rect 491200 413330 491256 413386
rect 491256 413330 491260 413386
rect 491196 413326 491260 413330
rect 491196 413306 491260 413310
rect 491196 413250 491200 413306
rect 491200 413250 491256 413306
rect 491256 413250 491260 413306
rect 491196 413246 491260 413250
rect 491196 413226 491260 413230
rect 491196 413170 491200 413226
rect 491200 413170 491256 413226
rect 491256 413170 491260 413226
rect 491196 413166 491260 413170
rect 491196 413146 491260 413150
rect 491196 413090 491200 413146
rect 491200 413090 491256 413146
rect 491256 413090 491260 413146
rect 491196 413086 491260 413090
rect 491196 413066 491260 413070
rect 491196 413010 491200 413066
rect 491200 413010 491256 413066
rect 491256 413010 491260 413066
rect 491196 413006 491260 413010
rect 491196 412986 491260 412990
rect 491196 412930 491200 412986
rect 491200 412930 491256 412986
rect 491256 412930 491260 412986
rect 491196 412926 491260 412930
rect 491196 412906 491260 412910
rect 491196 412850 491200 412906
rect 491200 412850 491256 412906
rect 491256 412850 491260 412906
rect 491196 412846 491260 412850
rect 491196 412826 491260 412830
rect 491196 412770 491200 412826
rect 491200 412770 491256 412826
rect 491256 412770 491260 412826
rect 491196 412766 491260 412770
rect 491196 412746 491260 412750
rect 491196 412690 491200 412746
rect 491200 412690 491256 412746
rect 491256 412690 491260 412746
rect 491196 412686 491260 412690
rect 491196 412666 491260 412670
rect 491196 412610 491200 412666
rect 491200 412610 491256 412666
rect 491256 412610 491260 412666
rect 491196 412606 491260 412610
rect 491196 412586 491260 412590
rect 491196 412530 491200 412586
rect 491200 412530 491256 412586
rect 491256 412530 491260 412586
rect 491196 412526 491260 412530
rect 491196 412506 491260 412510
rect 491196 412450 491200 412506
rect 491200 412450 491256 412506
rect 491256 412450 491260 412506
rect 491196 412446 491260 412450
rect 494956 414026 495020 414030
rect 494956 413970 494960 414026
rect 494960 413970 495016 414026
rect 495016 413970 495020 414026
rect 494956 413966 495020 413970
rect 494956 413946 495020 413950
rect 494956 413890 494960 413946
rect 494960 413890 495016 413946
rect 495016 413890 495020 413946
rect 494956 413886 495020 413890
rect 494956 413866 495020 413870
rect 494956 413810 494960 413866
rect 494960 413810 495016 413866
rect 495016 413810 495020 413866
rect 494956 413806 495020 413810
rect 494956 413786 495020 413790
rect 494956 413730 494960 413786
rect 494960 413730 495016 413786
rect 495016 413730 495020 413786
rect 494956 413726 495020 413730
rect 494956 413706 495020 413710
rect 494956 413650 494960 413706
rect 494960 413650 495016 413706
rect 495016 413650 495020 413706
rect 494956 413646 495020 413650
rect 494956 413626 495020 413630
rect 494956 413570 494960 413626
rect 494960 413570 495016 413626
rect 495016 413570 495020 413626
rect 494956 413566 495020 413570
rect 494956 413546 495020 413550
rect 494956 413490 494960 413546
rect 494960 413490 495016 413546
rect 495016 413490 495020 413546
rect 494956 413486 495020 413490
rect 494956 413466 495020 413470
rect 494956 413410 494960 413466
rect 494960 413410 495016 413466
rect 495016 413410 495020 413466
rect 494956 413406 495020 413410
rect 494956 413386 495020 413390
rect 494956 413330 494960 413386
rect 494960 413330 495016 413386
rect 495016 413330 495020 413386
rect 494956 413326 495020 413330
rect 494956 413306 495020 413310
rect 494956 413250 494960 413306
rect 494960 413250 495016 413306
rect 495016 413250 495020 413306
rect 494956 413246 495020 413250
rect 494956 413226 495020 413230
rect 494956 413170 494960 413226
rect 494960 413170 495016 413226
rect 495016 413170 495020 413226
rect 494956 413166 495020 413170
rect 494956 413146 495020 413150
rect 494956 413090 494960 413146
rect 494960 413090 495016 413146
rect 495016 413090 495020 413146
rect 494956 413086 495020 413090
rect 494956 413066 495020 413070
rect 494956 413010 494960 413066
rect 494960 413010 495016 413066
rect 495016 413010 495020 413066
rect 494956 413006 495020 413010
rect 494956 412986 495020 412990
rect 494956 412930 494960 412986
rect 494960 412930 495016 412986
rect 495016 412930 495020 412986
rect 494956 412926 495020 412930
rect 494956 412906 495020 412910
rect 494956 412850 494960 412906
rect 494960 412850 495016 412906
rect 495016 412850 495020 412906
rect 494956 412846 495020 412850
rect 494956 412826 495020 412830
rect 494956 412770 494960 412826
rect 494960 412770 495016 412826
rect 495016 412770 495020 412826
rect 494956 412766 495020 412770
rect 494956 412746 495020 412750
rect 494956 412690 494960 412746
rect 494960 412690 495016 412746
rect 495016 412690 495020 412746
rect 494956 412686 495020 412690
rect 494956 412666 495020 412670
rect 494956 412610 494960 412666
rect 494960 412610 495016 412666
rect 495016 412610 495020 412666
rect 494956 412606 495020 412610
rect 494956 412586 495020 412590
rect 494956 412530 494960 412586
rect 494960 412530 495016 412586
rect 495016 412530 495020 412586
rect 494956 412526 495020 412530
rect 494956 412506 495020 412510
rect 494956 412450 494960 412506
rect 494960 412450 495016 412506
rect 495016 412450 495020 412506
rect 494956 412446 495020 412450
rect 498716 414026 498780 414030
rect 498716 413970 498720 414026
rect 498720 413970 498776 414026
rect 498776 413970 498780 414026
rect 498716 413966 498780 413970
rect 498716 413946 498780 413950
rect 498716 413890 498720 413946
rect 498720 413890 498776 413946
rect 498776 413890 498780 413946
rect 498716 413886 498780 413890
rect 498716 413866 498780 413870
rect 498716 413810 498720 413866
rect 498720 413810 498776 413866
rect 498776 413810 498780 413866
rect 498716 413806 498780 413810
rect 498716 413786 498780 413790
rect 498716 413730 498720 413786
rect 498720 413730 498776 413786
rect 498776 413730 498780 413786
rect 498716 413726 498780 413730
rect 498716 413706 498780 413710
rect 498716 413650 498720 413706
rect 498720 413650 498776 413706
rect 498776 413650 498780 413706
rect 498716 413646 498780 413650
rect 498716 413626 498780 413630
rect 498716 413570 498720 413626
rect 498720 413570 498776 413626
rect 498776 413570 498780 413626
rect 498716 413566 498780 413570
rect 498716 413546 498780 413550
rect 498716 413490 498720 413546
rect 498720 413490 498776 413546
rect 498776 413490 498780 413546
rect 498716 413486 498780 413490
rect 498716 413466 498780 413470
rect 498716 413410 498720 413466
rect 498720 413410 498776 413466
rect 498776 413410 498780 413466
rect 498716 413406 498780 413410
rect 498716 413386 498780 413390
rect 498716 413330 498720 413386
rect 498720 413330 498776 413386
rect 498776 413330 498780 413386
rect 498716 413326 498780 413330
rect 498716 413306 498780 413310
rect 498716 413250 498720 413306
rect 498720 413250 498776 413306
rect 498776 413250 498780 413306
rect 498716 413246 498780 413250
rect 498716 413226 498780 413230
rect 498716 413170 498720 413226
rect 498720 413170 498776 413226
rect 498776 413170 498780 413226
rect 498716 413166 498780 413170
rect 498716 413146 498780 413150
rect 498716 413090 498720 413146
rect 498720 413090 498776 413146
rect 498776 413090 498780 413146
rect 498716 413086 498780 413090
rect 498716 413066 498780 413070
rect 498716 413010 498720 413066
rect 498720 413010 498776 413066
rect 498776 413010 498780 413066
rect 498716 413006 498780 413010
rect 498716 412986 498780 412990
rect 498716 412930 498720 412986
rect 498720 412930 498776 412986
rect 498776 412930 498780 412986
rect 498716 412926 498780 412930
rect 498716 412906 498780 412910
rect 498716 412850 498720 412906
rect 498720 412850 498776 412906
rect 498776 412850 498780 412906
rect 498716 412846 498780 412850
rect 498716 412826 498780 412830
rect 498716 412770 498720 412826
rect 498720 412770 498776 412826
rect 498776 412770 498780 412826
rect 498716 412766 498780 412770
rect 498716 412746 498780 412750
rect 498716 412690 498720 412746
rect 498720 412690 498776 412746
rect 498776 412690 498780 412746
rect 498716 412686 498780 412690
rect 498716 412666 498780 412670
rect 498716 412610 498720 412666
rect 498720 412610 498776 412666
rect 498776 412610 498780 412666
rect 498716 412606 498780 412610
rect 498716 412586 498780 412590
rect 498716 412530 498720 412586
rect 498720 412530 498776 412586
rect 498776 412530 498780 412586
rect 498716 412526 498780 412530
rect 498716 412506 498780 412510
rect 498716 412450 498720 412506
rect 498720 412450 498776 412506
rect 498776 412450 498780 412506
rect 498716 412446 498780 412450
rect 493076 411578 493140 411582
rect 493076 411522 493080 411578
rect 493080 411522 493136 411578
rect 493136 411522 493140 411578
rect 493076 411518 493140 411522
rect 493076 411498 493140 411502
rect 493076 411442 493080 411498
rect 493080 411442 493136 411498
rect 493136 411442 493140 411498
rect 493076 411438 493140 411442
rect 493076 411418 493140 411422
rect 493076 411362 493080 411418
rect 493080 411362 493136 411418
rect 493136 411362 493140 411418
rect 493076 411358 493140 411362
rect 493076 411338 493140 411342
rect 493076 411282 493080 411338
rect 493080 411282 493136 411338
rect 493136 411282 493140 411338
rect 493076 411278 493140 411282
rect 493076 411258 493140 411262
rect 493076 411202 493080 411258
rect 493080 411202 493136 411258
rect 493136 411202 493140 411258
rect 493076 411198 493140 411202
rect 493076 411178 493140 411182
rect 493076 411122 493080 411178
rect 493080 411122 493136 411178
rect 493136 411122 493140 411178
rect 493076 411118 493140 411122
rect 493076 411098 493140 411102
rect 493076 411042 493080 411098
rect 493080 411042 493136 411098
rect 493136 411042 493140 411098
rect 493076 411038 493140 411042
rect 493076 411018 493140 411022
rect 493076 410962 493080 411018
rect 493080 410962 493136 411018
rect 493136 410962 493140 411018
rect 493076 410958 493140 410962
rect 493076 410938 493140 410942
rect 493076 410882 493080 410938
rect 493080 410882 493136 410938
rect 493136 410882 493140 410938
rect 493076 410878 493140 410882
rect 493076 410858 493140 410862
rect 493076 410802 493080 410858
rect 493080 410802 493136 410858
rect 493136 410802 493140 410858
rect 493076 410798 493140 410802
rect 493076 410778 493140 410782
rect 493076 410722 493080 410778
rect 493080 410722 493136 410778
rect 493136 410722 493140 410778
rect 493076 410718 493140 410722
rect 493076 410698 493140 410702
rect 493076 410642 493080 410698
rect 493080 410642 493136 410698
rect 493136 410642 493140 410698
rect 493076 410638 493140 410642
rect 493076 410618 493140 410622
rect 493076 410562 493080 410618
rect 493080 410562 493136 410618
rect 493136 410562 493140 410618
rect 493076 410558 493140 410562
rect 493076 410538 493140 410542
rect 493076 410482 493080 410538
rect 493080 410482 493136 410538
rect 493136 410482 493140 410538
rect 493076 410478 493140 410482
rect 493076 410458 493140 410462
rect 493076 410402 493080 410458
rect 493080 410402 493136 410458
rect 493136 410402 493140 410458
rect 493076 410398 493140 410402
rect 493076 410378 493140 410382
rect 493076 410322 493080 410378
rect 493080 410322 493136 410378
rect 493136 410322 493140 410378
rect 493076 410318 493140 410322
rect 493076 410298 493140 410302
rect 493076 410242 493080 410298
rect 493080 410242 493136 410298
rect 493136 410242 493140 410298
rect 493076 410238 493140 410242
rect 493076 410218 493140 410222
rect 493076 410162 493080 410218
rect 493080 410162 493136 410218
rect 493136 410162 493140 410218
rect 493076 410158 493140 410162
rect 493076 410138 493140 410142
rect 493076 410082 493080 410138
rect 493080 410082 493136 410138
rect 493136 410082 493140 410138
rect 493076 410078 493140 410082
rect 493076 410058 493140 410062
rect 493076 410002 493080 410058
rect 493080 410002 493136 410058
rect 493136 410002 493140 410058
rect 493076 409998 493140 410002
rect 496836 411578 496900 411582
rect 496836 411522 496840 411578
rect 496840 411522 496896 411578
rect 496896 411522 496900 411578
rect 496836 411518 496900 411522
rect 496836 411498 496900 411502
rect 496836 411442 496840 411498
rect 496840 411442 496896 411498
rect 496896 411442 496900 411498
rect 496836 411438 496900 411442
rect 496836 411418 496900 411422
rect 496836 411362 496840 411418
rect 496840 411362 496896 411418
rect 496896 411362 496900 411418
rect 496836 411358 496900 411362
rect 496836 411338 496900 411342
rect 496836 411282 496840 411338
rect 496840 411282 496896 411338
rect 496896 411282 496900 411338
rect 496836 411278 496900 411282
rect 496836 411258 496900 411262
rect 496836 411202 496840 411258
rect 496840 411202 496896 411258
rect 496896 411202 496900 411258
rect 496836 411198 496900 411202
rect 496836 411178 496900 411182
rect 496836 411122 496840 411178
rect 496840 411122 496896 411178
rect 496896 411122 496900 411178
rect 496836 411118 496900 411122
rect 496836 411098 496900 411102
rect 496836 411042 496840 411098
rect 496840 411042 496896 411098
rect 496896 411042 496900 411098
rect 496836 411038 496900 411042
rect 496836 411018 496900 411022
rect 496836 410962 496840 411018
rect 496840 410962 496896 411018
rect 496896 410962 496900 411018
rect 496836 410958 496900 410962
rect 496836 410938 496900 410942
rect 496836 410882 496840 410938
rect 496840 410882 496896 410938
rect 496896 410882 496900 410938
rect 496836 410878 496900 410882
rect 496836 410858 496900 410862
rect 496836 410802 496840 410858
rect 496840 410802 496896 410858
rect 496896 410802 496900 410858
rect 496836 410798 496900 410802
rect 496836 410778 496900 410782
rect 496836 410722 496840 410778
rect 496840 410722 496896 410778
rect 496896 410722 496900 410778
rect 496836 410718 496900 410722
rect 496836 410698 496900 410702
rect 496836 410642 496840 410698
rect 496840 410642 496896 410698
rect 496896 410642 496900 410698
rect 496836 410638 496900 410642
rect 496836 410618 496900 410622
rect 496836 410562 496840 410618
rect 496840 410562 496896 410618
rect 496896 410562 496900 410618
rect 496836 410558 496900 410562
rect 496836 410538 496900 410542
rect 496836 410482 496840 410538
rect 496840 410482 496896 410538
rect 496896 410482 496900 410538
rect 496836 410478 496900 410482
rect 496836 410458 496900 410462
rect 496836 410402 496840 410458
rect 496840 410402 496896 410458
rect 496896 410402 496900 410458
rect 496836 410398 496900 410402
rect 496836 410378 496900 410382
rect 496836 410322 496840 410378
rect 496840 410322 496896 410378
rect 496896 410322 496900 410378
rect 496836 410318 496900 410322
rect 496836 410298 496900 410302
rect 496836 410242 496840 410298
rect 496840 410242 496896 410298
rect 496896 410242 496900 410298
rect 496836 410238 496900 410242
rect 496836 410218 496900 410222
rect 496836 410162 496840 410218
rect 496840 410162 496896 410218
rect 496896 410162 496900 410218
rect 496836 410158 496900 410162
rect 496836 410138 496900 410142
rect 496836 410082 496840 410138
rect 496840 410082 496896 410138
rect 496896 410082 496900 410138
rect 496836 410078 496900 410082
rect 496836 410058 496900 410062
rect 496836 410002 496840 410058
rect 496840 410002 496896 410058
rect 496896 410002 496900 410058
rect 496836 409998 496900 410002
rect 500596 411578 500660 411582
rect 500596 411522 500600 411578
rect 500600 411522 500656 411578
rect 500656 411522 500660 411578
rect 500596 411518 500660 411522
rect 500596 411498 500660 411502
rect 500596 411442 500600 411498
rect 500600 411442 500656 411498
rect 500656 411442 500660 411498
rect 500596 411438 500660 411442
rect 500596 411418 500660 411422
rect 500596 411362 500600 411418
rect 500600 411362 500656 411418
rect 500656 411362 500660 411418
rect 500596 411358 500660 411362
rect 500596 411338 500660 411342
rect 500596 411282 500600 411338
rect 500600 411282 500656 411338
rect 500656 411282 500660 411338
rect 500596 411278 500660 411282
rect 500596 411258 500660 411262
rect 500596 411202 500600 411258
rect 500600 411202 500656 411258
rect 500656 411202 500660 411258
rect 500596 411198 500660 411202
rect 500596 411178 500660 411182
rect 500596 411122 500600 411178
rect 500600 411122 500656 411178
rect 500656 411122 500660 411178
rect 500596 411118 500660 411122
rect 500596 411098 500660 411102
rect 500596 411042 500600 411098
rect 500600 411042 500656 411098
rect 500656 411042 500660 411098
rect 500596 411038 500660 411042
rect 500596 411018 500660 411022
rect 500596 410962 500600 411018
rect 500600 410962 500656 411018
rect 500656 410962 500660 411018
rect 500596 410958 500660 410962
rect 500596 410938 500660 410942
rect 500596 410882 500600 410938
rect 500600 410882 500656 410938
rect 500656 410882 500660 410938
rect 500596 410878 500660 410882
rect 500596 410858 500660 410862
rect 500596 410802 500600 410858
rect 500600 410802 500656 410858
rect 500656 410802 500660 410858
rect 500596 410798 500660 410802
rect 500596 410778 500660 410782
rect 500596 410722 500600 410778
rect 500600 410722 500656 410778
rect 500656 410722 500660 410778
rect 500596 410718 500660 410722
rect 500596 410698 500660 410702
rect 500596 410642 500600 410698
rect 500600 410642 500656 410698
rect 500656 410642 500660 410698
rect 500596 410638 500660 410642
rect 500596 410618 500660 410622
rect 500596 410562 500600 410618
rect 500600 410562 500656 410618
rect 500656 410562 500660 410618
rect 500596 410558 500660 410562
rect 500596 410538 500660 410542
rect 500596 410482 500600 410538
rect 500600 410482 500656 410538
rect 500656 410482 500660 410538
rect 500596 410478 500660 410482
rect 500596 410458 500660 410462
rect 500596 410402 500600 410458
rect 500600 410402 500656 410458
rect 500656 410402 500660 410458
rect 500596 410398 500660 410402
rect 500596 410378 500660 410382
rect 500596 410322 500600 410378
rect 500600 410322 500656 410378
rect 500656 410322 500660 410378
rect 500596 410318 500660 410322
rect 500596 410298 500660 410302
rect 500596 410242 500600 410298
rect 500600 410242 500656 410298
rect 500656 410242 500660 410298
rect 500596 410238 500660 410242
rect 500596 410218 500660 410222
rect 500596 410162 500600 410218
rect 500600 410162 500656 410218
rect 500656 410162 500660 410218
rect 500596 410158 500660 410162
rect 500596 410138 500660 410142
rect 500596 410082 500600 410138
rect 500600 410082 500656 410138
rect 500656 410082 500660 410138
rect 500596 410078 500660 410082
rect 500596 410058 500660 410062
rect 500596 410002 500600 410058
rect 500600 410002 500656 410058
rect 500656 410002 500660 410058
rect 500596 409998 500660 410002
rect 502476 414026 502540 414030
rect 502476 413970 502480 414026
rect 502480 413970 502536 414026
rect 502536 413970 502540 414026
rect 502476 413966 502540 413970
rect 502476 413946 502540 413950
rect 502476 413890 502480 413946
rect 502480 413890 502536 413946
rect 502536 413890 502540 413946
rect 502476 413886 502540 413890
rect 502476 413866 502540 413870
rect 502476 413810 502480 413866
rect 502480 413810 502536 413866
rect 502536 413810 502540 413866
rect 502476 413806 502540 413810
rect 502476 413786 502540 413790
rect 502476 413730 502480 413786
rect 502480 413730 502536 413786
rect 502536 413730 502540 413786
rect 502476 413726 502540 413730
rect 502476 413706 502540 413710
rect 502476 413650 502480 413706
rect 502480 413650 502536 413706
rect 502536 413650 502540 413706
rect 502476 413646 502540 413650
rect 502476 413626 502540 413630
rect 502476 413570 502480 413626
rect 502480 413570 502536 413626
rect 502536 413570 502540 413626
rect 502476 413566 502540 413570
rect 502476 413546 502540 413550
rect 502476 413490 502480 413546
rect 502480 413490 502536 413546
rect 502536 413490 502540 413546
rect 502476 413486 502540 413490
rect 502476 413466 502540 413470
rect 502476 413410 502480 413466
rect 502480 413410 502536 413466
rect 502536 413410 502540 413466
rect 502476 413406 502540 413410
rect 502476 413386 502540 413390
rect 502476 413330 502480 413386
rect 502480 413330 502536 413386
rect 502536 413330 502540 413386
rect 502476 413326 502540 413330
rect 502476 413306 502540 413310
rect 502476 413250 502480 413306
rect 502480 413250 502536 413306
rect 502536 413250 502540 413306
rect 502476 413246 502540 413250
rect 502476 413226 502540 413230
rect 502476 413170 502480 413226
rect 502480 413170 502536 413226
rect 502536 413170 502540 413226
rect 502476 413166 502540 413170
rect 502476 413146 502540 413150
rect 502476 413090 502480 413146
rect 502480 413090 502536 413146
rect 502536 413090 502540 413146
rect 502476 413086 502540 413090
rect 502476 413066 502540 413070
rect 502476 413010 502480 413066
rect 502480 413010 502536 413066
rect 502536 413010 502540 413066
rect 502476 413006 502540 413010
rect 502476 412986 502540 412990
rect 502476 412930 502480 412986
rect 502480 412930 502536 412986
rect 502536 412930 502540 412986
rect 502476 412926 502540 412930
rect 502476 412906 502540 412910
rect 502476 412850 502480 412906
rect 502480 412850 502536 412906
rect 502536 412850 502540 412906
rect 502476 412846 502540 412850
rect 502476 412826 502540 412830
rect 502476 412770 502480 412826
rect 502480 412770 502536 412826
rect 502536 412770 502540 412826
rect 502476 412766 502540 412770
rect 502476 412746 502540 412750
rect 502476 412690 502480 412746
rect 502480 412690 502536 412746
rect 502536 412690 502540 412746
rect 502476 412686 502540 412690
rect 502476 412666 502540 412670
rect 502476 412610 502480 412666
rect 502480 412610 502536 412666
rect 502536 412610 502540 412666
rect 502476 412606 502540 412610
rect 502476 412586 502540 412590
rect 502476 412530 502480 412586
rect 502480 412530 502536 412586
rect 502536 412530 502540 412586
rect 502476 412526 502540 412530
rect 502476 412506 502540 412510
rect 502476 412450 502480 412506
rect 502480 412450 502536 412506
rect 502536 412450 502540 412506
rect 502476 412446 502540 412450
rect 506236 414026 506300 414030
rect 506236 413970 506240 414026
rect 506240 413970 506296 414026
rect 506296 413970 506300 414026
rect 506236 413966 506300 413970
rect 506236 413946 506300 413950
rect 506236 413890 506240 413946
rect 506240 413890 506296 413946
rect 506296 413890 506300 413946
rect 506236 413886 506300 413890
rect 506236 413866 506300 413870
rect 506236 413810 506240 413866
rect 506240 413810 506296 413866
rect 506296 413810 506300 413866
rect 506236 413806 506300 413810
rect 506236 413786 506300 413790
rect 506236 413730 506240 413786
rect 506240 413730 506296 413786
rect 506296 413730 506300 413786
rect 506236 413726 506300 413730
rect 506236 413706 506300 413710
rect 506236 413650 506240 413706
rect 506240 413650 506296 413706
rect 506296 413650 506300 413706
rect 506236 413646 506300 413650
rect 506236 413626 506300 413630
rect 506236 413570 506240 413626
rect 506240 413570 506296 413626
rect 506296 413570 506300 413626
rect 506236 413566 506300 413570
rect 506236 413546 506300 413550
rect 506236 413490 506240 413546
rect 506240 413490 506296 413546
rect 506296 413490 506300 413546
rect 506236 413486 506300 413490
rect 506236 413466 506300 413470
rect 506236 413410 506240 413466
rect 506240 413410 506296 413466
rect 506296 413410 506300 413466
rect 506236 413406 506300 413410
rect 506236 413386 506300 413390
rect 506236 413330 506240 413386
rect 506240 413330 506296 413386
rect 506296 413330 506300 413386
rect 506236 413326 506300 413330
rect 506236 413306 506300 413310
rect 506236 413250 506240 413306
rect 506240 413250 506296 413306
rect 506296 413250 506300 413306
rect 506236 413246 506300 413250
rect 506236 413226 506300 413230
rect 506236 413170 506240 413226
rect 506240 413170 506296 413226
rect 506296 413170 506300 413226
rect 506236 413166 506300 413170
rect 506236 413146 506300 413150
rect 506236 413090 506240 413146
rect 506240 413090 506296 413146
rect 506296 413090 506300 413146
rect 506236 413086 506300 413090
rect 506236 413066 506300 413070
rect 506236 413010 506240 413066
rect 506240 413010 506296 413066
rect 506296 413010 506300 413066
rect 506236 413006 506300 413010
rect 506236 412986 506300 412990
rect 506236 412930 506240 412986
rect 506240 412930 506296 412986
rect 506296 412930 506300 412986
rect 506236 412926 506300 412930
rect 506236 412906 506300 412910
rect 506236 412850 506240 412906
rect 506240 412850 506296 412906
rect 506296 412850 506300 412906
rect 506236 412846 506300 412850
rect 506236 412826 506300 412830
rect 506236 412770 506240 412826
rect 506240 412770 506296 412826
rect 506296 412770 506300 412826
rect 506236 412766 506300 412770
rect 506236 412746 506300 412750
rect 506236 412690 506240 412746
rect 506240 412690 506296 412746
rect 506296 412690 506300 412746
rect 506236 412686 506300 412690
rect 506236 412666 506300 412670
rect 506236 412610 506240 412666
rect 506240 412610 506296 412666
rect 506296 412610 506300 412666
rect 506236 412606 506300 412610
rect 506236 412586 506300 412590
rect 506236 412530 506240 412586
rect 506240 412530 506296 412586
rect 506296 412530 506300 412586
rect 506236 412526 506300 412530
rect 506236 412506 506300 412510
rect 506236 412450 506240 412506
rect 506240 412450 506296 412506
rect 506296 412450 506300 412506
rect 506236 412446 506300 412450
rect 509996 414026 510060 414030
rect 509996 413970 510000 414026
rect 510000 413970 510056 414026
rect 510056 413970 510060 414026
rect 509996 413966 510060 413970
rect 509996 413946 510060 413950
rect 509996 413890 510000 413946
rect 510000 413890 510056 413946
rect 510056 413890 510060 413946
rect 509996 413886 510060 413890
rect 509996 413866 510060 413870
rect 509996 413810 510000 413866
rect 510000 413810 510056 413866
rect 510056 413810 510060 413866
rect 509996 413806 510060 413810
rect 509996 413786 510060 413790
rect 509996 413730 510000 413786
rect 510000 413730 510056 413786
rect 510056 413730 510060 413786
rect 509996 413726 510060 413730
rect 509996 413706 510060 413710
rect 509996 413650 510000 413706
rect 510000 413650 510056 413706
rect 510056 413650 510060 413706
rect 509996 413646 510060 413650
rect 509996 413626 510060 413630
rect 509996 413570 510000 413626
rect 510000 413570 510056 413626
rect 510056 413570 510060 413626
rect 509996 413566 510060 413570
rect 509996 413546 510060 413550
rect 509996 413490 510000 413546
rect 510000 413490 510056 413546
rect 510056 413490 510060 413546
rect 509996 413486 510060 413490
rect 509996 413466 510060 413470
rect 509996 413410 510000 413466
rect 510000 413410 510056 413466
rect 510056 413410 510060 413466
rect 509996 413406 510060 413410
rect 509996 413386 510060 413390
rect 509996 413330 510000 413386
rect 510000 413330 510056 413386
rect 510056 413330 510060 413386
rect 509996 413326 510060 413330
rect 509996 413306 510060 413310
rect 509996 413250 510000 413306
rect 510000 413250 510056 413306
rect 510056 413250 510060 413306
rect 509996 413246 510060 413250
rect 509996 413226 510060 413230
rect 509996 413170 510000 413226
rect 510000 413170 510056 413226
rect 510056 413170 510060 413226
rect 509996 413166 510060 413170
rect 509996 413146 510060 413150
rect 509996 413090 510000 413146
rect 510000 413090 510056 413146
rect 510056 413090 510060 413146
rect 509996 413086 510060 413090
rect 509996 413066 510060 413070
rect 509996 413010 510000 413066
rect 510000 413010 510056 413066
rect 510056 413010 510060 413066
rect 509996 413006 510060 413010
rect 509996 412986 510060 412990
rect 509996 412930 510000 412986
rect 510000 412930 510056 412986
rect 510056 412930 510060 412986
rect 509996 412926 510060 412930
rect 509996 412906 510060 412910
rect 509996 412850 510000 412906
rect 510000 412850 510056 412906
rect 510056 412850 510060 412906
rect 509996 412846 510060 412850
rect 509996 412826 510060 412830
rect 509996 412770 510000 412826
rect 510000 412770 510056 412826
rect 510056 412770 510060 412826
rect 509996 412766 510060 412770
rect 509996 412746 510060 412750
rect 509996 412690 510000 412746
rect 510000 412690 510056 412746
rect 510056 412690 510060 412746
rect 509996 412686 510060 412690
rect 509996 412666 510060 412670
rect 509996 412610 510000 412666
rect 510000 412610 510056 412666
rect 510056 412610 510060 412666
rect 509996 412606 510060 412610
rect 509996 412586 510060 412590
rect 509996 412530 510000 412586
rect 510000 412530 510056 412586
rect 510056 412530 510060 412586
rect 509996 412526 510060 412530
rect 509996 412506 510060 412510
rect 509996 412450 510000 412506
rect 510000 412450 510056 412506
rect 510056 412450 510060 412506
rect 509996 412446 510060 412450
rect 513756 414026 513820 414030
rect 513756 413970 513760 414026
rect 513760 413970 513816 414026
rect 513816 413970 513820 414026
rect 513756 413966 513820 413970
rect 513756 413946 513820 413950
rect 513756 413890 513760 413946
rect 513760 413890 513816 413946
rect 513816 413890 513820 413946
rect 513756 413886 513820 413890
rect 513756 413866 513820 413870
rect 513756 413810 513760 413866
rect 513760 413810 513816 413866
rect 513816 413810 513820 413866
rect 513756 413806 513820 413810
rect 513756 413786 513820 413790
rect 513756 413730 513760 413786
rect 513760 413730 513816 413786
rect 513816 413730 513820 413786
rect 513756 413726 513820 413730
rect 513756 413706 513820 413710
rect 513756 413650 513760 413706
rect 513760 413650 513816 413706
rect 513816 413650 513820 413706
rect 513756 413646 513820 413650
rect 513756 413626 513820 413630
rect 513756 413570 513760 413626
rect 513760 413570 513816 413626
rect 513816 413570 513820 413626
rect 513756 413566 513820 413570
rect 513756 413546 513820 413550
rect 513756 413490 513760 413546
rect 513760 413490 513816 413546
rect 513816 413490 513820 413546
rect 513756 413486 513820 413490
rect 513756 413466 513820 413470
rect 513756 413410 513760 413466
rect 513760 413410 513816 413466
rect 513816 413410 513820 413466
rect 513756 413406 513820 413410
rect 513756 413386 513820 413390
rect 513756 413330 513760 413386
rect 513760 413330 513816 413386
rect 513816 413330 513820 413386
rect 513756 413326 513820 413330
rect 513756 413306 513820 413310
rect 513756 413250 513760 413306
rect 513760 413250 513816 413306
rect 513816 413250 513820 413306
rect 513756 413246 513820 413250
rect 513756 413226 513820 413230
rect 513756 413170 513760 413226
rect 513760 413170 513816 413226
rect 513816 413170 513820 413226
rect 513756 413166 513820 413170
rect 513756 413146 513820 413150
rect 513756 413090 513760 413146
rect 513760 413090 513816 413146
rect 513816 413090 513820 413146
rect 513756 413086 513820 413090
rect 513756 413066 513820 413070
rect 513756 413010 513760 413066
rect 513760 413010 513816 413066
rect 513816 413010 513820 413066
rect 513756 413006 513820 413010
rect 513756 412986 513820 412990
rect 513756 412930 513760 412986
rect 513760 412930 513816 412986
rect 513816 412930 513820 412986
rect 513756 412926 513820 412930
rect 513756 412906 513820 412910
rect 513756 412850 513760 412906
rect 513760 412850 513816 412906
rect 513816 412850 513820 412906
rect 513756 412846 513820 412850
rect 513756 412826 513820 412830
rect 513756 412770 513760 412826
rect 513760 412770 513816 412826
rect 513816 412770 513820 412826
rect 513756 412766 513820 412770
rect 513756 412746 513820 412750
rect 513756 412690 513760 412746
rect 513760 412690 513816 412746
rect 513816 412690 513820 412746
rect 513756 412686 513820 412690
rect 513756 412666 513820 412670
rect 513756 412610 513760 412666
rect 513760 412610 513816 412666
rect 513816 412610 513820 412666
rect 513756 412606 513820 412610
rect 513756 412586 513820 412590
rect 513756 412530 513760 412586
rect 513760 412530 513816 412586
rect 513816 412530 513820 412586
rect 513756 412526 513820 412530
rect 513756 412506 513820 412510
rect 513756 412450 513760 412506
rect 513760 412450 513816 412506
rect 513816 412450 513820 412506
rect 513756 412446 513820 412450
rect 517516 414026 517580 414030
rect 517516 413970 517520 414026
rect 517520 413970 517576 414026
rect 517576 413970 517580 414026
rect 517516 413966 517580 413970
rect 517516 413946 517580 413950
rect 517516 413890 517520 413946
rect 517520 413890 517576 413946
rect 517576 413890 517580 413946
rect 517516 413886 517580 413890
rect 517516 413866 517580 413870
rect 517516 413810 517520 413866
rect 517520 413810 517576 413866
rect 517576 413810 517580 413866
rect 517516 413806 517580 413810
rect 517516 413786 517580 413790
rect 517516 413730 517520 413786
rect 517520 413730 517576 413786
rect 517576 413730 517580 413786
rect 517516 413726 517580 413730
rect 517516 413706 517580 413710
rect 517516 413650 517520 413706
rect 517520 413650 517576 413706
rect 517576 413650 517580 413706
rect 517516 413646 517580 413650
rect 517516 413626 517580 413630
rect 517516 413570 517520 413626
rect 517520 413570 517576 413626
rect 517576 413570 517580 413626
rect 517516 413566 517580 413570
rect 517516 413546 517580 413550
rect 517516 413490 517520 413546
rect 517520 413490 517576 413546
rect 517576 413490 517580 413546
rect 517516 413486 517580 413490
rect 517516 413466 517580 413470
rect 517516 413410 517520 413466
rect 517520 413410 517576 413466
rect 517576 413410 517580 413466
rect 517516 413406 517580 413410
rect 517516 413386 517580 413390
rect 517516 413330 517520 413386
rect 517520 413330 517576 413386
rect 517576 413330 517580 413386
rect 517516 413326 517580 413330
rect 517516 413306 517580 413310
rect 517516 413250 517520 413306
rect 517520 413250 517576 413306
rect 517576 413250 517580 413306
rect 517516 413246 517580 413250
rect 517516 413226 517580 413230
rect 517516 413170 517520 413226
rect 517520 413170 517576 413226
rect 517576 413170 517580 413226
rect 517516 413166 517580 413170
rect 517516 413146 517580 413150
rect 517516 413090 517520 413146
rect 517520 413090 517576 413146
rect 517576 413090 517580 413146
rect 517516 413086 517580 413090
rect 517516 413066 517580 413070
rect 517516 413010 517520 413066
rect 517520 413010 517576 413066
rect 517576 413010 517580 413066
rect 517516 413006 517580 413010
rect 517516 412986 517580 412990
rect 517516 412930 517520 412986
rect 517520 412930 517576 412986
rect 517576 412930 517580 412986
rect 517516 412926 517580 412930
rect 517516 412906 517580 412910
rect 517516 412850 517520 412906
rect 517520 412850 517576 412906
rect 517576 412850 517580 412906
rect 517516 412846 517580 412850
rect 517516 412826 517580 412830
rect 517516 412770 517520 412826
rect 517520 412770 517576 412826
rect 517576 412770 517580 412826
rect 517516 412766 517580 412770
rect 517516 412746 517580 412750
rect 517516 412690 517520 412746
rect 517520 412690 517576 412746
rect 517576 412690 517580 412746
rect 517516 412686 517580 412690
rect 517516 412666 517580 412670
rect 517516 412610 517520 412666
rect 517520 412610 517576 412666
rect 517576 412610 517580 412666
rect 517516 412606 517580 412610
rect 517516 412586 517580 412590
rect 517516 412530 517520 412586
rect 517520 412530 517576 412586
rect 517576 412530 517580 412586
rect 517516 412526 517580 412530
rect 517516 412506 517580 412510
rect 517516 412450 517520 412506
rect 517520 412450 517576 412506
rect 517576 412450 517580 412506
rect 517516 412446 517580 412450
rect 521276 414026 521340 414030
rect 521276 413970 521280 414026
rect 521280 413970 521336 414026
rect 521336 413970 521340 414026
rect 521276 413966 521340 413970
rect 521276 413946 521340 413950
rect 521276 413890 521280 413946
rect 521280 413890 521336 413946
rect 521336 413890 521340 413946
rect 521276 413886 521340 413890
rect 521276 413866 521340 413870
rect 521276 413810 521280 413866
rect 521280 413810 521336 413866
rect 521336 413810 521340 413866
rect 521276 413806 521340 413810
rect 521276 413786 521340 413790
rect 521276 413730 521280 413786
rect 521280 413730 521336 413786
rect 521336 413730 521340 413786
rect 521276 413726 521340 413730
rect 521276 413706 521340 413710
rect 521276 413650 521280 413706
rect 521280 413650 521336 413706
rect 521336 413650 521340 413706
rect 521276 413646 521340 413650
rect 521276 413626 521340 413630
rect 521276 413570 521280 413626
rect 521280 413570 521336 413626
rect 521336 413570 521340 413626
rect 521276 413566 521340 413570
rect 521276 413546 521340 413550
rect 521276 413490 521280 413546
rect 521280 413490 521336 413546
rect 521336 413490 521340 413546
rect 521276 413486 521340 413490
rect 521276 413466 521340 413470
rect 521276 413410 521280 413466
rect 521280 413410 521336 413466
rect 521336 413410 521340 413466
rect 521276 413406 521340 413410
rect 521276 413386 521340 413390
rect 521276 413330 521280 413386
rect 521280 413330 521336 413386
rect 521336 413330 521340 413386
rect 521276 413326 521340 413330
rect 521276 413306 521340 413310
rect 521276 413250 521280 413306
rect 521280 413250 521336 413306
rect 521336 413250 521340 413306
rect 521276 413246 521340 413250
rect 521276 413226 521340 413230
rect 521276 413170 521280 413226
rect 521280 413170 521336 413226
rect 521336 413170 521340 413226
rect 521276 413166 521340 413170
rect 521276 413146 521340 413150
rect 521276 413090 521280 413146
rect 521280 413090 521336 413146
rect 521336 413090 521340 413146
rect 521276 413086 521340 413090
rect 521276 413066 521340 413070
rect 521276 413010 521280 413066
rect 521280 413010 521336 413066
rect 521336 413010 521340 413066
rect 521276 413006 521340 413010
rect 521276 412986 521340 412990
rect 521276 412930 521280 412986
rect 521280 412930 521336 412986
rect 521336 412930 521340 412986
rect 521276 412926 521340 412930
rect 521276 412906 521340 412910
rect 521276 412850 521280 412906
rect 521280 412850 521336 412906
rect 521336 412850 521340 412906
rect 521276 412846 521340 412850
rect 521276 412826 521340 412830
rect 521276 412770 521280 412826
rect 521280 412770 521336 412826
rect 521336 412770 521340 412826
rect 521276 412766 521340 412770
rect 521276 412746 521340 412750
rect 521276 412690 521280 412746
rect 521280 412690 521336 412746
rect 521336 412690 521340 412746
rect 521276 412686 521340 412690
rect 521276 412666 521340 412670
rect 521276 412610 521280 412666
rect 521280 412610 521336 412666
rect 521336 412610 521340 412666
rect 521276 412606 521340 412610
rect 521276 412586 521340 412590
rect 521276 412530 521280 412586
rect 521280 412530 521336 412586
rect 521336 412530 521340 412586
rect 521276 412526 521340 412530
rect 521276 412506 521340 412510
rect 521276 412450 521280 412506
rect 521280 412450 521336 412506
rect 521336 412450 521340 412506
rect 521276 412446 521340 412450
rect 525036 414026 525100 414030
rect 525036 413970 525040 414026
rect 525040 413970 525096 414026
rect 525096 413970 525100 414026
rect 525036 413966 525100 413970
rect 525036 413946 525100 413950
rect 525036 413890 525040 413946
rect 525040 413890 525096 413946
rect 525096 413890 525100 413946
rect 525036 413886 525100 413890
rect 525036 413866 525100 413870
rect 525036 413810 525040 413866
rect 525040 413810 525096 413866
rect 525096 413810 525100 413866
rect 525036 413806 525100 413810
rect 525036 413786 525100 413790
rect 525036 413730 525040 413786
rect 525040 413730 525096 413786
rect 525096 413730 525100 413786
rect 525036 413726 525100 413730
rect 525036 413706 525100 413710
rect 525036 413650 525040 413706
rect 525040 413650 525096 413706
rect 525096 413650 525100 413706
rect 525036 413646 525100 413650
rect 525036 413626 525100 413630
rect 525036 413570 525040 413626
rect 525040 413570 525096 413626
rect 525096 413570 525100 413626
rect 525036 413566 525100 413570
rect 525036 413546 525100 413550
rect 525036 413490 525040 413546
rect 525040 413490 525096 413546
rect 525096 413490 525100 413546
rect 525036 413486 525100 413490
rect 525036 413466 525100 413470
rect 525036 413410 525040 413466
rect 525040 413410 525096 413466
rect 525096 413410 525100 413466
rect 525036 413406 525100 413410
rect 525036 413386 525100 413390
rect 525036 413330 525040 413386
rect 525040 413330 525096 413386
rect 525096 413330 525100 413386
rect 525036 413326 525100 413330
rect 525036 413306 525100 413310
rect 525036 413250 525040 413306
rect 525040 413250 525096 413306
rect 525096 413250 525100 413306
rect 525036 413246 525100 413250
rect 525036 413226 525100 413230
rect 525036 413170 525040 413226
rect 525040 413170 525096 413226
rect 525096 413170 525100 413226
rect 525036 413166 525100 413170
rect 525036 413146 525100 413150
rect 525036 413090 525040 413146
rect 525040 413090 525096 413146
rect 525096 413090 525100 413146
rect 525036 413086 525100 413090
rect 525036 413066 525100 413070
rect 525036 413010 525040 413066
rect 525040 413010 525096 413066
rect 525096 413010 525100 413066
rect 525036 413006 525100 413010
rect 525036 412986 525100 412990
rect 525036 412930 525040 412986
rect 525040 412930 525096 412986
rect 525096 412930 525100 412986
rect 525036 412926 525100 412930
rect 525036 412906 525100 412910
rect 525036 412850 525040 412906
rect 525040 412850 525096 412906
rect 525096 412850 525100 412906
rect 525036 412846 525100 412850
rect 525036 412826 525100 412830
rect 525036 412770 525040 412826
rect 525040 412770 525096 412826
rect 525096 412770 525100 412826
rect 525036 412766 525100 412770
rect 525036 412746 525100 412750
rect 525036 412690 525040 412746
rect 525040 412690 525096 412746
rect 525096 412690 525100 412746
rect 525036 412686 525100 412690
rect 525036 412666 525100 412670
rect 525036 412610 525040 412666
rect 525040 412610 525096 412666
rect 525096 412610 525100 412666
rect 525036 412606 525100 412610
rect 525036 412586 525100 412590
rect 525036 412530 525040 412586
rect 525040 412530 525096 412586
rect 525096 412530 525100 412586
rect 525036 412526 525100 412530
rect 525036 412506 525100 412510
rect 525036 412450 525040 412506
rect 525040 412450 525096 412506
rect 525096 412450 525100 412506
rect 525036 412446 525100 412450
rect 528796 414026 528860 414030
rect 528796 413970 528800 414026
rect 528800 413970 528856 414026
rect 528856 413970 528860 414026
rect 528796 413966 528860 413970
rect 528796 413946 528860 413950
rect 528796 413890 528800 413946
rect 528800 413890 528856 413946
rect 528856 413890 528860 413946
rect 528796 413886 528860 413890
rect 528796 413866 528860 413870
rect 528796 413810 528800 413866
rect 528800 413810 528856 413866
rect 528856 413810 528860 413866
rect 528796 413806 528860 413810
rect 528796 413786 528860 413790
rect 528796 413730 528800 413786
rect 528800 413730 528856 413786
rect 528856 413730 528860 413786
rect 528796 413726 528860 413730
rect 528796 413706 528860 413710
rect 528796 413650 528800 413706
rect 528800 413650 528856 413706
rect 528856 413650 528860 413706
rect 528796 413646 528860 413650
rect 528796 413626 528860 413630
rect 528796 413570 528800 413626
rect 528800 413570 528856 413626
rect 528856 413570 528860 413626
rect 528796 413566 528860 413570
rect 528796 413546 528860 413550
rect 528796 413490 528800 413546
rect 528800 413490 528856 413546
rect 528856 413490 528860 413546
rect 528796 413486 528860 413490
rect 528796 413466 528860 413470
rect 528796 413410 528800 413466
rect 528800 413410 528856 413466
rect 528856 413410 528860 413466
rect 528796 413406 528860 413410
rect 528796 413386 528860 413390
rect 528796 413330 528800 413386
rect 528800 413330 528856 413386
rect 528856 413330 528860 413386
rect 528796 413326 528860 413330
rect 528796 413306 528860 413310
rect 528796 413250 528800 413306
rect 528800 413250 528856 413306
rect 528856 413250 528860 413306
rect 528796 413246 528860 413250
rect 528796 413226 528860 413230
rect 528796 413170 528800 413226
rect 528800 413170 528856 413226
rect 528856 413170 528860 413226
rect 528796 413166 528860 413170
rect 528796 413146 528860 413150
rect 528796 413090 528800 413146
rect 528800 413090 528856 413146
rect 528856 413090 528860 413146
rect 528796 413086 528860 413090
rect 528796 413066 528860 413070
rect 528796 413010 528800 413066
rect 528800 413010 528856 413066
rect 528856 413010 528860 413066
rect 528796 413006 528860 413010
rect 528796 412986 528860 412990
rect 528796 412930 528800 412986
rect 528800 412930 528856 412986
rect 528856 412930 528860 412986
rect 528796 412926 528860 412930
rect 528796 412906 528860 412910
rect 528796 412850 528800 412906
rect 528800 412850 528856 412906
rect 528856 412850 528860 412906
rect 528796 412846 528860 412850
rect 528796 412826 528860 412830
rect 528796 412770 528800 412826
rect 528800 412770 528856 412826
rect 528856 412770 528860 412826
rect 528796 412766 528860 412770
rect 528796 412746 528860 412750
rect 528796 412690 528800 412746
rect 528800 412690 528856 412746
rect 528856 412690 528860 412746
rect 528796 412686 528860 412690
rect 528796 412666 528860 412670
rect 528796 412610 528800 412666
rect 528800 412610 528856 412666
rect 528856 412610 528860 412666
rect 528796 412606 528860 412610
rect 528796 412586 528860 412590
rect 528796 412530 528800 412586
rect 528800 412530 528856 412586
rect 528856 412530 528860 412586
rect 528796 412526 528860 412530
rect 528796 412506 528860 412510
rect 528796 412450 528800 412506
rect 528800 412450 528856 412506
rect 528856 412450 528860 412506
rect 528796 412446 528860 412450
rect 532556 414026 532620 414030
rect 532556 413970 532560 414026
rect 532560 413970 532616 414026
rect 532616 413970 532620 414026
rect 532556 413966 532620 413970
rect 532556 413946 532620 413950
rect 532556 413890 532560 413946
rect 532560 413890 532616 413946
rect 532616 413890 532620 413946
rect 532556 413886 532620 413890
rect 532556 413866 532620 413870
rect 532556 413810 532560 413866
rect 532560 413810 532616 413866
rect 532616 413810 532620 413866
rect 532556 413806 532620 413810
rect 532556 413786 532620 413790
rect 532556 413730 532560 413786
rect 532560 413730 532616 413786
rect 532616 413730 532620 413786
rect 532556 413726 532620 413730
rect 532556 413706 532620 413710
rect 532556 413650 532560 413706
rect 532560 413650 532616 413706
rect 532616 413650 532620 413706
rect 532556 413646 532620 413650
rect 532556 413626 532620 413630
rect 532556 413570 532560 413626
rect 532560 413570 532616 413626
rect 532616 413570 532620 413626
rect 532556 413566 532620 413570
rect 532556 413546 532620 413550
rect 532556 413490 532560 413546
rect 532560 413490 532616 413546
rect 532616 413490 532620 413546
rect 532556 413486 532620 413490
rect 532556 413466 532620 413470
rect 532556 413410 532560 413466
rect 532560 413410 532616 413466
rect 532616 413410 532620 413466
rect 532556 413406 532620 413410
rect 532556 413386 532620 413390
rect 532556 413330 532560 413386
rect 532560 413330 532616 413386
rect 532616 413330 532620 413386
rect 532556 413326 532620 413330
rect 532556 413306 532620 413310
rect 532556 413250 532560 413306
rect 532560 413250 532616 413306
rect 532616 413250 532620 413306
rect 532556 413246 532620 413250
rect 532556 413226 532620 413230
rect 532556 413170 532560 413226
rect 532560 413170 532616 413226
rect 532616 413170 532620 413226
rect 532556 413166 532620 413170
rect 532556 413146 532620 413150
rect 532556 413090 532560 413146
rect 532560 413090 532616 413146
rect 532616 413090 532620 413146
rect 532556 413086 532620 413090
rect 532556 413066 532620 413070
rect 532556 413010 532560 413066
rect 532560 413010 532616 413066
rect 532616 413010 532620 413066
rect 532556 413006 532620 413010
rect 532556 412986 532620 412990
rect 532556 412930 532560 412986
rect 532560 412930 532616 412986
rect 532616 412930 532620 412986
rect 532556 412926 532620 412930
rect 532556 412906 532620 412910
rect 532556 412850 532560 412906
rect 532560 412850 532616 412906
rect 532616 412850 532620 412906
rect 532556 412846 532620 412850
rect 532556 412826 532620 412830
rect 532556 412770 532560 412826
rect 532560 412770 532616 412826
rect 532616 412770 532620 412826
rect 532556 412766 532620 412770
rect 532556 412746 532620 412750
rect 532556 412690 532560 412746
rect 532560 412690 532616 412746
rect 532616 412690 532620 412746
rect 532556 412686 532620 412690
rect 532556 412666 532620 412670
rect 532556 412610 532560 412666
rect 532560 412610 532616 412666
rect 532616 412610 532620 412666
rect 532556 412606 532620 412610
rect 532556 412586 532620 412590
rect 532556 412530 532560 412586
rect 532560 412530 532616 412586
rect 532616 412530 532620 412586
rect 532556 412526 532620 412530
rect 532556 412506 532620 412510
rect 532556 412450 532560 412506
rect 532560 412450 532616 412506
rect 532616 412450 532620 412506
rect 532556 412446 532620 412450
rect 536316 414026 536380 414030
rect 536316 413970 536320 414026
rect 536320 413970 536376 414026
rect 536376 413970 536380 414026
rect 536316 413966 536380 413970
rect 536316 413946 536380 413950
rect 536316 413890 536320 413946
rect 536320 413890 536376 413946
rect 536376 413890 536380 413946
rect 536316 413886 536380 413890
rect 536316 413866 536380 413870
rect 536316 413810 536320 413866
rect 536320 413810 536376 413866
rect 536376 413810 536380 413866
rect 536316 413806 536380 413810
rect 536316 413786 536380 413790
rect 536316 413730 536320 413786
rect 536320 413730 536376 413786
rect 536376 413730 536380 413786
rect 536316 413726 536380 413730
rect 536316 413706 536380 413710
rect 536316 413650 536320 413706
rect 536320 413650 536376 413706
rect 536376 413650 536380 413706
rect 536316 413646 536380 413650
rect 536316 413626 536380 413630
rect 536316 413570 536320 413626
rect 536320 413570 536376 413626
rect 536376 413570 536380 413626
rect 536316 413566 536380 413570
rect 536316 413546 536380 413550
rect 536316 413490 536320 413546
rect 536320 413490 536376 413546
rect 536376 413490 536380 413546
rect 536316 413486 536380 413490
rect 536316 413466 536380 413470
rect 536316 413410 536320 413466
rect 536320 413410 536376 413466
rect 536376 413410 536380 413466
rect 536316 413406 536380 413410
rect 536316 413386 536380 413390
rect 536316 413330 536320 413386
rect 536320 413330 536376 413386
rect 536376 413330 536380 413386
rect 536316 413326 536380 413330
rect 536316 413306 536380 413310
rect 536316 413250 536320 413306
rect 536320 413250 536376 413306
rect 536376 413250 536380 413306
rect 536316 413246 536380 413250
rect 536316 413226 536380 413230
rect 536316 413170 536320 413226
rect 536320 413170 536376 413226
rect 536376 413170 536380 413226
rect 536316 413166 536380 413170
rect 536316 413146 536380 413150
rect 536316 413090 536320 413146
rect 536320 413090 536376 413146
rect 536376 413090 536380 413146
rect 536316 413086 536380 413090
rect 536316 413066 536380 413070
rect 536316 413010 536320 413066
rect 536320 413010 536376 413066
rect 536376 413010 536380 413066
rect 536316 413006 536380 413010
rect 536316 412986 536380 412990
rect 536316 412930 536320 412986
rect 536320 412930 536376 412986
rect 536376 412930 536380 412986
rect 536316 412926 536380 412930
rect 536316 412906 536380 412910
rect 536316 412850 536320 412906
rect 536320 412850 536376 412906
rect 536376 412850 536380 412906
rect 536316 412846 536380 412850
rect 536316 412826 536380 412830
rect 536316 412770 536320 412826
rect 536320 412770 536376 412826
rect 536376 412770 536380 412826
rect 536316 412766 536380 412770
rect 536316 412746 536380 412750
rect 536316 412690 536320 412746
rect 536320 412690 536376 412746
rect 536376 412690 536380 412746
rect 536316 412686 536380 412690
rect 536316 412666 536380 412670
rect 536316 412610 536320 412666
rect 536320 412610 536376 412666
rect 536376 412610 536380 412666
rect 536316 412606 536380 412610
rect 536316 412586 536380 412590
rect 536316 412530 536320 412586
rect 536320 412530 536376 412586
rect 536376 412530 536380 412586
rect 536316 412526 536380 412530
rect 536316 412506 536380 412510
rect 536316 412450 536320 412506
rect 536320 412450 536376 412506
rect 536376 412450 536380 412506
rect 536316 412446 536380 412450
rect 504356 411578 504420 411582
rect 504356 411522 504360 411578
rect 504360 411522 504416 411578
rect 504416 411522 504420 411578
rect 504356 411518 504420 411522
rect 504356 411498 504420 411502
rect 504356 411442 504360 411498
rect 504360 411442 504416 411498
rect 504416 411442 504420 411498
rect 504356 411438 504420 411442
rect 504356 411418 504420 411422
rect 504356 411362 504360 411418
rect 504360 411362 504416 411418
rect 504416 411362 504420 411418
rect 504356 411358 504420 411362
rect 504356 411338 504420 411342
rect 504356 411282 504360 411338
rect 504360 411282 504416 411338
rect 504416 411282 504420 411338
rect 504356 411278 504420 411282
rect 504356 411258 504420 411262
rect 504356 411202 504360 411258
rect 504360 411202 504416 411258
rect 504416 411202 504420 411258
rect 504356 411198 504420 411202
rect 504356 411178 504420 411182
rect 504356 411122 504360 411178
rect 504360 411122 504416 411178
rect 504416 411122 504420 411178
rect 504356 411118 504420 411122
rect 504356 411098 504420 411102
rect 504356 411042 504360 411098
rect 504360 411042 504416 411098
rect 504416 411042 504420 411098
rect 504356 411038 504420 411042
rect 504356 411018 504420 411022
rect 504356 410962 504360 411018
rect 504360 410962 504416 411018
rect 504416 410962 504420 411018
rect 504356 410958 504420 410962
rect 504356 410938 504420 410942
rect 504356 410882 504360 410938
rect 504360 410882 504416 410938
rect 504416 410882 504420 410938
rect 504356 410878 504420 410882
rect 504356 410858 504420 410862
rect 504356 410802 504360 410858
rect 504360 410802 504416 410858
rect 504416 410802 504420 410858
rect 504356 410798 504420 410802
rect 504356 410778 504420 410782
rect 504356 410722 504360 410778
rect 504360 410722 504416 410778
rect 504416 410722 504420 410778
rect 504356 410718 504420 410722
rect 504356 410698 504420 410702
rect 504356 410642 504360 410698
rect 504360 410642 504416 410698
rect 504416 410642 504420 410698
rect 504356 410638 504420 410642
rect 504356 410618 504420 410622
rect 504356 410562 504360 410618
rect 504360 410562 504416 410618
rect 504416 410562 504420 410618
rect 504356 410558 504420 410562
rect 504356 410538 504420 410542
rect 504356 410482 504360 410538
rect 504360 410482 504416 410538
rect 504416 410482 504420 410538
rect 504356 410478 504420 410482
rect 504356 410458 504420 410462
rect 504356 410402 504360 410458
rect 504360 410402 504416 410458
rect 504416 410402 504420 410458
rect 504356 410398 504420 410402
rect 504356 410378 504420 410382
rect 504356 410322 504360 410378
rect 504360 410322 504416 410378
rect 504416 410322 504420 410378
rect 504356 410318 504420 410322
rect 504356 410298 504420 410302
rect 504356 410242 504360 410298
rect 504360 410242 504416 410298
rect 504416 410242 504420 410298
rect 504356 410238 504420 410242
rect 504356 410218 504420 410222
rect 504356 410162 504360 410218
rect 504360 410162 504416 410218
rect 504416 410162 504420 410218
rect 504356 410158 504420 410162
rect 504356 410138 504420 410142
rect 504356 410082 504360 410138
rect 504360 410082 504416 410138
rect 504416 410082 504420 410138
rect 504356 410078 504420 410082
rect 504356 410058 504420 410062
rect 504356 410002 504360 410058
rect 504360 410002 504416 410058
rect 504416 410002 504420 410058
rect 504356 409998 504420 410002
rect 508116 411578 508180 411582
rect 508116 411522 508120 411578
rect 508120 411522 508176 411578
rect 508176 411522 508180 411578
rect 508116 411518 508180 411522
rect 508116 411498 508180 411502
rect 508116 411442 508120 411498
rect 508120 411442 508176 411498
rect 508176 411442 508180 411498
rect 508116 411438 508180 411442
rect 508116 411418 508180 411422
rect 508116 411362 508120 411418
rect 508120 411362 508176 411418
rect 508176 411362 508180 411418
rect 508116 411358 508180 411362
rect 508116 411338 508180 411342
rect 508116 411282 508120 411338
rect 508120 411282 508176 411338
rect 508176 411282 508180 411338
rect 508116 411278 508180 411282
rect 508116 411258 508180 411262
rect 508116 411202 508120 411258
rect 508120 411202 508176 411258
rect 508176 411202 508180 411258
rect 508116 411198 508180 411202
rect 508116 411178 508180 411182
rect 508116 411122 508120 411178
rect 508120 411122 508176 411178
rect 508176 411122 508180 411178
rect 508116 411118 508180 411122
rect 508116 411098 508180 411102
rect 508116 411042 508120 411098
rect 508120 411042 508176 411098
rect 508176 411042 508180 411098
rect 508116 411038 508180 411042
rect 508116 411018 508180 411022
rect 508116 410962 508120 411018
rect 508120 410962 508176 411018
rect 508176 410962 508180 411018
rect 508116 410958 508180 410962
rect 508116 410938 508180 410942
rect 508116 410882 508120 410938
rect 508120 410882 508176 410938
rect 508176 410882 508180 410938
rect 508116 410878 508180 410882
rect 508116 410858 508180 410862
rect 508116 410802 508120 410858
rect 508120 410802 508176 410858
rect 508176 410802 508180 410858
rect 508116 410798 508180 410802
rect 508116 410778 508180 410782
rect 508116 410722 508120 410778
rect 508120 410722 508176 410778
rect 508176 410722 508180 410778
rect 508116 410718 508180 410722
rect 508116 410698 508180 410702
rect 508116 410642 508120 410698
rect 508120 410642 508176 410698
rect 508176 410642 508180 410698
rect 508116 410638 508180 410642
rect 508116 410618 508180 410622
rect 508116 410562 508120 410618
rect 508120 410562 508176 410618
rect 508176 410562 508180 410618
rect 508116 410558 508180 410562
rect 508116 410538 508180 410542
rect 508116 410482 508120 410538
rect 508120 410482 508176 410538
rect 508176 410482 508180 410538
rect 508116 410478 508180 410482
rect 508116 410458 508180 410462
rect 508116 410402 508120 410458
rect 508120 410402 508176 410458
rect 508176 410402 508180 410458
rect 508116 410398 508180 410402
rect 508116 410378 508180 410382
rect 508116 410322 508120 410378
rect 508120 410322 508176 410378
rect 508176 410322 508180 410378
rect 508116 410318 508180 410322
rect 508116 410298 508180 410302
rect 508116 410242 508120 410298
rect 508120 410242 508176 410298
rect 508176 410242 508180 410298
rect 508116 410238 508180 410242
rect 508116 410218 508180 410222
rect 508116 410162 508120 410218
rect 508120 410162 508176 410218
rect 508176 410162 508180 410218
rect 508116 410158 508180 410162
rect 508116 410138 508180 410142
rect 508116 410082 508120 410138
rect 508120 410082 508176 410138
rect 508176 410082 508180 410138
rect 508116 410078 508180 410082
rect 508116 410058 508180 410062
rect 508116 410002 508120 410058
rect 508120 410002 508176 410058
rect 508176 410002 508180 410058
rect 508116 409998 508180 410002
rect 511876 411578 511940 411582
rect 511876 411522 511880 411578
rect 511880 411522 511936 411578
rect 511936 411522 511940 411578
rect 511876 411518 511940 411522
rect 511876 411498 511940 411502
rect 511876 411442 511880 411498
rect 511880 411442 511936 411498
rect 511936 411442 511940 411498
rect 511876 411438 511940 411442
rect 511876 411418 511940 411422
rect 511876 411362 511880 411418
rect 511880 411362 511936 411418
rect 511936 411362 511940 411418
rect 511876 411358 511940 411362
rect 511876 411338 511940 411342
rect 511876 411282 511880 411338
rect 511880 411282 511936 411338
rect 511936 411282 511940 411338
rect 511876 411278 511940 411282
rect 511876 411258 511940 411262
rect 511876 411202 511880 411258
rect 511880 411202 511936 411258
rect 511936 411202 511940 411258
rect 511876 411198 511940 411202
rect 511876 411178 511940 411182
rect 511876 411122 511880 411178
rect 511880 411122 511936 411178
rect 511936 411122 511940 411178
rect 511876 411118 511940 411122
rect 511876 411098 511940 411102
rect 511876 411042 511880 411098
rect 511880 411042 511936 411098
rect 511936 411042 511940 411098
rect 511876 411038 511940 411042
rect 511876 411018 511940 411022
rect 511876 410962 511880 411018
rect 511880 410962 511936 411018
rect 511936 410962 511940 411018
rect 511876 410958 511940 410962
rect 511876 410938 511940 410942
rect 511876 410882 511880 410938
rect 511880 410882 511936 410938
rect 511936 410882 511940 410938
rect 511876 410878 511940 410882
rect 511876 410858 511940 410862
rect 511876 410802 511880 410858
rect 511880 410802 511936 410858
rect 511936 410802 511940 410858
rect 511876 410798 511940 410802
rect 511876 410778 511940 410782
rect 511876 410722 511880 410778
rect 511880 410722 511936 410778
rect 511936 410722 511940 410778
rect 511876 410718 511940 410722
rect 511876 410698 511940 410702
rect 511876 410642 511880 410698
rect 511880 410642 511936 410698
rect 511936 410642 511940 410698
rect 511876 410638 511940 410642
rect 511876 410618 511940 410622
rect 511876 410562 511880 410618
rect 511880 410562 511936 410618
rect 511936 410562 511940 410618
rect 511876 410558 511940 410562
rect 511876 410538 511940 410542
rect 511876 410482 511880 410538
rect 511880 410482 511936 410538
rect 511936 410482 511940 410538
rect 511876 410478 511940 410482
rect 511876 410458 511940 410462
rect 511876 410402 511880 410458
rect 511880 410402 511936 410458
rect 511936 410402 511940 410458
rect 511876 410398 511940 410402
rect 511876 410378 511940 410382
rect 511876 410322 511880 410378
rect 511880 410322 511936 410378
rect 511936 410322 511940 410378
rect 511876 410318 511940 410322
rect 511876 410298 511940 410302
rect 511876 410242 511880 410298
rect 511880 410242 511936 410298
rect 511936 410242 511940 410298
rect 511876 410238 511940 410242
rect 511876 410218 511940 410222
rect 511876 410162 511880 410218
rect 511880 410162 511936 410218
rect 511936 410162 511940 410218
rect 511876 410158 511940 410162
rect 511876 410138 511940 410142
rect 511876 410082 511880 410138
rect 511880 410082 511936 410138
rect 511936 410082 511940 410138
rect 511876 410078 511940 410082
rect 511876 410058 511940 410062
rect 511876 410002 511880 410058
rect 511880 410002 511936 410058
rect 511936 410002 511940 410058
rect 511876 409998 511940 410002
rect 515636 411578 515700 411582
rect 515636 411522 515640 411578
rect 515640 411522 515696 411578
rect 515696 411522 515700 411578
rect 515636 411518 515700 411522
rect 515636 411498 515700 411502
rect 515636 411442 515640 411498
rect 515640 411442 515696 411498
rect 515696 411442 515700 411498
rect 515636 411438 515700 411442
rect 515636 411418 515700 411422
rect 515636 411362 515640 411418
rect 515640 411362 515696 411418
rect 515696 411362 515700 411418
rect 515636 411358 515700 411362
rect 515636 411338 515700 411342
rect 515636 411282 515640 411338
rect 515640 411282 515696 411338
rect 515696 411282 515700 411338
rect 515636 411278 515700 411282
rect 515636 411258 515700 411262
rect 515636 411202 515640 411258
rect 515640 411202 515696 411258
rect 515696 411202 515700 411258
rect 515636 411198 515700 411202
rect 515636 411178 515700 411182
rect 515636 411122 515640 411178
rect 515640 411122 515696 411178
rect 515696 411122 515700 411178
rect 515636 411118 515700 411122
rect 515636 411098 515700 411102
rect 515636 411042 515640 411098
rect 515640 411042 515696 411098
rect 515696 411042 515700 411098
rect 515636 411038 515700 411042
rect 515636 411018 515700 411022
rect 515636 410962 515640 411018
rect 515640 410962 515696 411018
rect 515696 410962 515700 411018
rect 515636 410958 515700 410962
rect 515636 410938 515700 410942
rect 515636 410882 515640 410938
rect 515640 410882 515696 410938
rect 515696 410882 515700 410938
rect 515636 410878 515700 410882
rect 515636 410858 515700 410862
rect 515636 410802 515640 410858
rect 515640 410802 515696 410858
rect 515696 410802 515700 410858
rect 515636 410798 515700 410802
rect 515636 410778 515700 410782
rect 515636 410722 515640 410778
rect 515640 410722 515696 410778
rect 515696 410722 515700 410778
rect 515636 410718 515700 410722
rect 515636 410698 515700 410702
rect 515636 410642 515640 410698
rect 515640 410642 515696 410698
rect 515696 410642 515700 410698
rect 515636 410638 515700 410642
rect 515636 410618 515700 410622
rect 515636 410562 515640 410618
rect 515640 410562 515696 410618
rect 515696 410562 515700 410618
rect 515636 410558 515700 410562
rect 515636 410538 515700 410542
rect 515636 410482 515640 410538
rect 515640 410482 515696 410538
rect 515696 410482 515700 410538
rect 515636 410478 515700 410482
rect 515636 410458 515700 410462
rect 515636 410402 515640 410458
rect 515640 410402 515696 410458
rect 515696 410402 515700 410458
rect 515636 410398 515700 410402
rect 515636 410378 515700 410382
rect 515636 410322 515640 410378
rect 515640 410322 515696 410378
rect 515696 410322 515700 410378
rect 515636 410318 515700 410322
rect 515636 410298 515700 410302
rect 515636 410242 515640 410298
rect 515640 410242 515696 410298
rect 515696 410242 515700 410298
rect 515636 410238 515700 410242
rect 515636 410218 515700 410222
rect 515636 410162 515640 410218
rect 515640 410162 515696 410218
rect 515696 410162 515700 410218
rect 515636 410158 515700 410162
rect 515636 410138 515700 410142
rect 515636 410082 515640 410138
rect 515640 410082 515696 410138
rect 515696 410082 515700 410138
rect 515636 410078 515700 410082
rect 515636 410058 515700 410062
rect 515636 410002 515640 410058
rect 515640 410002 515696 410058
rect 515696 410002 515700 410058
rect 515636 409998 515700 410002
rect 519396 411578 519460 411582
rect 519396 411522 519400 411578
rect 519400 411522 519456 411578
rect 519456 411522 519460 411578
rect 519396 411518 519460 411522
rect 519396 411498 519460 411502
rect 519396 411442 519400 411498
rect 519400 411442 519456 411498
rect 519456 411442 519460 411498
rect 519396 411438 519460 411442
rect 519396 411418 519460 411422
rect 519396 411362 519400 411418
rect 519400 411362 519456 411418
rect 519456 411362 519460 411418
rect 519396 411358 519460 411362
rect 519396 411338 519460 411342
rect 519396 411282 519400 411338
rect 519400 411282 519456 411338
rect 519456 411282 519460 411338
rect 519396 411278 519460 411282
rect 519396 411258 519460 411262
rect 519396 411202 519400 411258
rect 519400 411202 519456 411258
rect 519456 411202 519460 411258
rect 519396 411198 519460 411202
rect 519396 411178 519460 411182
rect 519396 411122 519400 411178
rect 519400 411122 519456 411178
rect 519456 411122 519460 411178
rect 519396 411118 519460 411122
rect 519396 411098 519460 411102
rect 519396 411042 519400 411098
rect 519400 411042 519456 411098
rect 519456 411042 519460 411098
rect 519396 411038 519460 411042
rect 519396 411018 519460 411022
rect 519396 410962 519400 411018
rect 519400 410962 519456 411018
rect 519456 410962 519460 411018
rect 519396 410958 519460 410962
rect 519396 410938 519460 410942
rect 519396 410882 519400 410938
rect 519400 410882 519456 410938
rect 519456 410882 519460 410938
rect 519396 410878 519460 410882
rect 519396 410858 519460 410862
rect 519396 410802 519400 410858
rect 519400 410802 519456 410858
rect 519456 410802 519460 410858
rect 519396 410798 519460 410802
rect 519396 410778 519460 410782
rect 519396 410722 519400 410778
rect 519400 410722 519456 410778
rect 519456 410722 519460 410778
rect 519396 410718 519460 410722
rect 519396 410698 519460 410702
rect 519396 410642 519400 410698
rect 519400 410642 519456 410698
rect 519456 410642 519460 410698
rect 519396 410638 519460 410642
rect 519396 410618 519460 410622
rect 519396 410562 519400 410618
rect 519400 410562 519456 410618
rect 519456 410562 519460 410618
rect 519396 410558 519460 410562
rect 519396 410538 519460 410542
rect 519396 410482 519400 410538
rect 519400 410482 519456 410538
rect 519456 410482 519460 410538
rect 519396 410478 519460 410482
rect 519396 410458 519460 410462
rect 519396 410402 519400 410458
rect 519400 410402 519456 410458
rect 519456 410402 519460 410458
rect 519396 410398 519460 410402
rect 519396 410378 519460 410382
rect 519396 410322 519400 410378
rect 519400 410322 519456 410378
rect 519456 410322 519460 410378
rect 519396 410318 519460 410322
rect 519396 410298 519460 410302
rect 519396 410242 519400 410298
rect 519400 410242 519456 410298
rect 519456 410242 519460 410298
rect 519396 410238 519460 410242
rect 519396 410218 519460 410222
rect 519396 410162 519400 410218
rect 519400 410162 519456 410218
rect 519456 410162 519460 410218
rect 519396 410158 519460 410162
rect 519396 410138 519460 410142
rect 519396 410082 519400 410138
rect 519400 410082 519456 410138
rect 519456 410082 519460 410138
rect 519396 410078 519460 410082
rect 519396 410058 519460 410062
rect 519396 410002 519400 410058
rect 519400 410002 519456 410058
rect 519456 410002 519460 410058
rect 519396 409998 519460 410002
rect 523156 411578 523220 411582
rect 523156 411522 523160 411578
rect 523160 411522 523216 411578
rect 523216 411522 523220 411578
rect 523156 411518 523220 411522
rect 523156 411498 523220 411502
rect 523156 411442 523160 411498
rect 523160 411442 523216 411498
rect 523216 411442 523220 411498
rect 523156 411438 523220 411442
rect 523156 411418 523220 411422
rect 523156 411362 523160 411418
rect 523160 411362 523216 411418
rect 523216 411362 523220 411418
rect 523156 411358 523220 411362
rect 523156 411338 523220 411342
rect 523156 411282 523160 411338
rect 523160 411282 523216 411338
rect 523216 411282 523220 411338
rect 523156 411278 523220 411282
rect 523156 411258 523220 411262
rect 523156 411202 523160 411258
rect 523160 411202 523216 411258
rect 523216 411202 523220 411258
rect 523156 411198 523220 411202
rect 523156 411178 523220 411182
rect 523156 411122 523160 411178
rect 523160 411122 523216 411178
rect 523216 411122 523220 411178
rect 523156 411118 523220 411122
rect 523156 411098 523220 411102
rect 523156 411042 523160 411098
rect 523160 411042 523216 411098
rect 523216 411042 523220 411098
rect 523156 411038 523220 411042
rect 523156 411018 523220 411022
rect 523156 410962 523160 411018
rect 523160 410962 523216 411018
rect 523216 410962 523220 411018
rect 523156 410958 523220 410962
rect 523156 410938 523220 410942
rect 523156 410882 523160 410938
rect 523160 410882 523216 410938
rect 523216 410882 523220 410938
rect 523156 410878 523220 410882
rect 523156 410858 523220 410862
rect 523156 410802 523160 410858
rect 523160 410802 523216 410858
rect 523216 410802 523220 410858
rect 523156 410798 523220 410802
rect 523156 410778 523220 410782
rect 523156 410722 523160 410778
rect 523160 410722 523216 410778
rect 523216 410722 523220 410778
rect 523156 410718 523220 410722
rect 523156 410698 523220 410702
rect 523156 410642 523160 410698
rect 523160 410642 523216 410698
rect 523216 410642 523220 410698
rect 523156 410638 523220 410642
rect 523156 410618 523220 410622
rect 523156 410562 523160 410618
rect 523160 410562 523216 410618
rect 523216 410562 523220 410618
rect 523156 410558 523220 410562
rect 523156 410538 523220 410542
rect 523156 410482 523160 410538
rect 523160 410482 523216 410538
rect 523216 410482 523220 410538
rect 523156 410478 523220 410482
rect 523156 410458 523220 410462
rect 523156 410402 523160 410458
rect 523160 410402 523216 410458
rect 523216 410402 523220 410458
rect 523156 410398 523220 410402
rect 523156 410378 523220 410382
rect 523156 410322 523160 410378
rect 523160 410322 523216 410378
rect 523216 410322 523220 410378
rect 523156 410318 523220 410322
rect 523156 410298 523220 410302
rect 523156 410242 523160 410298
rect 523160 410242 523216 410298
rect 523216 410242 523220 410298
rect 523156 410238 523220 410242
rect 523156 410218 523220 410222
rect 523156 410162 523160 410218
rect 523160 410162 523216 410218
rect 523216 410162 523220 410218
rect 523156 410158 523220 410162
rect 523156 410138 523220 410142
rect 523156 410082 523160 410138
rect 523160 410082 523216 410138
rect 523216 410082 523220 410138
rect 523156 410078 523220 410082
rect 523156 410058 523220 410062
rect 523156 410002 523160 410058
rect 523160 410002 523216 410058
rect 523216 410002 523220 410058
rect 523156 409998 523220 410002
rect 526916 411578 526980 411582
rect 526916 411522 526920 411578
rect 526920 411522 526976 411578
rect 526976 411522 526980 411578
rect 526916 411518 526980 411522
rect 526916 411498 526980 411502
rect 526916 411442 526920 411498
rect 526920 411442 526976 411498
rect 526976 411442 526980 411498
rect 526916 411438 526980 411442
rect 526916 411418 526980 411422
rect 526916 411362 526920 411418
rect 526920 411362 526976 411418
rect 526976 411362 526980 411418
rect 526916 411358 526980 411362
rect 526916 411338 526980 411342
rect 526916 411282 526920 411338
rect 526920 411282 526976 411338
rect 526976 411282 526980 411338
rect 526916 411278 526980 411282
rect 526916 411258 526980 411262
rect 526916 411202 526920 411258
rect 526920 411202 526976 411258
rect 526976 411202 526980 411258
rect 526916 411198 526980 411202
rect 526916 411178 526980 411182
rect 526916 411122 526920 411178
rect 526920 411122 526976 411178
rect 526976 411122 526980 411178
rect 526916 411118 526980 411122
rect 526916 411098 526980 411102
rect 526916 411042 526920 411098
rect 526920 411042 526976 411098
rect 526976 411042 526980 411098
rect 526916 411038 526980 411042
rect 526916 411018 526980 411022
rect 526916 410962 526920 411018
rect 526920 410962 526976 411018
rect 526976 410962 526980 411018
rect 526916 410958 526980 410962
rect 526916 410938 526980 410942
rect 526916 410882 526920 410938
rect 526920 410882 526976 410938
rect 526976 410882 526980 410938
rect 526916 410878 526980 410882
rect 526916 410858 526980 410862
rect 526916 410802 526920 410858
rect 526920 410802 526976 410858
rect 526976 410802 526980 410858
rect 526916 410798 526980 410802
rect 526916 410778 526980 410782
rect 526916 410722 526920 410778
rect 526920 410722 526976 410778
rect 526976 410722 526980 410778
rect 526916 410718 526980 410722
rect 526916 410698 526980 410702
rect 526916 410642 526920 410698
rect 526920 410642 526976 410698
rect 526976 410642 526980 410698
rect 526916 410638 526980 410642
rect 526916 410618 526980 410622
rect 526916 410562 526920 410618
rect 526920 410562 526976 410618
rect 526976 410562 526980 410618
rect 526916 410558 526980 410562
rect 526916 410538 526980 410542
rect 526916 410482 526920 410538
rect 526920 410482 526976 410538
rect 526976 410482 526980 410538
rect 526916 410478 526980 410482
rect 526916 410458 526980 410462
rect 526916 410402 526920 410458
rect 526920 410402 526976 410458
rect 526976 410402 526980 410458
rect 526916 410398 526980 410402
rect 526916 410378 526980 410382
rect 526916 410322 526920 410378
rect 526920 410322 526976 410378
rect 526976 410322 526980 410378
rect 526916 410318 526980 410322
rect 526916 410298 526980 410302
rect 526916 410242 526920 410298
rect 526920 410242 526976 410298
rect 526976 410242 526980 410298
rect 526916 410238 526980 410242
rect 526916 410218 526980 410222
rect 526916 410162 526920 410218
rect 526920 410162 526976 410218
rect 526976 410162 526980 410218
rect 526916 410158 526980 410162
rect 526916 410138 526980 410142
rect 526916 410082 526920 410138
rect 526920 410082 526976 410138
rect 526976 410082 526980 410138
rect 526916 410078 526980 410082
rect 526916 410058 526980 410062
rect 526916 410002 526920 410058
rect 526920 410002 526976 410058
rect 526976 410002 526980 410058
rect 526916 409998 526980 410002
rect 530676 411578 530740 411582
rect 530676 411522 530680 411578
rect 530680 411522 530736 411578
rect 530736 411522 530740 411578
rect 530676 411518 530740 411522
rect 530676 411498 530740 411502
rect 530676 411442 530680 411498
rect 530680 411442 530736 411498
rect 530736 411442 530740 411498
rect 530676 411438 530740 411442
rect 530676 411418 530740 411422
rect 530676 411362 530680 411418
rect 530680 411362 530736 411418
rect 530736 411362 530740 411418
rect 530676 411358 530740 411362
rect 530676 411338 530740 411342
rect 530676 411282 530680 411338
rect 530680 411282 530736 411338
rect 530736 411282 530740 411338
rect 530676 411278 530740 411282
rect 530676 411258 530740 411262
rect 530676 411202 530680 411258
rect 530680 411202 530736 411258
rect 530736 411202 530740 411258
rect 530676 411198 530740 411202
rect 530676 411178 530740 411182
rect 530676 411122 530680 411178
rect 530680 411122 530736 411178
rect 530736 411122 530740 411178
rect 530676 411118 530740 411122
rect 530676 411098 530740 411102
rect 530676 411042 530680 411098
rect 530680 411042 530736 411098
rect 530736 411042 530740 411098
rect 530676 411038 530740 411042
rect 530676 411018 530740 411022
rect 530676 410962 530680 411018
rect 530680 410962 530736 411018
rect 530736 410962 530740 411018
rect 530676 410958 530740 410962
rect 530676 410938 530740 410942
rect 530676 410882 530680 410938
rect 530680 410882 530736 410938
rect 530736 410882 530740 410938
rect 530676 410878 530740 410882
rect 530676 410858 530740 410862
rect 530676 410802 530680 410858
rect 530680 410802 530736 410858
rect 530736 410802 530740 410858
rect 530676 410798 530740 410802
rect 530676 410778 530740 410782
rect 530676 410722 530680 410778
rect 530680 410722 530736 410778
rect 530736 410722 530740 410778
rect 530676 410718 530740 410722
rect 530676 410698 530740 410702
rect 530676 410642 530680 410698
rect 530680 410642 530736 410698
rect 530736 410642 530740 410698
rect 530676 410638 530740 410642
rect 530676 410618 530740 410622
rect 530676 410562 530680 410618
rect 530680 410562 530736 410618
rect 530736 410562 530740 410618
rect 530676 410558 530740 410562
rect 530676 410538 530740 410542
rect 530676 410482 530680 410538
rect 530680 410482 530736 410538
rect 530736 410482 530740 410538
rect 530676 410478 530740 410482
rect 530676 410458 530740 410462
rect 530676 410402 530680 410458
rect 530680 410402 530736 410458
rect 530736 410402 530740 410458
rect 530676 410398 530740 410402
rect 530676 410378 530740 410382
rect 530676 410322 530680 410378
rect 530680 410322 530736 410378
rect 530736 410322 530740 410378
rect 530676 410318 530740 410322
rect 530676 410298 530740 410302
rect 530676 410242 530680 410298
rect 530680 410242 530736 410298
rect 530736 410242 530740 410298
rect 530676 410238 530740 410242
rect 530676 410218 530740 410222
rect 530676 410162 530680 410218
rect 530680 410162 530736 410218
rect 530736 410162 530740 410218
rect 530676 410158 530740 410162
rect 530676 410138 530740 410142
rect 530676 410082 530680 410138
rect 530680 410082 530736 410138
rect 530736 410082 530740 410138
rect 530676 410078 530740 410082
rect 530676 410058 530740 410062
rect 530676 410002 530680 410058
rect 530680 410002 530736 410058
rect 530736 410002 530740 410058
rect 530676 409998 530740 410002
rect 534436 411578 534500 411582
rect 534436 411522 534440 411578
rect 534440 411522 534496 411578
rect 534496 411522 534500 411578
rect 534436 411518 534500 411522
rect 534436 411498 534500 411502
rect 534436 411442 534440 411498
rect 534440 411442 534496 411498
rect 534496 411442 534500 411498
rect 534436 411438 534500 411442
rect 534436 411418 534500 411422
rect 534436 411362 534440 411418
rect 534440 411362 534496 411418
rect 534496 411362 534500 411418
rect 534436 411358 534500 411362
rect 534436 411338 534500 411342
rect 534436 411282 534440 411338
rect 534440 411282 534496 411338
rect 534496 411282 534500 411338
rect 534436 411278 534500 411282
rect 534436 411258 534500 411262
rect 534436 411202 534440 411258
rect 534440 411202 534496 411258
rect 534496 411202 534500 411258
rect 534436 411198 534500 411202
rect 534436 411178 534500 411182
rect 534436 411122 534440 411178
rect 534440 411122 534496 411178
rect 534496 411122 534500 411178
rect 534436 411118 534500 411122
rect 534436 411098 534500 411102
rect 534436 411042 534440 411098
rect 534440 411042 534496 411098
rect 534496 411042 534500 411098
rect 534436 411038 534500 411042
rect 534436 411018 534500 411022
rect 534436 410962 534440 411018
rect 534440 410962 534496 411018
rect 534496 410962 534500 411018
rect 534436 410958 534500 410962
rect 534436 410938 534500 410942
rect 534436 410882 534440 410938
rect 534440 410882 534496 410938
rect 534496 410882 534500 410938
rect 534436 410878 534500 410882
rect 534436 410858 534500 410862
rect 534436 410802 534440 410858
rect 534440 410802 534496 410858
rect 534496 410802 534500 410858
rect 534436 410798 534500 410802
rect 534436 410778 534500 410782
rect 534436 410722 534440 410778
rect 534440 410722 534496 410778
rect 534496 410722 534500 410778
rect 534436 410718 534500 410722
rect 534436 410698 534500 410702
rect 534436 410642 534440 410698
rect 534440 410642 534496 410698
rect 534496 410642 534500 410698
rect 534436 410638 534500 410642
rect 534436 410618 534500 410622
rect 534436 410562 534440 410618
rect 534440 410562 534496 410618
rect 534496 410562 534500 410618
rect 534436 410558 534500 410562
rect 534436 410538 534500 410542
rect 534436 410482 534440 410538
rect 534440 410482 534496 410538
rect 534496 410482 534500 410538
rect 534436 410478 534500 410482
rect 534436 410458 534500 410462
rect 534436 410402 534440 410458
rect 534440 410402 534496 410458
rect 534496 410402 534500 410458
rect 534436 410398 534500 410402
rect 534436 410378 534500 410382
rect 534436 410322 534440 410378
rect 534440 410322 534496 410378
rect 534496 410322 534500 410378
rect 534436 410318 534500 410322
rect 534436 410298 534500 410302
rect 534436 410242 534440 410298
rect 534440 410242 534496 410298
rect 534496 410242 534500 410298
rect 534436 410238 534500 410242
rect 534436 410218 534500 410222
rect 534436 410162 534440 410218
rect 534440 410162 534496 410218
rect 534496 410162 534500 410218
rect 534436 410158 534500 410162
rect 534436 410138 534500 410142
rect 534436 410082 534440 410138
rect 534440 410082 534496 410138
rect 534496 410082 534500 410138
rect 534436 410078 534500 410082
rect 534436 410058 534500 410062
rect 534436 410002 534440 410058
rect 534440 410002 534496 410058
rect 534496 410002 534500 410058
rect 534436 409998 534500 410002
rect 494766 408964 494830 409008
rect 494766 408944 494770 408964
rect 494770 408944 494826 408964
rect 494826 408944 494830 408964
rect 494766 408908 494770 408928
rect 494770 408908 494826 408928
rect 494826 408908 494830 408928
rect 494766 408864 494830 408908
rect 493366 408358 493430 408422
rect 493446 408358 493510 408422
rect 493526 408358 493590 408422
rect 493606 408358 493670 408422
rect 493686 408358 493750 408422
rect 493766 408358 493830 408422
rect 493846 408358 493910 408422
rect 494066 408358 494130 408422
rect 494146 408358 494210 408422
rect 494226 408358 494290 408422
rect 494306 408358 494370 408422
rect 494386 408358 494450 408422
rect 494466 408358 494530 408422
rect 494546 408358 494610 408422
rect 493366 407639 493430 407703
rect 493446 407639 493510 407703
rect 493526 407639 493590 407703
rect 493606 407639 493670 407703
rect 493686 407639 493750 407703
rect 493766 407639 493830 407703
rect 493846 407639 493910 407703
rect 494066 407639 494130 407703
rect 494146 407639 494210 407703
rect 494226 407639 494290 407703
rect 494306 407639 494370 407703
rect 494386 407639 494450 407703
rect 494466 407639 494530 407703
rect 494546 407639 494610 407703
rect 493366 406920 493430 406984
rect 493446 406920 493510 406984
rect 493526 406920 493590 406984
rect 493606 406920 493670 406984
rect 493686 406920 493750 406984
rect 493766 406920 493830 406984
rect 493846 406920 493910 406984
rect 494066 406920 494130 406984
rect 494146 406920 494210 406984
rect 494226 406920 494290 406984
rect 494306 406920 494370 406984
rect 494386 406920 494450 406984
rect 494466 406920 494530 406984
rect 494546 406920 494610 406984
rect 493366 406201 493430 406265
rect 493446 406201 493510 406265
rect 493526 406201 493590 406265
rect 493606 406201 493670 406265
rect 493686 406201 493750 406265
rect 493766 406201 493830 406265
rect 493846 406201 493910 406265
rect 494066 406201 494130 406265
rect 494146 406201 494210 406265
rect 494226 406201 494290 406265
rect 494306 406201 494370 406265
rect 494386 406201 494450 406265
rect 494466 406201 494530 406265
rect 494546 406201 494610 406265
rect 493366 405482 493430 405546
rect 493446 405482 493510 405546
rect 493526 405482 493590 405546
rect 493606 405482 493670 405546
rect 493686 405482 493750 405546
rect 493766 405482 493830 405546
rect 493846 405482 493910 405546
rect 494066 405482 494130 405546
rect 494146 405482 494210 405546
rect 494226 405482 494290 405546
rect 494306 405482 494370 405546
rect 494386 405482 494450 405546
rect 494466 405482 494530 405546
rect 494546 405482 494610 405546
rect 493366 404763 493430 404827
rect 493446 404763 493510 404827
rect 493526 404763 493590 404827
rect 493606 404763 493670 404827
rect 493686 404763 493750 404827
rect 493766 404763 493830 404827
rect 493846 404763 493910 404827
rect 494066 404763 494130 404827
rect 494146 404763 494210 404827
rect 494226 404763 494290 404827
rect 494306 404763 494370 404827
rect 494386 404763 494450 404827
rect 494466 404763 494530 404827
rect 494546 404763 494610 404827
rect 493366 404044 493430 404108
rect 493446 404044 493510 404108
rect 493526 404044 493590 404108
rect 493606 404044 493670 404108
rect 493686 404044 493750 404108
rect 493766 404044 493830 404108
rect 493846 404044 493910 404108
rect 494066 404044 494130 404108
rect 494146 404044 494210 404108
rect 494226 404044 494290 404108
rect 494306 404044 494370 404108
rect 494386 404044 494450 404108
rect 494466 404044 494530 404108
rect 494546 404044 494610 404108
rect 493366 403325 493430 403389
rect 493446 403325 493510 403389
rect 493526 403325 493590 403389
rect 493606 403325 493670 403389
rect 493686 403325 493750 403389
rect 493766 403325 493830 403389
rect 493846 403325 493910 403389
rect 494066 403325 494130 403389
rect 494146 403325 494210 403389
rect 494226 403325 494290 403389
rect 494306 403325 494370 403389
rect 494386 403325 494450 403389
rect 494466 403325 494530 403389
rect 494546 403325 494610 403389
rect 493366 402606 493430 402670
rect 493446 402606 493510 402670
rect 493526 402606 493590 402670
rect 493606 402606 493670 402670
rect 493686 402606 493750 402670
rect 493766 402606 493830 402670
rect 493846 402606 493910 402670
rect 494066 402606 494130 402670
rect 494146 402606 494210 402670
rect 494226 402606 494290 402670
rect 494306 402606 494370 402670
rect 494386 402606 494450 402670
rect 494466 402606 494530 402670
rect 494546 402606 494610 402670
rect 493366 401887 493430 401951
rect 493446 401887 493510 401951
rect 493526 401887 493590 401951
rect 493606 401887 493670 401951
rect 493686 401887 493750 401951
rect 493766 401887 493830 401951
rect 493846 401887 493910 401951
rect 494066 401887 494130 401951
rect 494146 401887 494210 401951
rect 494226 401887 494290 401951
rect 494306 401887 494370 401951
rect 494386 401887 494450 401951
rect 494466 401887 494530 401951
rect 494546 401887 494610 401951
rect 498526 408964 498590 409008
rect 498526 408944 498530 408964
rect 498530 408944 498586 408964
rect 498586 408944 498590 408964
rect 498526 408908 498530 408928
rect 498530 408908 498586 408928
rect 498586 408908 498590 408928
rect 498526 408864 498590 408908
rect 497126 408358 497190 408422
rect 497206 408358 497270 408422
rect 497286 408358 497350 408422
rect 497366 408358 497430 408422
rect 497446 408358 497510 408422
rect 497526 408358 497590 408422
rect 497606 408358 497670 408422
rect 497826 408358 497890 408422
rect 497906 408358 497970 408422
rect 497986 408358 498050 408422
rect 498066 408358 498130 408422
rect 498146 408358 498210 408422
rect 498226 408358 498290 408422
rect 498306 408358 498370 408422
rect 500658 407976 500722 408040
rect 502286 408572 502350 408616
rect 502286 408552 502290 408572
rect 502290 408552 502346 408572
rect 502346 408552 502350 408572
rect 502286 408516 502290 408536
rect 502290 408516 502346 408536
rect 502346 408516 502350 408536
rect 502286 408472 502350 408516
rect 497126 407639 497190 407703
rect 497206 407639 497270 407703
rect 497286 407639 497350 407703
rect 497366 407639 497430 407703
rect 497446 407639 497510 407703
rect 497526 407639 497590 407703
rect 497606 407639 497670 407703
rect 497826 407639 497890 407703
rect 497906 407639 497970 407703
rect 497986 407639 498050 407703
rect 498066 407639 498130 407703
rect 498146 407639 498210 407703
rect 498226 407639 498290 407703
rect 498306 407639 498370 407703
rect 497126 406920 497190 406984
rect 497206 406920 497270 406984
rect 497286 406920 497350 406984
rect 497366 406920 497430 406984
rect 497446 406920 497510 406984
rect 497526 406920 497590 406984
rect 497606 406920 497670 406984
rect 497826 406920 497890 406984
rect 497906 406920 497970 406984
rect 497986 406920 498050 406984
rect 498066 406920 498130 406984
rect 498146 406920 498210 406984
rect 498226 406920 498290 406984
rect 498306 406920 498370 406984
rect 500886 407966 500950 408030
rect 500966 407966 501030 408030
rect 501046 407966 501110 408030
rect 501126 407966 501190 408030
rect 501206 407966 501270 408030
rect 501286 407966 501350 408030
rect 501366 407966 501430 408030
rect 501586 407966 501650 408030
rect 501666 407966 501730 408030
rect 501746 407966 501810 408030
rect 501826 407966 501890 408030
rect 501906 407966 501970 408030
rect 501986 407966 502050 408030
rect 502066 407966 502130 408030
rect 500886 407247 500950 407311
rect 500966 407247 501030 407311
rect 501046 407247 501110 407311
rect 501126 407247 501190 407311
rect 501206 407247 501270 407311
rect 501286 407247 501350 407311
rect 501366 407247 501430 407311
rect 501586 407247 501650 407311
rect 501666 407247 501730 407311
rect 501746 407247 501810 407311
rect 501826 407247 501890 407311
rect 501906 407247 501970 407311
rect 501986 407247 502050 407311
rect 502066 407247 502130 407311
rect 498706 406656 498770 406660
rect 498706 406600 498710 406656
rect 498710 406600 498766 406656
rect 498766 406600 498770 406656
rect 498706 406596 498770 406600
rect 500886 406528 500950 406592
rect 500966 406528 501030 406592
rect 501046 406528 501110 406592
rect 501126 406528 501190 406592
rect 501206 406528 501270 406592
rect 501286 406528 501350 406592
rect 501366 406528 501430 406592
rect 501586 406528 501650 406592
rect 501666 406528 501730 406592
rect 501746 406528 501810 406592
rect 501826 406528 501890 406592
rect 501906 406528 501970 406592
rect 501986 406528 502050 406592
rect 502066 406528 502130 406592
rect 497126 406201 497190 406265
rect 497206 406201 497270 406265
rect 497286 406201 497350 406265
rect 497366 406201 497430 406265
rect 497446 406201 497510 406265
rect 497526 406201 497590 406265
rect 497606 406201 497670 406265
rect 497826 406201 497890 406265
rect 497906 406201 497970 406265
rect 497986 406201 498050 406265
rect 498066 406201 498130 406265
rect 498146 406201 498210 406265
rect 498226 406201 498290 406265
rect 498306 406201 498370 406265
rect 497126 405482 497190 405546
rect 497206 405482 497270 405546
rect 497286 405482 497350 405546
rect 497366 405482 497430 405546
rect 497446 405482 497510 405546
rect 497526 405482 497590 405546
rect 497606 405482 497670 405546
rect 497826 405482 497890 405546
rect 497906 405482 497970 405546
rect 497986 405482 498050 405546
rect 498066 405482 498130 405546
rect 498146 405482 498210 405546
rect 498226 405482 498290 405546
rect 498306 405482 498370 405546
rect 497126 404763 497190 404827
rect 497206 404763 497270 404827
rect 497286 404763 497350 404827
rect 497366 404763 497430 404827
rect 497446 404763 497510 404827
rect 497526 404763 497590 404827
rect 497606 404763 497670 404827
rect 497826 404763 497890 404827
rect 497906 404763 497970 404827
rect 497986 404763 498050 404827
rect 498066 404763 498130 404827
rect 498146 404763 498210 404827
rect 498226 404763 498290 404827
rect 498306 404763 498370 404827
rect 497126 404044 497190 404108
rect 497206 404044 497270 404108
rect 497286 404044 497350 404108
rect 497366 404044 497430 404108
rect 497446 404044 497510 404108
rect 497526 404044 497590 404108
rect 497606 404044 497670 404108
rect 497826 404044 497890 404108
rect 497906 404044 497970 404108
rect 497986 404044 498050 404108
rect 498066 404044 498130 404108
rect 498146 404044 498210 404108
rect 498226 404044 498290 404108
rect 498306 404044 498370 404108
rect 497126 403325 497190 403389
rect 497206 403325 497270 403389
rect 497286 403325 497350 403389
rect 497366 403325 497430 403389
rect 497446 403325 497510 403389
rect 497526 403325 497590 403389
rect 497606 403325 497670 403389
rect 497826 403325 497890 403389
rect 497906 403325 497970 403389
rect 497986 403325 498050 403389
rect 498066 403325 498130 403389
rect 498146 403325 498210 403389
rect 498226 403325 498290 403389
rect 498306 403325 498370 403389
rect 497126 402606 497190 402670
rect 497206 402606 497270 402670
rect 497286 402606 497350 402670
rect 497366 402606 497430 402670
rect 497446 402606 497510 402670
rect 497526 402606 497590 402670
rect 497606 402606 497670 402670
rect 497826 402606 497890 402670
rect 497906 402606 497970 402670
rect 497986 402606 498050 402670
rect 498066 402606 498130 402670
rect 498146 402606 498210 402670
rect 498226 402606 498290 402670
rect 498306 402606 498370 402670
rect 497126 401887 497190 401951
rect 497206 401887 497270 401951
rect 497286 401887 497350 401951
rect 497366 401887 497430 401951
rect 497446 401887 497510 401951
rect 497526 401887 497590 401951
rect 497606 401887 497670 401951
rect 497826 401887 497890 401951
rect 497906 401887 497970 401951
rect 497986 401887 498050 401951
rect 498066 401887 498130 401951
rect 498146 401887 498210 401951
rect 498226 401887 498290 401951
rect 498306 401887 498370 401951
rect 500886 405809 500950 405873
rect 500966 405809 501030 405873
rect 501046 405809 501110 405873
rect 501126 405809 501190 405873
rect 501206 405809 501270 405873
rect 501286 405809 501350 405873
rect 501366 405809 501430 405873
rect 501586 405809 501650 405873
rect 501666 405809 501730 405873
rect 501746 405809 501810 405873
rect 501826 405809 501890 405873
rect 501906 405809 501970 405873
rect 501986 405809 502050 405873
rect 502066 405809 502130 405873
rect 500886 405090 500950 405154
rect 500966 405090 501030 405154
rect 501046 405090 501110 405154
rect 501126 405090 501190 405154
rect 501206 405090 501270 405154
rect 501286 405090 501350 405154
rect 501366 405090 501430 405154
rect 501586 405090 501650 405154
rect 501666 405090 501730 405154
rect 501746 405090 501810 405154
rect 501826 405090 501890 405154
rect 501906 405090 501970 405154
rect 501986 405090 502050 405154
rect 502066 405090 502130 405154
rect 500886 404371 500950 404435
rect 500966 404371 501030 404435
rect 501046 404371 501110 404435
rect 501126 404371 501190 404435
rect 501206 404371 501270 404435
rect 501286 404371 501350 404435
rect 501366 404371 501430 404435
rect 501586 404371 501650 404435
rect 501666 404371 501730 404435
rect 501746 404371 501810 404435
rect 501826 404371 501890 404435
rect 501906 404371 501970 404435
rect 501986 404371 502050 404435
rect 502066 404371 502130 404435
rect 500886 403652 500950 403716
rect 500966 403652 501030 403716
rect 501046 403652 501110 403716
rect 501126 403652 501190 403716
rect 501206 403652 501270 403716
rect 501286 403652 501350 403716
rect 501366 403652 501430 403716
rect 501586 403652 501650 403716
rect 501666 403652 501730 403716
rect 501746 403652 501810 403716
rect 501826 403652 501890 403716
rect 501906 403652 501970 403716
rect 501986 403652 502050 403716
rect 502066 403652 502130 403716
rect 500886 402933 500950 402997
rect 500966 402933 501030 402997
rect 501046 402933 501110 402997
rect 501126 402933 501190 402997
rect 501206 402933 501270 402997
rect 501286 402933 501350 402997
rect 501366 402933 501430 402997
rect 501586 402933 501650 402997
rect 501666 402933 501730 402997
rect 501746 402933 501810 402997
rect 501826 402933 501890 402997
rect 501906 402933 501970 402997
rect 501986 402933 502050 402997
rect 502066 402933 502130 402997
rect 500886 402214 500950 402278
rect 500966 402214 501030 402278
rect 501046 402214 501110 402278
rect 501126 402214 501190 402278
rect 501206 402214 501270 402278
rect 501286 402214 501350 402278
rect 501366 402214 501430 402278
rect 501586 402214 501650 402278
rect 501666 402214 501730 402278
rect 501746 402214 501810 402278
rect 501826 402214 501890 402278
rect 501906 402214 501970 402278
rect 501986 402214 502050 402278
rect 502066 402214 502130 402278
rect 494766 401516 494830 401560
rect 494766 401496 494770 401516
rect 494770 401496 494826 401516
rect 494826 401496 494830 401516
rect 498218 401490 498282 401554
rect 500886 401495 500950 401559
rect 500966 401495 501030 401559
rect 501046 401495 501110 401559
rect 501126 401495 501190 401559
rect 501206 401495 501270 401559
rect 501286 401495 501350 401559
rect 501366 401495 501430 401559
rect 501586 401495 501650 401559
rect 501666 401495 501730 401559
rect 501746 401495 501810 401559
rect 501826 401495 501890 401559
rect 501906 401495 501970 401559
rect 501986 401495 502050 401559
rect 502066 401495 502130 401559
rect 494766 401460 494770 401480
rect 494770 401460 494826 401480
rect 494826 401460 494830 401480
rect 494766 401416 494830 401460
rect 493366 400910 493430 400974
rect 493446 400910 493510 400974
rect 493526 400910 493590 400974
rect 493606 400910 493670 400974
rect 493686 400910 493750 400974
rect 493766 400910 493830 400974
rect 493846 400910 493910 400974
rect 494066 400910 494130 400974
rect 494146 400910 494210 400974
rect 494226 400910 494290 400974
rect 494306 400910 494370 400974
rect 494386 400910 494450 400974
rect 494466 400910 494530 400974
rect 494546 400910 494610 400974
rect 493366 400191 493430 400255
rect 493446 400191 493510 400255
rect 493526 400191 493590 400255
rect 493606 400191 493670 400255
rect 493686 400191 493750 400255
rect 493766 400191 493830 400255
rect 493846 400191 493910 400255
rect 494066 400191 494130 400255
rect 494146 400191 494210 400255
rect 494226 400191 494290 400255
rect 494306 400191 494370 400255
rect 494386 400191 494450 400255
rect 494466 400191 494530 400255
rect 494546 400191 494610 400255
rect 504806 401352 504870 401416
rect 493366 399472 493430 399536
rect 493446 399472 493510 399536
rect 493526 399472 493590 399536
rect 493606 399472 493670 399536
rect 493686 399472 493750 399536
rect 493766 399472 493830 399536
rect 493846 399472 493910 399536
rect 494066 399472 494130 399536
rect 494146 399472 494210 399536
rect 494226 399472 494290 399536
rect 494306 399472 494370 399536
rect 494386 399472 494450 399536
rect 494466 399472 494530 399536
rect 494546 399472 494610 399536
rect 493366 398753 493430 398817
rect 493446 398753 493510 398817
rect 493526 398753 493590 398817
rect 493606 398753 493670 398817
rect 493686 398753 493750 398817
rect 493766 398753 493830 398817
rect 493846 398753 493910 398817
rect 494066 398753 494130 398817
rect 494146 398753 494210 398817
rect 494226 398753 494290 398817
rect 494306 398753 494370 398817
rect 494386 398753 494450 398817
rect 494466 398753 494530 398817
rect 494546 398753 494610 398817
rect 493366 398034 493430 398098
rect 493446 398034 493510 398098
rect 493526 398034 493590 398098
rect 493606 398034 493670 398098
rect 493686 398034 493750 398098
rect 493766 398034 493830 398098
rect 493846 398034 493910 398098
rect 494066 398034 494130 398098
rect 494146 398034 494210 398098
rect 494226 398034 494290 398098
rect 494306 398034 494370 398098
rect 494386 398034 494450 398098
rect 494466 398034 494530 398098
rect 494546 398034 494610 398098
rect 493366 397315 493430 397379
rect 493446 397315 493510 397379
rect 493526 397315 493590 397379
rect 493606 397315 493670 397379
rect 493686 397315 493750 397379
rect 493766 397315 493830 397379
rect 493846 397315 493910 397379
rect 494066 397315 494130 397379
rect 494146 397315 494210 397379
rect 494226 397315 494290 397379
rect 494306 397315 494370 397379
rect 494386 397315 494450 397379
rect 494466 397315 494530 397379
rect 494546 397315 494610 397379
rect 494924 397272 494988 397276
rect 494924 397216 494928 397272
rect 494928 397216 494984 397272
rect 494984 397216 494988 397272
rect 494924 397212 494988 397216
rect 493366 396596 493430 396660
rect 493446 396596 493510 396660
rect 493526 396596 493590 396660
rect 493606 396596 493670 396660
rect 493686 396596 493750 396660
rect 493766 396596 493830 396660
rect 493846 396596 493910 396660
rect 494066 396596 494130 396660
rect 494146 396596 494210 396660
rect 494226 396596 494290 396660
rect 494306 396596 494370 396660
rect 494386 396596 494450 396660
rect 494466 396596 494530 396660
rect 494546 396596 494610 396660
rect 493366 395877 493430 395941
rect 493446 395877 493510 395941
rect 493526 395877 493590 395941
rect 493606 395877 493670 395941
rect 493686 395877 493750 395941
rect 493766 395877 493830 395941
rect 493846 395877 493910 395941
rect 494066 395877 494130 395941
rect 494146 395877 494210 395941
rect 494226 395877 494290 395941
rect 494306 395877 494370 395941
rect 494386 395877 494450 395941
rect 494466 395877 494530 395941
rect 494546 395877 494610 395941
rect 493366 395158 493430 395222
rect 493446 395158 493510 395222
rect 493526 395158 493590 395222
rect 493606 395158 493670 395222
rect 493686 395158 493750 395222
rect 493766 395158 493830 395222
rect 493846 395158 493910 395222
rect 494066 395158 494130 395222
rect 494146 395158 494210 395222
rect 494226 395158 494290 395222
rect 494306 395158 494370 395222
rect 494386 395158 494450 395222
rect 494466 395158 494530 395222
rect 494546 395158 494610 395222
rect 493366 394439 493430 394503
rect 493446 394439 493510 394503
rect 493526 394439 493590 394503
rect 493606 394439 493670 394503
rect 493686 394439 493750 394503
rect 493766 394439 493830 394503
rect 493846 394439 493910 394503
rect 494066 394439 494130 394503
rect 494146 394439 494210 394503
rect 494226 394439 494290 394503
rect 494306 394439 494370 394503
rect 494386 394439 494450 394503
rect 494466 394439 494530 394503
rect 494546 394439 494610 394503
rect 502286 399752 502350 399796
rect 502286 399732 502290 399752
rect 502290 399732 502346 399752
rect 502346 399732 502350 399752
rect 502286 399696 502290 399716
rect 502290 399696 502346 399716
rect 502346 399696 502350 399716
rect 502286 399652 502350 399696
rect 502366 399480 502430 399484
rect 502366 399424 502370 399480
rect 502370 399424 502426 399480
rect 502426 399424 502430 399480
rect 502366 399420 502430 399424
rect 500886 399146 500950 399210
rect 500966 399146 501030 399210
rect 501046 399146 501110 399210
rect 501126 399146 501190 399210
rect 501206 399146 501270 399210
rect 501286 399146 501350 399210
rect 501366 399146 501430 399210
rect 501586 399146 501650 399210
rect 501666 399146 501730 399210
rect 501746 399146 501810 399210
rect 501826 399146 501890 399210
rect 501906 399146 501970 399210
rect 501986 399146 502050 399210
rect 502066 399146 502130 399210
rect 500886 398427 500950 398491
rect 500966 398427 501030 398491
rect 501046 398427 501110 398491
rect 501126 398427 501190 398491
rect 501206 398427 501270 398491
rect 501286 398427 501350 398491
rect 501366 398427 501430 398491
rect 501586 398427 501650 398491
rect 501666 398427 501730 398491
rect 501746 398427 501810 398491
rect 501826 398427 501890 398491
rect 501906 398427 501970 398491
rect 501986 398427 502050 398491
rect 502066 398427 502130 398491
rect 500886 397708 500950 397772
rect 500966 397708 501030 397772
rect 501046 397708 501110 397772
rect 501126 397708 501190 397772
rect 501206 397708 501270 397772
rect 501286 397708 501350 397772
rect 501366 397708 501430 397772
rect 501586 397708 501650 397772
rect 501666 397708 501730 397772
rect 501746 397708 501810 397772
rect 501826 397708 501890 397772
rect 501906 397708 501970 397772
rect 501986 397708 502050 397772
rect 502066 397708 502130 397772
rect 500886 396989 500950 397053
rect 500966 396989 501030 397053
rect 501046 396989 501110 397053
rect 501126 396989 501190 397053
rect 501206 396989 501270 397053
rect 501286 396989 501350 397053
rect 501366 396989 501430 397053
rect 501586 396989 501650 397053
rect 501666 396989 501730 397053
rect 501746 396989 501810 397053
rect 501826 396989 501890 397053
rect 501906 396989 501970 397053
rect 501986 396989 502050 397053
rect 502066 396989 502130 397053
rect 500886 396270 500950 396334
rect 500966 396270 501030 396334
rect 501046 396270 501110 396334
rect 501126 396270 501190 396334
rect 501206 396270 501270 396334
rect 501286 396270 501350 396334
rect 501366 396270 501430 396334
rect 501586 396270 501650 396334
rect 501666 396270 501730 396334
rect 501746 396270 501810 396334
rect 501826 396270 501890 396334
rect 501906 396270 501970 396334
rect 501986 396270 502050 396334
rect 502066 396270 502130 396334
rect 500886 395551 500950 395615
rect 500966 395551 501030 395615
rect 501046 395551 501110 395615
rect 501126 395551 501190 395615
rect 501206 395551 501270 395615
rect 501286 395551 501350 395615
rect 501366 395551 501430 395615
rect 501586 395551 501650 395615
rect 501666 395551 501730 395615
rect 501746 395551 501810 395615
rect 501826 395551 501890 395615
rect 501906 395551 501970 395615
rect 501986 395551 502050 395615
rect 502066 395551 502130 395615
rect 500886 394832 500950 394896
rect 500966 394832 501030 394896
rect 501046 394832 501110 394896
rect 501126 394832 501190 394896
rect 501206 394832 501270 394896
rect 501286 394832 501350 394896
rect 501366 394832 501430 394896
rect 501586 394832 501650 394896
rect 501666 394832 501730 394896
rect 501746 394832 501810 394896
rect 501826 394832 501890 394896
rect 501906 394832 501970 394896
rect 501986 394832 502050 394896
rect 502066 394832 502130 394896
rect 500886 394113 500950 394177
rect 500966 394113 501030 394177
rect 501046 394113 501110 394177
rect 501126 394113 501190 394177
rect 501206 394113 501270 394177
rect 501286 394113 501350 394177
rect 501366 394113 501430 394177
rect 501586 394113 501650 394177
rect 501666 394113 501730 394177
rect 501746 394113 501810 394177
rect 501826 394113 501890 394177
rect 501906 394113 501970 394177
rect 501986 394113 502050 394177
rect 502066 394113 502130 394177
rect 500886 393394 500950 393458
rect 500966 393394 501030 393458
rect 501046 393394 501110 393458
rect 501126 393394 501190 393458
rect 501206 393394 501270 393458
rect 501286 393394 501350 393458
rect 501366 393394 501430 393458
rect 501586 393394 501650 393458
rect 501666 393394 501730 393458
rect 501746 393394 501810 393458
rect 501826 393394 501890 393458
rect 501906 393394 501970 393458
rect 501986 393394 502050 393458
rect 502066 393394 502130 393458
rect 500658 392708 500662 392722
rect 500662 392708 500718 392722
rect 500718 392708 500722 392722
rect 500658 392658 500722 392708
rect 500886 392675 500950 392739
rect 500966 392675 501030 392739
rect 501046 392675 501110 392739
rect 501126 392675 501190 392739
rect 501206 392675 501270 392739
rect 501286 392675 501350 392739
rect 501366 392675 501430 392739
rect 501586 392675 501650 392739
rect 501666 392675 501730 392739
rect 501746 392675 501810 392739
rect 501826 392675 501890 392739
rect 501906 392675 501970 392739
rect 501986 392675 502050 392739
rect 502066 392675 502130 392739
rect 559736 403192 559926 403368
rect 573538 402980 573888 403312
rect 509806 388678 509870 388722
rect 509806 388658 509810 388678
rect 509810 388658 509866 388678
rect 509866 388658 509870 388678
rect 509806 388622 509810 388642
rect 509810 388622 509866 388642
rect 509866 388622 509870 388642
rect 509806 388578 509870 388622
rect 508406 388072 508470 388136
rect 508486 388072 508550 388136
rect 508566 388072 508630 388136
rect 508646 388072 508710 388136
rect 508726 388072 508790 388136
rect 508806 388072 508870 388136
rect 508886 388072 508950 388136
rect 509106 388072 509170 388136
rect 509186 388072 509250 388136
rect 509266 388072 509330 388136
rect 509346 388072 509410 388136
rect 509426 388072 509490 388136
rect 509506 388072 509570 388136
rect 509586 388072 509650 388136
rect 508406 387353 508470 387417
rect 508486 387353 508550 387417
rect 508566 387353 508630 387417
rect 508646 387353 508710 387417
rect 508726 387353 508790 387417
rect 508806 387353 508870 387417
rect 508886 387353 508950 387417
rect 509106 387353 509170 387417
rect 509186 387353 509250 387417
rect 509266 387353 509330 387417
rect 509346 387353 509410 387417
rect 509426 387353 509490 387417
rect 509506 387353 509570 387417
rect 509586 387353 509650 387417
rect 508406 386634 508470 386698
rect 508486 386634 508550 386698
rect 508566 386634 508630 386698
rect 508646 386634 508710 386698
rect 508726 386634 508790 386698
rect 508806 386634 508870 386698
rect 508886 386634 508950 386698
rect 509106 386634 509170 386698
rect 509186 386634 509250 386698
rect 509266 386634 509330 386698
rect 509346 386634 509410 386698
rect 509426 386634 509490 386698
rect 509506 386634 509570 386698
rect 509586 386634 509650 386698
rect 508406 385915 508470 385979
rect 508486 385915 508550 385979
rect 508566 385915 508630 385979
rect 508646 385915 508710 385979
rect 508726 385915 508790 385979
rect 508806 385915 508870 385979
rect 508886 385915 508950 385979
rect 509106 385915 509170 385979
rect 509186 385915 509250 385979
rect 509266 385915 509330 385979
rect 509346 385915 509410 385979
rect 509426 385915 509490 385979
rect 509506 385915 509570 385979
rect 509586 385915 509650 385979
rect 505050 385206 505114 385270
rect 508406 385196 508470 385260
rect 508486 385196 508550 385260
rect 508566 385196 508630 385260
rect 508646 385196 508710 385260
rect 508726 385196 508790 385260
rect 508806 385196 508870 385260
rect 508886 385196 508950 385260
rect 509106 385196 509170 385260
rect 509186 385196 509250 385260
rect 509266 385196 509330 385260
rect 509346 385196 509410 385260
rect 509426 385196 509490 385260
rect 509506 385196 509570 385260
rect 509586 385196 509650 385260
rect 516274 385206 516338 385270
rect 506046 384954 506110 384998
rect 506046 384934 506050 384954
rect 506050 384934 506106 384954
rect 506106 384934 506110 384954
rect 506046 384898 506050 384918
rect 506050 384898 506106 384918
rect 506106 384898 506110 384918
rect 506046 384854 506110 384898
rect 504646 384348 504710 384412
rect 504726 384348 504790 384412
rect 504806 384348 504870 384412
rect 504886 384348 504950 384412
rect 504966 384348 505030 384412
rect 505046 384348 505110 384412
rect 505126 384348 505190 384412
rect 505346 384348 505410 384412
rect 505426 384348 505490 384412
rect 505506 384348 505570 384412
rect 505586 384348 505650 384412
rect 505666 384348 505730 384412
rect 505746 384348 505810 384412
rect 505826 384348 505890 384412
rect 504646 383629 504710 383693
rect 504726 383629 504790 383693
rect 504806 383629 504870 383693
rect 504886 383629 504950 383693
rect 504966 383629 505030 383693
rect 505046 383629 505110 383693
rect 505126 383629 505190 383693
rect 505346 383629 505410 383693
rect 505426 383629 505490 383693
rect 505506 383629 505570 383693
rect 505586 383629 505650 383693
rect 505666 383629 505730 383693
rect 505746 383629 505810 383693
rect 505826 383629 505890 383693
rect 504646 382910 504710 382974
rect 504726 382910 504790 382974
rect 504806 382910 504870 382974
rect 504886 382910 504950 382974
rect 504966 382910 505030 382974
rect 505046 382910 505110 382974
rect 505126 382910 505190 382974
rect 505346 382910 505410 382974
rect 505426 382910 505490 382974
rect 505506 382910 505570 382974
rect 505586 382910 505650 382974
rect 505666 382910 505730 382974
rect 505746 382910 505810 382974
rect 505826 382910 505890 382974
rect 504646 382191 504710 382255
rect 504726 382191 504790 382255
rect 504806 382191 504870 382255
rect 504886 382191 504950 382255
rect 504966 382191 505030 382255
rect 505046 382191 505110 382255
rect 505126 382191 505190 382255
rect 505346 382191 505410 382255
rect 505426 382191 505490 382255
rect 505506 382191 505570 382255
rect 505586 382191 505650 382255
rect 505666 382191 505730 382255
rect 505746 382191 505810 382255
rect 505826 382191 505890 382255
rect 504440 381540 504504 381544
rect 504440 381484 504444 381540
rect 504444 381484 504500 381540
rect 504500 381484 504504 381540
rect 504440 381480 504504 381484
rect 508406 384477 508470 384541
rect 508486 384477 508550 384541
rect 508566 384477 508630 384541
rect 508646 384477 508710 384541
rect 508726 384477 508790 384541
rect 508806 384477 508870 384541
rect 508886 384477 508950 384541
rect 509106 384477 509170 384541
rect 509186 384477 509250 384541
rect 509266 384477 509330 384541
rect 509346 384477 509410 384541
rect 509426 384477 509490 384541
rect 509506 384477 509570 384541
rect 509586 384477 509650 384541
rect 508406 383758 508470 383822
rect 508486 383758 508550 383822
rect 508566 383758 508630 383822
rect 508646 383758 508710 383822
rect 508726 383758 508790 383822
rect 508806 383758 508870 383822
rect 508886 383758 508950 383822
rect 509106 383758 509170 383822
rect 509186 383758 509250 383822
rect 509266 383758 509330 383822
rect 509346 383758 509410 383822
rect 509426 383758 509490 383822
rect 509506 383758 509570 383822
rect 509586 383758 509650 383822
rect 508406 383039 508470 383103
rect 508486 383039 508550 383103
rect 508566 383039 508630 383103
rect 508646 383039 508710 383103
rect 508726 383039 508790 383103
rect 508806 383039 508870 383103
rect 508886 383039 508950 383103
rect 509106 383039 509170 383103
rect 509186 383039 509250 383103
rect 509266 383039 509330 383103
rect 509346 383039 509410 383103
rect 509426 383039 509490 383103
rect 509506 383039 509570 383103
rect 509586 383039 509650 383103
rect 508406 382320 508470 382384
rect 508486 382320 508550 382384
rect 508566 382320 508630 382384
rect 508646 382320 508710 382384
rect 508726 382320 508790 382384
rect 508806 382320 508870 382384
rect 508886 382320 508950 382384
rect 509106 382320 509170 382384
rect 509186 382320 509250 382384
rect 509266 382320 509330 382384
rect 509346 382320 509410 382384
rect 509426 382320 509490 382384
rect 509506 382320 509570 382384
rect 509586 382320 509650 382384
rect 508222 381618 508286 381682
rect 508406 381601 508470 381665
rect 508486 381601 508550 381665
rect 508566 381601 508630 381665
rect 508646 381601 508710 381665
rect 508726 381601 508790 381665
rect 508806 381601 508870 381665
rect 508886 381601 508950 381665
rect 509106 381601 509170 381665
rect 509186 381601 509250 381665
rect 509266 381601 509330 381665
rect 509346 381601 509410 381665
rect 509426 381601 509490 381665
rect 509506 381601 509570 381665
rect 509586 381601 509650 381665
rect 513566 384954 513630 384998
rect 513566 384934 513570 384954
rect 513570 384934 513626 384954
rect 513626 384934 513630 384954
rect 513566 384898 513570 384918
rect 513570 384898 513626 384918
rect 513626 384898 513630 384918
rect 513566 384854 513630 384898
rect 512166 384348 512230 384412
rect 512246 384348 512310 384412
rect 512326 384348 512390 384412
rect 512406 384348 512470 384412
rect 512486 384348 512550 384412
rect 512566 384348 512630 384412
rect 512646 384348 512710 384412
rect 512866 384348 512930 384412
rect 512946 384348 513010 384412
rect 513026 384348 513090 384412
rect 513106 384348 513170 384412
rect 513186 384348 513250 384412
rect 513266 384348 513330 384412
rect 513346 384348 513410 384412
rect 512166 383629 512230 383693
rect 512246 383629 512310 383693
rect 512326 383629 512390 383693
rect 512406 383629 512470 383693
rect 512486 383629 512550 383693
rect 512566 383629 512630 383693
rect 512646 383629 512710 383693
rect 512866 383629 512930 383693
rect 512946 383629 513010 383693
rect 513026 383629 513090 383693
rect 513106 383629 513170 383693
rect 513186 383629 513250 383693
rect 513266 383629 513330 383693
rect 513346 383629 513410 383693
rect 512166 382910 512230 382974
rect 512246 382910 512310 382974
rect 512326 382910 512390 382974
rect 512406 382910 512470 382974
rect 512486 382910 512550 382974
rect 512566 382910 512630 382974
rect 512646 382910 512710 382974
rect 512866 382910 512930 382974
rect 512946 382910 513010 382974
rect 513026 382910 513090 382974
rect 513106 382910 513170 382974
rect 513186 382910 513250 382974
rect 513266 382910 513330 382974
rect 513346 382910 513410 382974
rect 512166 382191 512230 382255
rect 512246 382191 512310 382255
rect 512326 382191 512390 382255
rect 512406 382191 512470 382255
rect 512486 382191 512550 382255
rect 512566 382191 512630 382255
rect 512646 382191 512710 382255
rect 512866 382191 512930 382255
rect 512946 382191 513010 382255
rect 513026 382191 513090 382255
rect 513106 382191 513170 382255
rect 513186 382191 513250 382255
rect 513266 382191 513330 382255
rect 513346 382191 513410 382255
rect 504646 381472 504710 381536
rect 504726 381472 504790 381536
rect 504806 381472 504870 381536
rect 504886 381472 504950 381536
rect 504966 381472 505030 381536
rect 505046 381472 505110 381536
rect 505126 381472 505190 381536
rect 505346 381472 505410 381536
rect 505426 381472 505490 381536
rect 505506 381472 505570 381536
rect 505586 381472 505650 381536
rect 505666 381472 505730 381536
rect 505746 381472 505810 381536
rect 505826 381472 505890 381536
rect 511882 381540 511946 381544
rect 511882 381484 511886 381540
rect 511886 381484 511942 381540
rect 511942 381484 511946 381540
rect 511882 381480 511946 381484
rect 517326 384954 517390 384998
rect 517326 384934 517330 384954
rect 517330 384934 517386 384954
rect 517386 384934 517390 384954
rect 517326 384898 517330 384918
rect 517330 384898 517386 384918
rect 517386 384898 517390 384918
rect 517326 384854 517390 384898
rect 515926 384348 515990 384412
rect 516006 384348 516070 384412
rect 516086 384348 516150 384412
rect 516166 384348 516230 384412
rect 516246 384348 516310 384412
rect 516326 384348 516390 384412
rect 516406 384348 516470 384412
rect 516626 384348 516690 384412
rect 516706 384348 516770 384412
rect 516786 384348 516850 384412
rect 516866 384348 516930 384412
rect 516946 384348 517010 384412
rect 517026 384348 517090 384412
rect 517106 384348 517170 384412
rect 515926 383629 515990 383693
rect 516006 383629 516070 383693
rect 516086 383629 516150 383693
rect 516166 383629 516230 383693
rect 516246 383629 516310 383693
rect 516326 383629 516390 383693
rect 516406 383629 516470 383693
rect 516626 383629 516690 383693
rect 516706 383629 516770 383693
rect 516786 383629 516850 383693
rect 516866 383629 516930 383693
rect 516946 383629 517010 383693
rect 517026 383629 517090 383693
rect 517106 383629 517170 383693
rect 515926 382910 515990 382974
rect 516006 382910 516070 382974
rect 516086 382910 516150 382974
rect 516166 382910 516230 382974
rect 516246 382910 516310 382974
rect 516326 382910 516390 382974
rect 516406 382910 516470 382974
rect 516626 382910 516690 382974
rect 516706 382910 516770 382974
rect 516786 382910 516850 382974
rect 516866 382910 516930 382974
rect 516946 382910 517010 382974
rect 517026 382910 517090 382974
rect 517106 382910 517170 382974
rect 515926 382191 515990 382255
rect 516006 382191 516070 382255
rect 516086 382191 516150 382255
rect 516166 382191 516230 382255
rect 516246 382191 516310 382255
rect 516326 382191 516390 382255
rect 516406 382191 516470 382255
rect 516626 382191 516690 382255
rect 516706 382191 516770 382255
rect 516786 382191 516850 382255
rect 516866 382191 516930 382255
rect 516946 382191 517010 382255
rect 517026 382191 517090 382255
rect 517106 382191 517170 382255
rect 512166 381472 512230 381536
rect 512246 381472 512310 381536
rect 512326 381472 512390 381536
rect 512406 381472 512470 381536
rect 512486 381472 512550 381536
rect 512566 381472 512630 381536
rect 512646 381472 512710 381536
rect 512866 381472 512930 381536
rect 512946 381472 513010 381536
rect 513026 381472 513090 381536
rect 513106 381472 513170 381536
rect 513186 381472 513250 381536
rect 513266 381472 513330 381536
rect 513346 381472 513410 381536
rect 515664 381540 515728 381544
rect 515664 381484 515668 381540
rect 515668 381484 515724 381540
rect 515724 381484 515728 381540
rect 515664 381480 515728 381484
rect 504646 380753 504710 380817
rect 504726 380753 504790 380817
rect 504806 380753 504870 380817
rect 504886 380753 504950 380817
rect 504966 380753 505030 380817
rect 505046 380753 505110 380817
rect 505126 380753 505190 380817
rect 505346 380753 505410 380817
rect 505426 380753 505490 380817
rect 505506 380753 505570 380817
rect 505586 380753 505650 380817
rect 505666 380753 505730 380817
rect 505746 380753 505810 380817
rect 505826 380753 505890 380817
rect 508222 380790 508286 380854
rect 504646 380034 504710 380098
rect 504726 380034 504790 380098
rect 504806 380034 504870 380098
rect 504886 380034 504950 380098
rect 504966 380034 505030 380098
rect 505046 380034 505110 380098
rect 505126 380034 505190 380098
rect 505346 380034 505410 380098
rect 505426 380034 505490 380098
rect 505506 380034 505570 380098
rect 505586 380034 505650 380098
rect 505666 380034 505730 380098
rect 505746 380034 505810 380098
rect 505826 380034 505890 380098
rect 504646 379315 504710 379379
rect 504726 379315 504790 379379
rect 504806 379315 504870 379379
rect 504886 379315 504950 379379
rect 504966 379315 505030 379379
rect 505046 379315 505110 379379
rect 505126 379315 505190 379379
rect 505346 379315 505410 379379
rect 505426 379315 505490 379379
rect 505506 379315 505570 379379
rect 505586 379315 505650 379379
rect 505666 379315 505730 379379
rect 505746 379315 505810 379379
rect 505826 379315 505890 379379
rect 504646 378596 504710 378660
rect 504726 378596 504790 378660
rect 504806 378596 504870 378660
rect 504886 378596 504950 378660
rect 504966 378596 505030 378660
rect 505046 378596 505110 378660
rect 505126 378596 505190 378660
rect 505346 378596 505410 378660
rect 505426 378596 505490 378660
rect 505506 378596 505570 378660
rect 505586 378596 505650 378660
rect 505666 378596 505730 378660
rect 505746 378596 505810 378660
rect 505826 378596 505890 378660
rect 504646 377877 504710 377941
rect 504726 377877 504790 377941
rect 504806 377877 504870 377941
rect 504886 377877 504950 377941
rect 504966 377877 505030 377941
rect 505046 377877 505110 377941
rect 505126 377877 505190 377941
rect 505346 377877 505410 377941
rect 505426 377877 505490 377941
rect 505506 377877 505570 377941
rect 505586 377877 505650 377941
rect 505666 377877 505730 377941
rect 505746 377877 505810 377941
rect 505826 377877 505890 377941
rect 509806 381230 509870 381274
rect 509806 381210 509810 381230
rect 509810 381210 509866 381230
rect 509866 381210 509870 381230
rect 509806 381174 509810 381194
rect 509810 381174 509866 381194
rect 509866 381174 509870 381194
rect 509806 381130 509870 381174
rect 508406 380624 508470 380688
rect 508486 380624 508550 380688
rect 508566 380624 508630 380688
rect 508646 380624 508710 380688
rect 508726 380624 508790 380688
rect 508806 380624 508870 380688
rect 508886 380624 508950 380688
rect 509106 380624 509170 380688
rect 509186 380624 509250 380688
rect 509266 380624 509330 380688
rect 509346 380624 509410 380688
rect 509426 380624 509490 380688
rect 509506 380624 509570 380688
rect 509586 380624 509650 380688
rect 508406 379905 508470 379969
rect 508486 379905 508550 379969
rect 508566 379905 508630 379969
rect 508646 379905 508710 379969
rect 508726 379905 508790 379969
rect 508806 379905 508870 379969
rect 508886 379905 508950 379969
rect 509106 379905 509170 379969
rect 509186 379905 509250 379969
rect 509266 379905 509330 379969
rect 509346 379905 509410 379969
rect 509426 379905 509490 379969
rect 509506 379905 509570 379969
rect 509586 379905 509650 379969
rect 508406 379186 508470 379250
rect 508486 379186 508550 379250
rect 508566 379186 508630 379250
rect 508646 379186 508710 379250
rect 508726 379186 508790 379250
rect 508806 379186 508870 379250
rect 508886 379186 508950 379250
rect 509106 379186 509170 379250
rect 509186 379186 509250 379250
rect 509266 379186 509330 379250
rect 509346 379186 509410 379250
rect 509426 379186 509490 379250
rect 509506 379186 509570 379250
rect 509586 379186 509650 379250
rect 508406 378467 508470 378531
rect 508486 378467 508550 378531
rect 508566 378467 508630 378531
rect 508646 378467 508710 378531
rect 508726 378467 508790 378531
rect 508806 378467 508870 378531
rect 508886 378467 508950 378531
rect 509106 378467 509170 378531
rect 509186 378467 509250 378531
rect 509266 378467 509330 378531
rect 509346 378467 509410 378531
rect 509426 378467 509490 378531
rect 509506 378467 509570 378531
rect 509586 378467 509650 378531
rect 512166 380753 512230 380817
rect 512246 380753 512310 380817
rect 512326 380753 512390 380817
rect 512406 380753 512470 380817
rect 512486 380753 512550 380817
rect 512566 380753 512630 380817
rect 512646 380753 512710 380817
rect 512866 380753 512930 380817
rect 512946 380753 513010 380817
rect 513026 380753 513090 380817
rect 513106 380753 513170 380817
rect 513186 380753 513250 380817
rect 513266 380753 513330 380817
rect 513346 380753 513410 380817
rect 512166 380034 512230 380098
rect 512246 380034 512310 380098
rect 512326 380034 512390 380098
rect 512406 380034 512470 380098
rect 512486 380034 512550 380098
rect 512566 380034 512630 380098
rect 512646 380034 512710 380098
rect 512866 380034 512930 380098
rect 512946 380034 513010 380098
rect 513026 380034 513090 380098
rect 513106 380034 513170 380098
rect 513186 380034 513250 380098
rect 513266 380034 513330 380098
rect 513346 380034 513410 380098
rect 512166 379315 512230 379379
rect 512246 379315 512310 379379
rect 512326 379315 512390 379379
rect 512406 379315 512470 379379
rect 512486 379315 512550 379379
rect 512566 379315 512630 379379
rect 512646 379315 512710 379379
rect 512866 379315 512930 379379
rect 512946 379315 513010 379379
rect 513026 379315 513090 379379
rect 513106 379315 513170 379379
rect 513186 379315 513250 379379
rect 513266 379315 513330 379379
rect 513346 379315 513410 379379
rect 512166 378596 512230 378660
rect 512246 378596 512310 378660
rect 512326 378596 512390 378660
rect 512406 378596 512470 378660
rect 512486 378596 512550 378660
rect 512566 378596 512630 378660
rect 512646 378596 512710 378660
rect 512866 378596 512930 378660
rect 512946 378596 513010 378660
rect 513026 378596 513090 378660
rect 513106 378596 513170 378660
rect 513186 378596 513250 378660
rect 513266 378596 513330 378660
rect 513346 378596 513410 378660
rect 512166 377877 512230 377941
rect 512246 377877 512310 377941
rect 512326 377877 512390 377941
rect 512406 377877 512470 377941
rect 512486 377877 512550 377941
rect 512566 377877 512630 377941
rect 512646 377877 512710 377941
rect 512866 377877 512930 377941
rect 512946 377877 513010 377941
rect 513026 377877 513090 377941
rect 513106 377877 513170 377941
rect 513186 377877 513250 377941
rect 513266 377877 513330 377941
rect 513346 377877 513410 377941
rect 515926 381472 515990 381536
rect 516006 381472 516070 381536
rect 516086 381472 516150 381536
rect 516166 381472 516230 381536
rect 516246 381472 516310 381536
rect 516326 381472 516390 381536
rect 516406 381472 516470 381536
rect 516626 381472 516690 381536
rect 516706 381472 516770 381536
rect 516786 381472 516850 381536
rect 516866 381472 516930 381536
rect 516946 381472 517010 381536
rect 517026 381472 517090 381536
rect 517106 381472 517170 381536
rect 515926 380753 515990 380817
rect 516006 380753 516070 380817
rect 516086 380753 516150 380817
rect 516166 380753 516230 380817
rect 516246 380753 516310 380817
rect 516326 380753 516390 380817
rect 516406 380753 516470 380817
rect 516626 380753 516690 380817
rect 516706 380753 516770 380817
rect 516786 380753 516850 380817
rect 516866 380753 516930 380817
rect 516946 380753 517010 380817
rect 517026 380753 517090 380817
rect 517106 380753 517170 380817
rect 515926 380034 515990 380098
rect 516006 380034 516070 380098
rect 516086 380034 516150 380098
rect 516166 380034 516230 380098
rect 516246 380034 516310 380098
rect 516326 380034 516390 380098
rect 516406 380034 516470 380098
rect 516626 380034 516690 380098
rect 516706 380034 516770 380098
rect 516786 380034 516850 380098
rect 516866 380034 516930 380098
rect 516946 380034 517010 380098
rect 517026 380034 517090 380098
rect 517106 380034 517170 380098
rect 515926 379315 515990 379379
rect 516006 379315 516070 379379
rect 516086 379315 516150 379379
rect 516166 379315 516230 379379
rect 516246 379315 516310 379379
rect 516326 379315 516390 379379
rect 516406 379315 516470 379379
rect 516626 379315 516690 379379
rect 516706 379315 516770 379379
rect 516786 379315 516850 379379
rect 516866 379315 516930 379379
rect 516946 379315 517010 379379
rect 517026 379315 517090 379379
rect 517106 379315 517170 379379
rect 515926 378596 515990 378660
rect 516006 378596 516070 378660
rect 516086 378596 516150 378660
rect 516166 378596 516230 378660
rect 516246 378596 516310 378660
rect 516326 378596 516390 378660
rect 516406 378596 516470 378660
rect 516626 378596 516690 378660
rect 516706 378596 516770 378660
rect 516786 378596 516850 378660
rect 516866 378596 516930 378660
rect 516946 378596 517010 378660
rect 517026 378596 517090 378660
rect 517106 378596 517170 378660
rect 515926 377877 515990 377941
rect 516006 377877 516070 377941
rect 516086 377877 516150 377941
rect 516166 377877 516230 377941
rect 516246 377877 516310 377941
rect 516326 377877 516390 377941
rect 516406 377877 516470 377941
rect 516626 377877 516690 377941
rect 516706 377877 516770 377941
rect 516786 377877 516850 377941
rect 516866 377877 516930 377941
rect 516946 377877 517010 377941
rect 517026 377877 517090 377941
rect 517106 377877 517170 377941
rect 508406 377748 508470 377812
rect 508486 377748 508550 377812
rect 508566 377748 508630 377812
rect 508646 377748 508710 377812
rect 508726 377748 508790 377812
rect 508806 377748 508870 377812
rect 508886 377748 508950 377812
rect 509106 377748 509170 377812
rect 509186 377748 509250 377812
rect 509266 377748 509330 377812
rect 509346 377748 509410 377812
rect 509426 377748 509490 377812
rect 509506 377748 509570 377812
rect 509586 377748 509650 377812
rect 506026 377400 506090 377404
rect 506026 377344 506030 377400
rect 506030 377344 506086 377400
rect 506086 377344 506090 377400
rect 506026 377340 506090 377344
rect 508406 377029 508470 377093
rect 508486 377029 508550 377093
rect 508566 377029 508630 377093
rect 508646 377029 508710 377093
rect 508726 377029 508790 377093
rect 508806 377029 508870 377093
rect 508886 377029 508950 377093
rect 509106 377029 509170 377093
rect 509186 377029 509250 377093
rect 509266 377029 509330 377093
rect 509346 377029 509410 377093
rect 509426 377029 509490 377093
rect 509506 377029 509570 377093
rect 509586 377029 509650 377093
rect 508406 376310 508470 376374
rect 508486 376310 508550 376374
rect 508566 376310 508630 376374
rect 508646 376310 508710 376374
rect 508726 376310 508790 376374
rect 508806 376310 508870 376374
rect 508886 376310 508950 376374
rect 509106 376310 509170 376374
rect 509186 376310 509250 376374
rect 509266 376310 509330 376374
rect 509346 376310 509410 376374
rect 509426 376310 509490 376374
rect 509506 376310 509570 376374
rect 509586 376310 509650 376374
rect 508406 375591 508470 375655
rect 508486 375591 508550 375655
rect 508566 375591 508630 375655
rect 508646 375591 508710 375655
rect 508726 375591 508790 375655
rect 508806 375591 508870 375655
rect 508886 375591 508950 375655
rect 509106 375591 509170 375655
rect 509186 375591 509250 375655
rect 509266 375591 509330 375655
rect 509346 375591 509410 375655
rect 509426 375591 509490 375655
rect 509506 375591 509570 375655
rect 509586 375591 509650 375655
rect 508406 374872 508470 374936
rect 508486 374872 508550 374936
rect 508566 374872 508630 374936
rect 508646 374872 508710 374936
rect 508726 374872 508790 374936
rect 508806 374872 508870 374936
rect 508886 374872 508950 374936
rect 509106 374872 509170 374936
rect 509186 374872 509250 374936
rect 509266 374872 509330 374936
rect 509346 374872 509410 374936
rect 509426 374872 509490 374936
rect 509506 374872 509570 374936
rect 509586 374872 509650 374936
rect 508406 374153 508470 374217
rect 508486 374153 508550 374217
rect 508566 374153 508630 374217
rect 508646 374153 508710 374217
rect 508726 374153 508790 374217
rect 508806 374153 508870 374217
rect 508886 374153 508950 374217
rect 509106 374153 509170 374217
rect 509186 374153 509250 374217
rect 509266 374153 509330 374217
rect 509346 374153 509410 374217
rect 509426 374153 509490 374217
rect 509506 374153 509570 374217
rect 509586 374153 509650 374217
rect 493076 361470 493140 361474
rect 493076 361414 493080 361470
rect 493080 361414 493136 361470
rect 493136 361414 493140 361470
rect 493076 361410 493140 361414
rect 493076 361390 493140 361394
rect 493076 361334 493080 361390
rect 493080 361334 493136 361390
rect 493136 361334 493140 361390
rect 493076 361330 493140 361334
rect 493076 361310 493140 361314
rect 493076 361254 493080 361310
rect 493080 361254 493136 361310
rect 493136 361254 493140 361310
rect 493076 361250 493140 361254
rect 493076 361230 493140 361234
rect 493076 361174 493080 361230
rect 493080 361174 493136 361230
rect 493136 361174 493140 361230
rect 493076 361170 493140 361174
rect 493076 361150 493140 361154
rect 493076 361094 493080 361150
rect 493080 361094 493136 361150
rect 493136 361094 493140 361150
rect 493076 361090 493140 361094
rect 493076 361070 493140 361074
rect 493076 361014 493080 361070
rect 493080 361014 493136 361070
rect 493136 361014 493140 361070
rect 493076 361010 493140 361014
rect 493076 360990 493140 360994
rect 493076 360934 493080 360990
rect 493080 360934 493136 360990
rect 493136 360934 493140 360990
rect 493076 360930 493140 360934
rect 493076 360910 493140 360914
rect 493076 360854 493080 360910
rect 493080 360854 493136 360910
rect 493136 360854 493140 360910
rect 493076 360850 493140 360854
rect 493076 360830 493140 360834
rect 493076 360774 493080 360830
rect 493080 360774 493136 360830
rect 493136 360774 493140 360830
rect 493076 360770 493140 360774
rect 493076 360750 493140 360754
rect 493076 360694 493080 360750
rect 493080 360694 493136 360750
rect 493136 360694 493140 360750
rect 493076 360690 493140 360694
rect 493076 360670 493140 360674
rect 493076 360614 493080 360670
rect 493080 360614 493136 360670
rect 493136 360614 493140 360670
rect 493076 360610 493140 360614
rect 493076 360590 493140 360594
rect 493076 360534 493080 360590
rect 493080 360534 493136 360590
rect 493136 360534 493140 360590
rect 493076 360530 493140 360534
rect 493076 360510 493140 360514
rect 493076 360454 493080 360510
rect 493080 360454 493136 360510
rect 493136 360454 493140 360510
rect 493076 360450 493140 360454
rect 493076 360430 493140 360434
rect 493076 360374 493080 360430
rect 493080 360374 493136 360430
rect 493136 360374 493140 360430
rect 493076 360370 493140 360374
rect 493076 360350 493140 360354
rect 493076 360294 493080 360350
rect 493080 360294 493136 360350
rect 493136 360294 493140 360350
rect 493076 360290 493140 360294
rect 493076 360270 493140 360274
rect 493076 360214 493080 360270
rect 493080 360214 493136 360270
rect 493136 360214 493140 360270
rect 493076 360210 493140 360214
rect 493076 360190 493140 360194
rect 493076 360134 493080 360190
rect 493080 360134 493136 360190
rect 493136 360134 493140 360190
rect 493076 360130 493140 360134
rect 493076 360110 493140 360114
rect 493076 360054 493080 360110
rect 493080 360054 493136 360110
rect 493136 360054 493140 360110
rect 493076 360050 493140 360054
rect 493076 360030 493140 360034
rect 493076 359974 493080 360030
rect 493080 359974 493136 360030
rect 493136 359974 493140 360030
rect 493076 359970 493140 359974
rect 493076 359950 493140 359954
rect 493076 359894 493080 359950
rect 493080 359894 493136 359950
rect 493136 359894 493140 359950
rect 493076 359890 493140 359894
rect 496836 361470 496900 361474
rect 496836 361414 496840 361470
rect 496840 361414 496896 361470
rect 496896 361414 496900 361470
rect 496836 361410 496900 361414
rect 496836 361390 496900 361394
rect 496836 361334 496840 361390
rect 496840 361334 496896 361390
rect 496896 361334 496900 361390
rect 496836 361330 496900 361334
rect 496836 361310 496900 361314
rect 496836 361254 496840 361310
rect 496840 361254 496896 361310
rect 496896 361254 496900 361310
rect 496836 361250 496900 361254
rect 496836 361230 496900 361234
rect 496836 361174 496840 361230
rect 496840 361174 496896 361230
rect 496896 361174 496900 361230
rect 496836 361170 496900 361174
rect 496836 361150 496900 361154
rect 496836 361094 496840 361150
rect 496840 361094 496896 361150
rect 496896 361094 496900 361150
rect 496836 361090 496900 361094
rect 496836 361070 496900 361074
rect 496836 361014 496840 361070
rect 496840 361014 496896 361070
rect 496896 361014 496900 361070
rect 496836 361010 496900 361014
rect 496836 360990 496900 360994
rect 496836 360934 496840 360990
rect 496840 360934 496896 360990
rect 496896 360934 496900 360990
rect 496836 360930 496900 360934
rect 496836 360910 496900 360914
rect 496836 360854 496840 360910
rect 496840 360854 496896 360910
rect 496896 360854 496900 360910
rect 496836 360850 496900 360854
rect 496836 360830 496900 360834
rect 496836 360774 496840 360830
rect 496840 360774 496896 360830
rect 496896 360774 496900 360830
rect 496836 360770 496900 360774
rect 496836 360750 496900 360754
rect 496836 360694 496840 360750
rect 496840 360694 496896 360750
rect 496896 360694 496900 360750
rect 496836 360690 496900 360694
rect 496836 360670 496900 360674
rect 496836 360614 496840 360670
rect 496840 360614 496896 360670
rect 496896 360614 496900 360670
rect 496836 360610 496900 360614
rect 496836 360590 496900 360594
rect 496836 360534 496840 360590
rect 496840 360534 496896 360590
rect 496896 360534 496900 360590
rect 496836 360530 496900 360534
rect 496836 360510 496900 360514
rect 496836 360454 496840 360510
rect 496840 360454 496896 360510
rect 496896 360454 496900 360510
rect 496836 360450 496900 360454
rect 496836 360430 496900 360434
rect 496836 360374 496840 360430
rect 496840 360374 496896 360430
rect 496896 360374 496900 360430
rect 496836 360370 496900 360374
rect 496836 360350 496900 360354
rect 496836 360294 496840 360350
rect 496840 360294 496896 360350
rect 496896 360294 496900 360350
rect 496836 360290 496900 360294
rect 496836 360270 496900 360274
rect 496836 360214 496840 360270
rect 496840 360214 496896 360270
rect 496896 360214 496900 360270
rect 496836 360210 496900 360214
rect 496836 360190 496900 360194
rect 496836 360134 496840 360190
rect 496840 360134 496896 360190
rect 496896 360134 496900 360190
rect 496836 360130 496900 360134
rect 496836 360110 496900 360114
rect 496836 360054 496840 360110
rect 496840 360054 496896 360110
rect 496896 360054 496900 360110
rect 496836 360050 496900 360054
rect 496836 360030 496900 360034
rect 496836 359974 496840 360030
rect 496840 359974 496896 360030
rect 496896 359974 496900 360030
rect 496836 359970 496900 359974
rect 496836 359950 496900 359954
rect 496836 359894 496840 359950
rect 496840 359894 496896 359950
rect 496896 359894 496900 359950
rect 496836 359890 496900 359894
rect 500596 361470 500660 361474
rect 500596 361414 500600 361470
rect 500600 361414 500656 361470
rect 500656 361414 500660 361470
rect 500596 361410 500660 361414
rect 500596 361390 500660 361394
rect 500596 361334 500600 361390
rect 500600 361334 500656 361390
rect 500656 361334 500660 361390
rect 500596 361330 500660 361334
rect 500596 361310 500660 361314
rect 500596 361254 500600 361310
rect 500600 361254 500656 361310
rect 500656 361254 500660 361310
rect 500596 361250 500660 361254
rect 500596 361230 500660 361234
rect 500596 361174 500600 361230
rect 500600 361174 500656 361230
rect 500656 361174 500660 361230
rect 500596 361170 500660 361174
rect 500596 361150 500660 361154
rect 500596 361094 500600 361150
rect 500600 361094 500656 361150
rect 500656 361094 500660 361150
rect 500596 361090 500660 361094
rect 500596 361070 500660 361074
rect 500596 361014 500600 361070
rect 500600 361014 500656 361070
rect 500656 361014 500660 361070
rect 500596 361010 500660 361014
rect 500596 360990 500660 360994
rect 500596 360934 500600 360990
rect 500600 360934 500656 360990
rect 500656 360934 500660 360990
rect 500596 360930 500660 360934
rect 500596 360910 500660 360914
rect 500596 360854 500600 360910
rect 500600 360854 500656 360910
rect 500656 360854 500660 360910
rect 500596 360850 500660 360854
rect 500596 360830 500660 360834
rect 500596 360774 500600 360830
rect 500600 360774 500656 360830
rect 500656 360774 500660 360830
rect 500596 360770 500660 360774
rect 500596 360750 500660 360754
rect 500596 360694 500600 360750
rect 500600 360694 500656 360750
rect 500656 360694 500660 360750
rect 500596 360690 500660 360694
rect 500596 360670 500660 360674
rect 500596 360614 500600 360670
rect 500600 360614 500656 360670
rect 500656 360614 500660 360670
rect 500596 360610 500660 360614
rect 500596 360590 500660 360594
rect 500596 360534 500600 360590
rect 500600 360534 500656 360590
rect 500656 360534 500660 360590
rect 500596 360530 500660 360534
rect 500596 360510 500660 360514
rect 500596 360454 500600 360510
rect 500600 360454 500656 360510
rect 500656 360454 500660 360510
rect 500596 360450 500660 360454
rect 500596 360430 500660 360434
rect 500596 360374 500600 360430
rect 500600 360374 500656 360430
rect 500656 360374 500660 360430
rect 500596 360370 500660 360374
rect 500596 360350 500660 360354
rect 500596 360294 500600 360350
rect 500600 360294 500656 360350
rect 500656 360294 500660 360350
rect 500596 360290 500660 360294
rect 500596 360270 500660 360274
rect 500596 360214 500600 360270
rect 500600 360214 500656 360270
rect 500656 360214 500660 360270
rect 500596 360210 500660 360214
rect 500596 360190 500660 360194
rect 500596 360134 500600 360190
rect 500600 360134 500656 360190
rect 500656 360134 500660 360190
rect 500596 360130 500660 360134
rect 500596 360110 500660 360114
rect 500596 360054 500600 360110
rect 500600 360054 500656 360110
rect 500656 360054 500660 360110
rect 500596 360050 500660 360054
rect 500596 360030 500660 360034
rect 500596 359974 500600 360030
rect 500600 359974 500656 360030
rect 500656 359974 500660 360030
rect 500596 359970 500660 359974
rect 500596 359950 500660 359954
rect 500596 359894 500600 359950
rect 500600 359894 500656 359950
rect 500656 359894 500660 359950
rect 500596 359890 500660 359894
rect 504356 361470 504420 361474
rect 504356 361414 504360 361470
rect 504360 361414 504416 361470
rect 504416 361414 504420 361470
rect 504356 361410 504420 361414
rect 504356 361390 504420 361394
rect 504356 361334 504360 361390
rect 504360 361334 504416 361390
rect 504416 361334 504420 361390
rect 504356 361330 504420 361334
rect 504356 361310 504420 361314
rect 504356 361254 504360 361310
rect 504360 361254 504416 361310
rect 504416 361254 504420 361310
rect 504356 361250 504420 361254
rect 504356 361230 504420 361234
rect 504356 361174 504360 361230
rect 504360 361174 504416 361230
rect 504416 361174 504420 361230
rect 504356 361170 504420 361174
rect 504356 361150 504420 361154
rect 504356 361094 504360 361150
rect 504360 361094 504416 361150
rect 504416 361094 504420 361150
rect 504356 361090 504420 361094
rect 504356 361070 504420 361074
rect 504356 361014 504360 361070
rect 504360 361014 504416 361070
rect 504416 361014 504420 361070
rect 504356 361010 504420 361014
rect 504356 360990 504420 360994
rect 504356 360934 504360 360990
rect 504360 360934 504416 360990
rect 504416 360934 504420 360990
rect 504356 360930 504420 360934
rect 504356 360910 504420 360914
rect 504356 360854 504360 360910
rect 504360 360854 504416 360910
rect 504416 360854 504420 360910
rect 504356 360850 504420 360854
rect 504356 360830 504420 360834
rect 504356 360774 504360 360830
rect 504360 360774 504416 360830
rect 504416 360774 504420 360830
rect 504356 360770 504420 360774
rect 504356 360750 504420 360754
rect 504356 360694 504360 360750
rect 504360 360694 504416 360750
rect 504416 360694 504420 360750
rect 504356 360690 504420 360694
rect 504356 360670 504420 360674
rect 504356 360614 504360 360670
rect 504360 360614 504416 360670
rect 504416 360614 504420 360670
rect 504356 360610 504420 360614
rect 504356 360590 504420 360594
rect 504356 360534 504360 360590
rect 504360 360534 504416 360590
rect 504416 360534 504420 360590
rect 504356 360530 504420 360534
rect 504356 360510 504420 360514
rect 504356 360454 504360 360510
rect 504360 360454 504416 360510
rect 504416 360454 504420 360510
rect 504356 360450 504420 360454
rect 504356 360430 504420 360434
rect 504356 360374 504360 360430
rect 504360 360374 504416 360430
rect 504416 360374 504420 360430
rect 504356 360370 504420 360374
rect 504356 360350 504420 360354
rect 504356 360294 504360 360350
rect 504360 360294 504416 360350
rect 504416 360294 504420 360350
rect 504356 360290 504420 360294
rect 504356 360270 504420 360274
rect 504356 360214 504360 360270
rect 504360 360214 504416 360270
rect 504416 360214 504420 360270
rect 504356 360210 504420 360214
rect 504356 360190 504420 360194
rect 504356 360134 504360 360190
rect 504360 360134 504416 360190
rect 504416 360134 504420 360190
rect 504356 360130 504420 360134
rect 504356 360110 504420 360114
rect 504356 360054 504360 360110
rect 504360 360054 504416 360110
rect 504416 360054 504420 360110
rect 504356 360050 504420 360054
rect 504356 360030 504420 360034
rect 504356 359974 504360 360030
rect 504360 359974 504416 360030
rect 504416 359974 504420 360030
rect 504356 359970 504420 359974
rect 504356 359950 504420 359954
rect 504356 359894 504360 359950
rect 504360 359894 504416 359950
rect 504416 359894 504420 359950
rect 504356 359890 504420 359894
rect 508116 361470 508180 361474
rect 508116 361414 508120 361470
rect 508120 361414 508176 361470
rect 508176 361414 508180 361470
rect 508116 361410 508180 361414
rect 508116 361390 508180 361394
rect 508116 361334 508120 361390
rect 508120 361334 508176 361390
rect 508176 361334 508180 361390
rect 508116 361330 508180 361334
rect 508116 361310 508180 361314
rect 508116 361254 508120 361310
rect 508120 361254 508176 361310
rect 508176 361254 508180 361310
rect 508116 361250 508180 361254
rect 508116 361230 508180 361234
rect 508116 361174 508120 361230
rect 508120 361174 508176 361230
rect 508176 361174 508180 361230
rect 508116 361170 508180 361174
rect 508116 361150 508180 361154
rect 508116 361094 508120 361150
rect 508120 361094 508176 361150
rect 508176 361094 508180 361150
rect 508116 361090 508180 361094
rect 508116 361070 508180 361074
rect 508116 361014 508120 361070
rect 508120 361014 508176 361070
rect 508176 361014 508180 361070
rect 508116 361010 508180 361014
rect 508116 360990 508180 360994
rect 508116 360934 508120 360990
rect 508120 360934 508176 360990
rect 508176 360934 508180 360990
rect 508116 360930 508180 360934
rect 508116 360910 508180 360914
rect 508116 360854 508120 360910
rect 508120 360854 508176 360910
rect 508176 360854 508180 360910
rect 508116 360850 508180 360854
rect 508116 360830 508180 360834
rect 508116 360774 508120 360830
rect 508120 360774 508176 360830
rect 508176 360774 508180 360830
rect 508116 360770 508180 360774
rect 508116 360750 508180 360754
rect 508116 360694 508120 360750
rect 508120 360694 508176 360750
rect 508176 360694 508180 360750
rect 508116 360690 508180 360694
rect 508116 360670 508180 360674
rect 508116 360614 508120 360670
rect 508120 360614 508176 360670
rect 508176 360614 508180 360670
rect 508116 360610 508180 360614
rect 508116 360590 508180 360594
rect 508116 360534 508120 360590
rect 508120 360534 508176 360590
rect 508176 360534 508180 360590
rect 508116 360530 508180 360534
rect 508116 360510 508180 360514
rect 508116 360454 508120 360510
rect 508120 360454 508176 360510
rect 508176 360454 508180 360510
rect 508116 360450 508180 360454
rect 508116 360430 508180 360434
rect 508116 360374 508120 360430
rect 508120 360374 508176 360430
rect 508176 360374 508180 360430
rect 508116 360370 508180 360374
rect 508116 360350 508180 360354
rect 508116 360294 508120 360350
rect 508120 360294 508176 360350
rect 508176 360294 508180 360350
rect 508116 360290 508180 360294
rect 508116 360270 508180 360274
rect 508116 360214 508120 360270
rect 508120 360214 508176 360270
rect 508176 360214 508180 360270
rect 508116 360210 508180 360214
rect 508116 360190 508180 360194
rect 508116 360134 508120 360190
rect 508120 360134 508176 360190
rect 508176 360134 508180 360190
rect 508116 360130 508180 360134
rect 508116 360110 508180 360114
rect 508116 360054 508120 360110
rect 508120 360054 508176 360110
rect 508176 360054 508180 360110
rect 508116 360050 508180 360054
rect 508116 360030 508180 360034
rect 508116 359974 508120 360030
rect 508120 359974 508176 360030
rect 508176 359974 508180 360030
rect 508116 359970 508180 359974
rect 508116 359950 508180 359954
rect 508116 359894 508120 359950
rect 508120 359894 508176 359950
rect 508176 359894 508180 359950
rect 508116 359890 508180 359894
rect 511876 361470 511940 361474
rect 511876 361414 511880 361470
rect 511880 361414 511936 361470
rect 511936 361414 511940 361470
rect 511876 361410 511940 361414
rect 511876 361390 511940 361394
rect 511876 361334 511880 361390
rect 511880 361334 511936 361390
rect 511936 361334 511940 361390
rect 511876 361330 511940 361334
rect 511876 361310 511940 361314
rect 511876 361254 511880 361310
rect 511880 361254 511936 361310
rect 511936 361254 511940 361310
rect 511876 361250 511940 361254
rect 511876 361230 511940 361234
rect 511876 361174 511880 361230
rect 511880 361174 511936 361230
rect 511936 361174 511940 361230
rect 511876 361170 511940 361174
rect 511876 361150 511940 361154
rect 511876 361094 511880 361150
rect 511880 361094 511936 361150
rect 511936 361094 511940 361150
rect 511876 361090 511940 361094
rect 511876 361070 511940 361074
rect 511876 361014 511880 361070
rect 511880 361014 511936 361070
rect 511936 361014 511940 361070
rect 511876 361010 511940 361014
rect 511876 360990 511940 360994
rect 511876 360934 511880 360990
rect 511880 360934 511936 360990
rect 511936 360934 511940 360990
rect 511876 360930 511940 360934
rect 511876 360910 511940 360914
rect 511876 360854 511880 360910
rect 511880 360854 511936 360910
rect 511936 360854 511940 360910
rect 511876 360850 511940 360854
rect 511876 360830 511940 360834
rect 511876 360774 511880 360830
rect 511880 360774 511936 360830
rect 511936 360774 511940 360830
rect 511876 360770 511940 360774
rect 511876 360750 511940 360754
rect 511876 360694 511880 360750
rect 511880 360694 511936 360750
rect 511936 360694 511940 360750
rect 511876 360690 511940 360694
rect 511876 360670 511940 360674
rect 511876 360614 511880 360670
rect 511880 360614 511936 360670
rect 511936 360614 511940 360670
rect 511876 360610 511940 360614
rect 511876 360590 511940 360594
rect 511876 360534 511880 360590
rect 511880 360534 511936 360590
rect 511936 360534 511940 360590
rect 511876 360530 511940 360534
rect 511876 360510 511940 360514
rect 511876 360454 511880 360510
rect 511880 360454 511936 360510
rect 511936 360454 511940 360510
rect 511876 360450 511940 360454
rect 511876 360430 511940 360434
rect 511876 360374 511880 360430
rect 511880 360374 511936 360430
rect 511936 360374 511940 360430
rect 511876 360370 511940 360374
rect 511876 360350 511940 360354
rect 511876 360294 511880 360350
rect 511880 360294 511936 360350
rect 511936 360294 511940 360350
rect 511876 360290 511940 360294
rect 511876 360270 511940 360274
rect 511876 360214 511880 360270
rect 511880 360214 511936 360270
rect 511936 360214 511940 360270
rect 511876 360210 511940 360214
rect 511876 360190 511940 360194
rect 511876 360134 511880 360190
rect 511880 360134 511936 360190
rect 511936 360134 511940 360190
rect 511876 360130 511940 360134
rect 511876 360110 511940 360114
rect 511876 360054 511880 360110
rect 511880 360054 511936 360110
rect 511936 360054 511940 360110
rect 511876 360050 511940 360054
rect 511876 360030 511940 360034
rect 511876 359974 511880 360030
rect 511880 359974 511936 360030
rect 511936 359974 511940 360030
rect 511876 359970 511940 359974
rect 511876 359950 511940 359954
rect 511876 359894 511880 359950
rect 511880 359894 511936 359950
rect 511936 359894 511940 359950
rect 511876 359890 511940 359894
rect 515636 361470 515700 361474
rect 515636 361414 515640 361470
rect 515640 361414 515696 361470
rect 515696 361414 515700 361470
rect 515636 361410 515700 361414
rect 515636 361390 515700 361394
rect 515636 361334 515640 361390
rect 515640 361334 515696 361390
rect 515696 361334 515700 361390
rect 515636 361330 515700 361334
rect 515636 361310 515700 361314
rect 515636 361254 515640 361310
rect 515640 361254 515696 361310
rect 515696 361254 515700 361310
rect 515636 361250 515700 361254
rect 515636 361230 515700 361234
rect 515636 361174 515640 361230
rect 515640 361174 515696 361230
rect 515696 361174 515700 361230
rect 515636 361170 515700 361174
rect 515636 361150 515700 361154
rect 515636 361094 515640 361150
rect 515640 361094 515696 361150
rect 515696 361094 515700 361150
rect 515636 361090 515700 361094
rect 515636 361070 515700 361074
rect 515636 361014 515640 361070
rect 515640 361014 515696 361070
rect 515696 361014 515700 361070
rect 515636 361010 515700 361014
rect 515636 360990 515700 360994
rect 515636 360934 515640 360990
rect 515640 360934 515696 360990
rect 515696 360934 515700 360990
rect 515636 360930 515700 360934
rect 515636 360910 515700 360914
rect 515636 360854 515640 360910
rect 515640 360854 515696 360910
rect 515696 360854 515700 360910
rect 515636 360850 515700 360854
rect 515636 360830 515700 360834
rect 515636 360774 515640 360830
rect 515640 360774 515696 360830
rect 515696 360774 515700 360830
rect 515636 360770 515700 360774
rect 515636 360750 515700 360754
rect 515636 360694 515640 360750
rect 515640 360694 515696 360750
rect 515696 360694 515700 360750
rect 515636 360690 515700 360694
rect 515636 360670 515700 360674
rect 515636 360614 515640 360670
rect 515640 360614 515696 360670
rect 515696 360614 515700 360670
rect 515636 360610 515700 360614
rect 515636 360590 515700 360594
rect 515636 360534 515640 360590
rect 515640 360534 515696 360590
rect 515696 360534 515700 360590
rect 515636 360530 515700 360534
rect 515636 360510 515700 360514
rect 515636 360454 515640 360510
rect 515640 360454 515696 360510
rect 515696 360454 515700 360510
rect 515636 360450 515700 360454
rect 515636 360430 515700 360434
rect 515636 360374 515640 360430
rect 515640 360374 515696 360430
rect 515696 360374 515700 360430
rect 515636 360370 515700 360374
rect 515636 360350 515700 360354
rect 515636 360294 515640 360350
rect 515640 360294 515696 360350
rect 515696 360294 515700 360350
rect 515636 360290 515700 360294
rect 515636 360270 515700 360274
rect 515636 360214 515640 360270
rect 515640 360214 515696 360270
rect 515696 360214 515700 360270
rect 515636 360210 515700 360214
rect 515636 360190 515700 360194
rect 515636 360134 515640 360190
rect 515640 360134 515696 360190
rect 515696 360134 515700 360190
rect 515636 360130 515700 360134
rect 515636 360110 515700 360114
rect 515636 360054 515640 360110
rect 515640 360054 515696 360110
rect 515696 360054 515700 360110
rect 515636 360050 515700 360054
rect 515636 360030 515700 360034
rect 515636 359974 515640 360030
rect 515640 359974 515696 360030
rect 515696 359974 515700 360030
rect 515636 359970 515700 359974
rect 515636 359950 515700 359954
rect 515636 359894 515640 359950
rect 515640 359894 515696 359950
rect 515696 359894 515700 359950
rect 515636 359890 515700 359894
rect 519396 361470 519460 361474
rect 519396 361414 519400 361470
rect 519400 361414 519456 361470
rect 519456 361414 519460 361470
rect 519396 361410 519460 361414
rect 519396 361390 519460 361394
rect 519396 361334 519400 361390
rect 519400 361334 519456 361390
rect 519456 361334 519460 361390
rect 519396 361330 519460 361334
rect 519396 361310 519460 361314
rect 519396 361254 519400 361310
rect 519400 361254 519456 361310
rect 519456 361254 519460 361310
rect 519396 361250 519460 361254
rect 519396 361230 519460 361234
rect 519396 361174 519400 361230
rect 519400 361174 519456 361230
rect 519456 361174 519460 361230
rect 519396 361170 519460 361174
rect 519396 361150 519460 361154
rect 519396 361094 519400 361150
rect 519400 361094 519456 361150
rect 519456 361094 519460 361150
rect 519396 361090 519460 361094
rect 519396 361070 519460 361074
rect 519396 361014 519400 361070
rect 519400 361014 519456 361070
rect 519456 361014 519460 361070
rect 519396 361010 519460 361014
rect 519396 360990 519460 360994
rect 519396 360934 519400 360990
rect 519400 360934 519456 360990
rect 519456 360934 519460 360990
rect 519396 360930 519460 360934
rect 519396 360910 519460 360914
rect 519396 360854 519400 360910
rect 519400 360854 519456 360910
rect 519456 360854 519460 360910
rect 519396 360850 519460 360854
rect 519396 360830 519460 360834
rect 519396 360774 519400 360830
rect 519400 360774 519456 360830
rect 519456 360774 519460 360830
rect 519396 360770 519460 360774
rect 519396 360750 519460 360754
rect 519396 360694 519400 360750
rect 519400 360694 519456 360750
rect 519456 360694 519460 360750
rect 519396 360690 519460 360694
rect 519396 360670 519460 360674
rect 519396 360614 519400 360670
rect 519400 360614 519456 360670
rect 519456 360614 519460 360670
rect 519396 360610 519460 360614
rect 519396 360590 519460 360594
rect 519396 360534 519400 360590
rect 519400 360534 519456 360590
rect 519456 360534 519460 360590
rect 519396 360530 519460 360534
rect 519396 360510 519460 360514
rect 519396 360454 519400 360510
rect 519400 360454 519456 360510
rect 519456 360454 519460 360510
rect 519396 360450 519460 360454
rect 519396 360430 519460 360434
rect 519396 360374 519400 360430
rect 519400 360374 519456 360430
rect 519456 360374 519460 360430
rect 519396 360370 519460 360374
rect 519396 360350 519460 360354
rect 519396 360294 519400 360350
rect 519400 360294 519456 360350
rect 519456 360294 519460 360350
rect 519396 360290 519460 360294
rect 519396 360270 519460 360274
rect 519396 360214 519400 360270
rect 519400 360214 519456 360270
rect 519456 360214 519460 360270
rect 519396 360210 519460 360214
rect 519396 360190 519460 360194
rect 519396 360134 519400 360190
rect 519400 360134 519456 360190
rect 519456 360134 519460 360190
rect 519396 360130 519460 360134
rect 519396 360110 519460 360114
rect 519396 360054 519400 360110
rect 519400 360054 519456 360110
rect 519456 360054 519460 360110
rect 519396 360050 519460 360054
rect 519396 360030 519460 360034
rect 519396 359974 519400 360030
rect 519400 359974 519456 360030
rect 519456 359974 519460 360030
rect 519396 359970 519460 359974
rect 519396 359950 519460 359954
rect 519396 359894 519400 359950
rect 519400 359894 519456 359950
rect 519456 359894 519460 359950
rect 519396 359890 519460 359894
rect 523156 361470 523220 361474
rect 523156 361414 523160 361470
rect 523160 361414 523216 361470
rect 523216 361414 523220 361470
rect 523156 361410 523220 361414
rect 523156 361390 523220 361394
rect 523156 361334 523160 361390
rect 523160 361334 523216 361390
rect 523216 361334 523220 361390
rect 523156 361330 523220 361334
rect 523156 361310 523220 361314
rect 523156 361254 523160 361310
rect 523160 361254 523216 361310
rect 523216 361254 523220 361310
rect 523156 361250 523220 361254
rect 523156 361230 523220 361234
rect 523156 361174 523160 361230
rect 523160 361174 523216 361230
rect 523216 361174 523220 361230
rect 523156 361170 523220 361174
rect 523156 361150 523220 361154
rect 523156 361094 523160 361150
rect 523160 361094 523216 361150
rect 523216 361094 523220 361150
rect 523156 361090 523220 361094
rect 523156 361070 523220 361074
rect 523156 361014 523160 361070
rect 523160 361014 523216 361070
rect 523216 361014 523220 361070
rect 523156 361010 523220 361014
rect 523156 360990 523220 360994
rect 523156 360934 523160 360990
rect 523160 360934 523216 360990
rect 523216 360934 523220 360990
rect 523156 360930 523220 360934
rect 523156 360910 523220 360914
rect 523156 360854 523160 360910
rect 523160 360854 523216 360910
rect 523216 360854 523220 360910
rect 523156 360850 523220 360854
rect 523156 360830 523220 360834
rect 523156 360774 523160 360830
rect 523160 360774 523216 360830
rect 523216 360774 523220 360830
rect 523156 360770 523220 360774
rect 523156 360750 523220 360754
rect 523156 360694 523160 360750
rect 523160 360694 523216 360750
rect 523216 360694 523220 360750
rect 523156 360690 523220 360694
rect 523156 360670 523220 360674
rect 523156 360614 523160 360670
rect 523160 360614 523216 360670
rect 523216 360614 523220 360670
rect 523156 360610 523220 360614
rect 523156 360590 523220 360594
rect 523156 360534 523160 360590
rect 523160 360534 523216 360590
rect 523216 360534 523220 360590
rect 523156 360530 523220 360534
rect 523156 360510 523220 360514
rect 523156 360454 523160 360510
rect 523160 360454 523216 360510
rect 523216 360454 523220 360510
rect 523156 360450 523220 360454
rect 523156 360430 523220 360434
rect 523156 360374 523160 360430
rect 523160 360374 523216 360430
rect 523216 360374 523220 360430
rect 523156 360370 523220 360374
rect 523156 360350 523220 360354
rect 523156 360294 523160 360350
rect 523160 360294 523216 360350
rect 523216 360294 523220 360350
rect 523156 360290 523220 360294
rect 523156 360270 523220 360274
rect 523156 360214 523160 360270
rect 523160 360214 523216 360270
rect 523216 360214 523220 360270
rect 523156 360210 523220 360214
rect 523156 360190 523220 360194
rect 523156 360134 523160 360190
rect 523160 360134 523216 360190
rect 523216 360134 523220 360190
rect 523156 360130 523220 360134
rect 523156 360110 523220 360114
rect 523156 360054 523160 360110
rect 523160 360054 523216 360110
rect 523216 360054 523220 360110
rect 523156 360050 523220 360054
rect 523156 360030 523220 360034
rect 523156 359974 523160 360030
rect 523160 359974 523216 360030
rect 523216 359974 523220 360030
rect 523156 359970 523220 359974
rect 523156 359950 523220 359954
rect 523156 359894 523160 359950
rect 523160 359894 523216 359950
rect 523216 359894 523220 359950
rect 523156 359890 523220 359894
rect 526916 361470 526980 361474
rect 526916 361414 526920 361470
rect 526920 361414 526976 361470
rect 526976 361414 526980 361470
rect 526916 361410 526980 361414
rect 526916 361390 526980 361394
rect 526916 361334 526920 361390
rect 526920 361334 526976 361390
rect 526976 361334 526980 361390
rect 526916 361330 526980 361334
rect 526916 361310 526980 361314
rect 526916 361254 526920 361310
rect 526920 361254 526976 361310
rect 526976 361254 526980 361310
rect 526916 361250 526980 361254
rect 526916 361230 526980 361234
rect 526916 361174 526920 361230
rect 526920 361174 526976 361230
rect 526976 361174 526980 361230
rect 526916 361170 526980 361174
rect 526916 361150 526980 361154
rect 526916 361094 526920 361150
rect 526920 361094 526976 361150
rect 526976 361094 526980 361150
rect 526916 361090 526980 361094
rect 526916 361070 526980 361074
rect 526916 361014 526920 361070
rect 526920 361014 526976 361070
rect 526976 361014 526980 361070
rect 526916 361010 526980 361014
rect 526916 360990 526980 360994
rect 526916 360934 526920 360990
rect 526920 360934 526976 360990
rect 526976 360934 526980 360990
rect 526916 360930 526980 360934
rect 526916 360910 526980 360914
rect 526916 360854 526920 360910
rect 526920 360854 526976 360910
rect 526976 360854 526980 360910
rect 526916 360850 526980 360854
rect 526916 360830 526980 360834
rect 526916 360774 526920 360830
rect 526920 360774 526976 360830
rect 526976 360774 526980 360830
rect 526916 360770 526980 360774
rect 526916 360750 526980 360754
rect 526916 360694 526920 360750
rect 526920 360694 526976 360750
rect 526976 360694 526980 360750
rect 526916 360690 526980 360694
rect 526916 360670 526980 360674
rect 526916 360614 526920 360670
rect 526920 360614 526976 360670
rect 526976 360614 526980 360670
rect 526916 360610 526980 360614
rect 526916 360590 526980 360594
rect 526916 360534 526920 360590
rect 526920 360534 526976 360590
rect 526976 360534 526980 360590
rect 526916 360530 526980 360534
rect 526916 360510 526980 360514
rect 526916 360454 526920 360510
rect 526920 360454 526976 360510
rect 526976 360454 526980 360510
rect 526916 360450 526980 360454
rect 526916 360430 526980 360434
rect 526916 360374 526920 360430
rect 526920 360374 526976 360430
rect 526976 360374 526980 360430
rect 526916 360370 526980 360374
rect 526916 360350 526980 360354
rect 526916 360294 526920 360350
rect 526920 360294 526976 360350
rect 526976 360294 526980 360350
rect 526916 360290 526980 360294
rect 526916 360270 526980 360274
rect 526916 360214 526920 360270
rect 526920 360214 526976 360270
rect 526976 360214 526980 360270
rect 526916 360210 526980 360214
rect 526916 360190 526980 360194
rect 526916 360134 526920 360190
rect 526920 360134 526976 360190
rect 526976 360134 526980 360190
rect 526916 360130 526980 360134
rect 526916 360110 526980 360114
rect 526916 360054 526920 360110
rect 526920 360054 526976 360110
rect 526976 360054 526980 360110
rect 526916 360050 526980 360054
rect 526916 360030 526980 360034
rect 526916 359974 526920 360030
rect 526920 359974 526976 360030
rect 526976 359974 526980 360030
rect 526916 359970 526980 359974
rect 526916 359950 526980 359954
rect 526916 359894 526920 359950
rect 526920 359894 526976 359950
rect 526976 359894 526980 359950
rect 526916 359890 526980 359894
rect 530676 361470 530740 361474
rect 530676 361414 530680 361470
rect 530680 361414 530736 361470
rect 530736 361414 530740 361470
rect 530676 361410 530740 361414
rect 530676 361390 530740 361394
rect 530676 361334 530680 361390
rect 530680 361334 530736 361390
rect 530736 361334 530740 361390
rect 530676 361330 530740 361334
rect 530676 361310 530740 361314
rect 530676 361254 530680 361310
rect 530680 361254 530736 361310
rect 530736 361254 530740 361310
rect 530676 361250 530740 361254
rect 530676 361230 530740 361234
rect 530676 361174 530680 361230
rect 530680 361174 530736 361230
rect 530736 361174 530740 361230
rect 530676 361170 530740 361174
rect 530676 361150 530740 361154
rect 530676 361094 530680 361150
rect 530680 361094 530736 361150
rect 530736 361094 530740 361150
rect 530676 361090 530740 361094
rect 530676 361070 530740 361074
rect 530676 361014 530680 361070
rect 530680 361014 530736 361070
rect 530736 361014 530740 361070
rect 530676 361010 530740 361014
rect 530676 360990 530740 360994
rect 530676 360934 530680 360990
rect 530680 360934 530736 360990
rect 530736 360934 530740 360990
rect 530676 360930 530740 360934
rect 530676 360910 530740 360914
rect 530676 360854 530680 360910
rect 530680 360854 530736 360910
rect 530736 360854 530740 360910
rect 530676 360850 530740 360854
rect 530676 360830 530740 360834
rect 530676 360774 530680 360830
rect 530680 360774 530736 360830
rect 530736 360774 530740 360830
rect 530676 360770 530740 360774
rect 530676 360750 530740 360754
rect 530676 360694 530680 360750
rect 530680 360694 530736 360750
rect 530736 360694 530740 360750
rect 530676 360690 530740 360694
rect 530676 360670 530740 360674
rect 530676 360614 530680 360670
rect 530680 360614 530736 360670
rect 530736 360614 530740 360670
rect 530676 360610 530740 360614
rect 530676 360590 530740 360594
rect 530676 360534 530680 360590
rect 530680 360534 530736 360590
rect 530736 360534 530740 360590
rect 530676 360530 530740 360534
rect 530676 360510 530740 360514
rect 530676 360454 530680 360510
rect 530680 360454 530736 360510
rect 530736 360454 530740 360510
rect 530676 360450 530740 360454
rect 530676 360430 530740 360434
rect 530676 360374 530680 360430
rect 530680 360374 530736 360430
rect 530736 360374 530740 360430
rect 530676 360370 530740 360374
rect 530676 360350 530740 360354
rect 530676 360294 530680 360350
rect 530680 360294 530736 360350
rect 530736 360294 530740 360350
rect 530676 360290 530740 360294
rect 530676 360270 530740 360274
rect 530676 360214 530680 360270
rect 530680 360214 530736 360270
rect 530736 360214 530740 360270
rect 530676 360210 530740 360214
rect 530676 360190 530740 360194
rect 530676 360134 530680 360190
rect 530680 360134 530736 360190
rect 530736 360134 530740 360190
rect 530676 360130 530740 360134
rect 530676 360110 530740 360114
rect 530676 360054 530680 360110
rect 530680 360054 530736 360110
rect 530736 360054 530740 360110
rect 530676 360050 530740 360054
rect 530676 360030 530740 360034
rect 530676 359974 530680 360030
rect 530680 359974 530736 360030
rect 530736 359974 530740 360030
rect 530676 359970 530740 359974
rect 530676 359950 530740 359954
rect 530676 359894 530680 359950
rect 530680 359894 530736 359950
rect 530736 359894 530740 359950
rect 530676 359890 530740 359894
rect 534436 361470 534500 361474
rect 534436 361414 534440 361470
rect 534440 361414 534496 361470
rect 534496 361414 534500 361470
rect 534436 361410 534500 361414
rect 534436 361390 534500 361394
rect 534436 361334 534440 361390
rect 534440 361334 534496 361390
rect 534496 361334 534500 361390
rect 534436 361330 534500 361334
rect 534436 361310 534500 361314
rect 534436 361254 534440 361310
rect 534440 361254 534496 361310
rect 534496 361254 534500 361310
rect 534436 361250 534500 361254
rect 534436 361230 534500 361234
rect 534436 361174 534440 361230
rect 534440 361174 534496 361230
rect 534496 361174 534500 361230
rect 534436 361170 534500 361174
rect 534436 361150 534500 361154
rect 534436 361094 534440 361150
rect 534440 361094 534496 361150
rect 534496 361094 534500 361150
rect 534436 361090 534500 361094
rect 534436 361070 534500 361074
rect 534436 361014 534440 361070
rect 534440 361014 534496 361070
rect 534496 361014 534500 361070
rect 534436 361010 534500 361014
rect 534436 360990 534500 360994
rect 534436 360934 534440 360990
rect 534440 360934 534496 360990
rect 534496 360934 534500 360990
rect 534436 360930 534500 360934
rect 534436 360910 534500 360914
rect 534436 360854 534440 360910
rect 534440 360854 534496 360910
rect 534496 360854 534500 360910
rect 534436 360850 534500 360854
rect 534436 360830 534500 360834
rect 534436 360774 534440 360830
rect 534440 360774 534496 360830
rect 534496 360774 534500 360830
rect 534436 360770 534500 360774
rect 534436 360750 534500 360754
rect 534436 360694 534440 360750
rect 534440 360694 534496 360750
rect 534496 360694 534500 360750
rect 534436 360690 534500 360694
rect 534436 360670 534500 360674
rect 534436 360614 534440 360670
rect 534440 360614 534496 360670
rect 534496 360614 534500 360670
rect 534436 360610 534500 360614
rect 534436 360590 534500 360594
rect 534436 360534 534440 360590
rect 534440 360534 534496 360590
rect 534496 360534 534500 360590
rect 534436 360530 534500 360534
rect 534436 360510 534500 360514
rect 534436 360454 534440 360510
rect 534440 360454 534496 360510
rect 534496 360454 534500 360510
rect 534436 360450 534500 360454
rect 534436 360430 534500 360434
rect 534436 360374 534440 360430
rect 534440 360374 534496 360430
rect 534496 360374 534500 360430
rect 534436 360370 534500 360374
rect 534436 360350 534500 360354
rect 534436 360294 534440 360350
rect 534440 360294 534496 360350
rect 534496 360294 534500 360350
rect 534436 360290 534500 360294
rect 534436 360270 534500 360274
rect 534436 360214 534440 360270
rect 534440 360214 534496 360270
rect 534496 360214 534500 360270
rect 534436 360210 534500 360214
rect 534436 360190 534500 360194
rect 534436 360134 534440 360190
rect 534440 360134 534496 360190
rect 534496 360134 534500 360190
rect 534436 360130 534500 360134
rect 534436 360110 534500 360114
rect 534436 360054 534440 360110
rect 534440 360054 534496 360110
rect 534496 360054 534500 360110
rect 534436 360050 534500 360054
rect 534436 360030 534500 360034
rect 534436 359974 534440 360030
rect 534440 359974 534496 360030
rect 534496 359974 534500 360030
rect 534436 359970 534500 359974
rect 534436 359950 534500 359954
rect 534436 359894 534440 359950
rect 534440 359894 534496 359950
rect 534496 359894 534500 359950
rect 534436 359890 534500 359894
rect 491196 359022 491260 359026
rect 491196 358966 491200 359022
rect 491200 358966 491256 359022
rect 491256 358966 491260 359022
rect 491196 358962 491260 358966
rect 491196 358942 491260 358946
rect 491196 358886 491200 358942
rect 491200 358886 491256 358942
rect 491256 358886 491260 358942
rect 491196 358882 491260 358886
rect 491196 358862 491260 358866
rect 491196 358806 491200 358862
rect 491200 358806 491256 358862
rect 491256 358806 491260 358862
rect 491196 358802 491260 358806
rect 491196 358782 491260 358786
rect 491196 358726 491200 358782
rect 491200 358726 491256 358782
rect 491256 358726 491260 358782
rect 491196 358722 491260 358726
rect 491196 358702 491260 358706
rect 491196 358646 491200 358702
rect 491200 358646 491256 358702
rect 491256 358646 491260 358702
rect 491196 358642 491260 358646
rect 491196 358622 491260 358626
rect 491196 358566 491200 358622
rect 491200 358566 491256 358622
rect 491256 358566 491260 358622
rect 491196 358562 491260 358566
rect 491196 358542 491260 358546
rect 491196 358486 491200 358542
rect 491200 358486 491256 358542
rect 491256 358486 491260 358542
rect 491196 358482 491260 358486
rect 491196 358462 491260 358466
rect 491196 358406 491200 358462
rect 491200 358406 491256 358462
rect 491256 358406 491260 358462
rect 491196 358402 491260 358406
rect 491196 358382 491260 358386
rect 491196 358326 491200 358382
rect 491200 358326 491256 358382
rect 491256 358326 491260 358382
rect 491196 358322 491260 358326
rect 491196 358302 491260 358306
rect 491196 358246 491200 358302
rect 491200 358246 491256 358302
rect 491256 358246 491260 358302
rect 491196 358242 491260 358246
rect 491196 358222 491260 358226
rect 491196 358166 491200 358222
rect 491200 358166 491256 358222
rect 491256 358166 491260 358222
rect 491196 358162 491260 358166
rect 491196 358142 491260 358146
rect 491196 358086 491200 358142
rect 491200 358086 491256 358142
rect 491256 358086 491260 358142
rect 491196 358082 491260 358086
rect 491196 358062 491260 358066
rect 491196 358006 491200 358062
rect 491200 358006 491256 358062
rect 491256 358006 491260 358062
rect 491196 358002 491260 358006
rect 491196 357982 491260 357986
rect 491196 357926 491200 357982
rect 491200 357926 491256 357982
rect 491256 357926 491260 357982
rect 491196 357922 491260 357926
rect 491196 357902 491260 357906
rect 491196 357846 491200 357902
rect 491200 357846 491256 357902
rect 491256 357846 491260 357902
rect 491196 357842 491260 357846
rect 491196 357822 491260 357826
rect 491196 357766 491200 357822
rect 491200 357766 491256 357822
rect 491256 357766 491260 357822
rect 491196 357762 491260 357766
rect 491196 357742 491260 357746
rect 491196 357686 491200 357742
rect 491200 357686 491256 357742
rect 491256 357686 491260 357742
rect 491196 357682 491260 357686
rect 491196 357662 491260 357666
rect 491196 357606 491200 357662
rect 491200 357606 491256 357662
rect 491256 357606 491260 357662
rect 491196 357602 491260 357606
rect 491196 357582 491260 357586
rect 491196 357526 491200 357582
rect 491200 357526 491256 357582
rect 491256 357526 491260 357582
rect 491196 357522 491260 357526
rect 491196 357502 491260 357506
rect 491196 357446 491200 357502
rect 491200 357446 491256 357502
rect 491256 357446 491260 357502
rect 491196 357442 491260 357446
rect 494956 359022 495020 359026
rect 494956 358966 494960 359022
rect 494960 358966 495016 359022
rect 495016 358966 495020 359022
rect 494956 358962 495020 358966
rect 494956 358942 495020 358946
rect 494956 358886 494960 358942
rect 494960 358886 495016 358942
rect 495016 358886 495020 358942
rect 494956 358882 495020 358886
rect 494956 358862 495020 358866
rect 494956 358806 494960 358862
rect 494960 358806 495016 358862
rect 495016 358806 495020 358862
rect 494956 358802 495020 358806
rect 494956 358782 495020 358786
rect 494956 358726 494960 358782
rect 494960 358726 495016 358782
rect 495016 358726 495020 358782
rect 494956 358722 495020 358726
rect 494956 358702 495020 358706
rect 494956 358646 494960 358702
rect 494960 358646 495016 358702
rect 495016 358646 495020 358702
rect 494956 358642 495020 358646
rect 494956 358622 495020 358626
rect 494956 358566 494960 358622
rect 494960 358566 495016 358622
rect 495016 358566 495020 358622
rect 494956 358562 495020 358566
rect 494956 358542 495020 358546
rect 494956 358486 494960 358542
rect 494960 358486 495016 358542
rect 495016 358486 495020 358542
rect 494956 358482 495020 358486
rect 494956 358462 495020 358466
rect 494956 358406 494960 358462
rect 494960 358406 495016 358462
rect 495016 358406 495020 358462
rect 494956 358402 495020 358406
rect 494956 358382 495020 358386
rect 494956 358326 494960 358382
rect 494960 358326 495016 358382
rect 495016 358326 495020 358382
rect 494956 358322 495020 358326
rect 494956 358302 495020 358306
rect 494956 358246 494960 358302
rect 494960 358246 495016 358302
rect 495016 358246 495020 358302
rect 494956 358242 495020 358246
rect 494956 358222 495020 358226
rect 494956 358166 494960 358222
rect 494960 358166 495016 358222
rect 495016 358166 495020 358222
rect 494956 358162 495020 358166
rect 494956 358142 495020 358146
rect 494956 358086 494960 358142
rect 494960 358086 495016 358142
rect 495016 358086 495020 358142
rect 494956 358082 495020 358086
rect 494956 358062 495020 358066
rect 494956 358006 494960 358062
rect 494960 358006 495016 358062
rect 495016 358006 495020 358062
rect 494956 358002 495020 358006
rect 494956 357982 495020 357986
rect 494956 357926 494960 357982
rect 494960 357926 495016 357982
rect 495016 357926 495020 357982
rect 494956 357922 495020 357926
rect 494956 357902 495020 357906
rect 494956 357846 494960 357902
rect 494960 357846 495016 357902
rect 495016 357846 495020 357902
rect 494956 357842 495020 357846
rect 494956 357822 495020 357826
rect 494956 357766 494960 357822
rect 494960 357766 495016 357822
rect 495016 357766 495020 357822
rect 494956 357762 495020 357766
rect 494956 357742 495020 357746
rect 494956 357686 494960 357742
rect 494960 357686 495016 357742
rect 495016 357686 495020 357742
rect 494956 357682 495020 357686
rect 494956 357662 495020 357666
rect 494956 357606 494960 357662
rect 494960 357606 495016 357662
rect 495016 357606 495020 357662
rect 494956 357602 495020 357606
rect 494956 357582 495020 357586
rect 494956 357526 494960 357582
rect 494960 357526 495016 357582
rect 495016 357526 495020 357582
rect 494956 357522 495020 357526
rect 494956 357502 495020 357506
rect 494956 357446 494960 357502
rect 494960 357446 495016 357502
rect 495016 357446 495020 357502
rect 494956 357442 495020 357446
rect 498716 359022 498780 359026
rect 498716 358966 498720 359022
rect 498720 358966 498776 359022
rect 498776 358966 498780 359022
rect 498716 358962 498780 358966
rect 498716 358942 498780 358946
rect 498716 358886 498720 358942
rect 498720 358886 498776 358942
rect 498776 358886 498780 358942
rect 498716 358882 498780 358886
rect 498716 358862 498780 358866
rect 498716 358806 498720 358862
rect 498720 358806 498776 358862
rect 498776 358806 498780 358862
rect 498716 358802 498780 358806
rect 498716 358782 498780 358786
rect 498716 358726 498720 358782
rect 498720 358726 498776 358782
rect 498776 358726 498780 358782
rect 498716 358722 498780 358726
rect 498716 358702 498780 358706
rect 498716 358646 498720 358702
rect 498720 358646 498776 358702
rect 498776 358646 498780 358702
rect 498716 358642 498780 358646
rect 498716 358622 498780 358626
rect 498716 358566 498720 358622
rect 498720 358566 498776 358622
rect 498776 358566 498780 358622
rect 498716 358562 498780 358566
rect 498716 358542 498780 358546
rect 498716 358486 498720 358542
rect 498720 358486 498776 358542
rect 498776 358486 498780 358542
rect 498716 358482 498780 358486
rect 498716 358462 498780 358466
rect 498716 358406 498720 358462
rect 498720 358406 498776 358462
rect 498776 358406 498780 358462
rect 498716 358402 498780 358406
rect 498716 358382 498780 358386
rect 498716 358326 498720 358382
rect 498720 358326 498776 358382
rect 498776 358326 498780 358382
rect 498716 358322 498780 358326
rect 498716 358302 498780 358306
rect 498716 358246 498720 358302
rect 498720 358246 498776 358302
rect 498776 358246 498780 358302
rect 498716 358242 498780 358246
rect 498716 358222 498780 358226
rect 498716 358166 498720 358222
rect 498720 358166 498776 358222
rect 498776 358166 498780 358222
rect 498716 358162 498780 358166
rect 498716 358142 498780 358146
rect 498716 358086 498720 358142
rect 498720 358086 498776 358142
rect 498776 358086 498780 358142
rect 498716 358082 498780 358086
rect 498716 358062 498780 358066
rect 498716 358006 498720 358062
rect 498720 358006 498776 358062
rect 498776 358006 498780 358062
rect 498716 358002 498780 358006
rect 498716 357982 498780 357986
rect 498716 357926 498720 357982
rect 498720 357926 498776 357982
rect 498776 357926 498780 357982
rect 498716 357922 498780 357926
rect 498716 357902 498780 357906
rect 498716 357846 498720 357902
rect 498720 357846 498776 357902
rect 498776 357846 498780 357902
rect 498716 357842 498780 357846
rect 498716 357822 498780 357826
rect 498716 357766 498720 357822
rect 498720 357766 498776 357822
rect 498776 357766 498780 357822
rect 498716 357762 498780 357766
rect 498716 357742 498780 357746
rect 498716 357686 498720 357742
rect 498720 357686 498776 357742
rect 498776 357686 498780 357742
rect 498716 357682 498780 357686
rect 498716 357662 498780 357666
rect 498716 357606 498720 357662
rect 498720 357606 498776 357662
rect 498776 357606 498780 357662
rect 498716 357602 498780 357606
rect 498716 357582 498780 357586
rect 498716 357526 498720 357582
rect 498720 357526 498776 357582
rect 498776 357526 498780 357582
rect 498716 357522 498780 357526
rect 498716 357502 498780 357506
rect 498716 357446 498720 357502
rect 498720 357446 498776 357502
rect 498776 357446 498780 357502
rect 498716 357442 498780 357446
rect 502476 359022 502540 359026
rect 502476 358966 502480 359022
rect 502480 358966 502536 359022
rect 502536 358966 502540 359022
rect 502476 358962 502540 358966
rect 502476 358942 502540 358946
rect 502476 358886 502480 358942
rect 502480 358886 502536 358942
rect 502536 358886 502540 358942
rect 502476 358882 502540 358886
rect 502476 358862 502540 358866
rect 502476 358806 502480 358862
rect 502480 358806 502536 358862
rect 502536 358806 502540 358862
rect 502476 358802 502540 358806
rect 502476 358782 502540 358786
rect 502476 358726 502480 358782
rect 502480 358726 502536 358782
rect 502536 358726 502540 358782
rect 502476 358722 502540 358726
rect 502476 358702 502540 358706
rect 502476 358646 502480 358702
rect 502480 358646 502536 358702
rect 502536 358646 502540 358702
rect 502476 358642 502540 358646
rect 502476 358622 502540 358626
rect 502476 358566 502480 358622
rect 502480 358566 502536 358622
rect 502536 358566 502540 358622
rect 502476 358562 502540 358566
rect 502476 358542 502540 358546
rect 502476 358486 502480 358542
rect 502480 358486 502536 358542
rect 502536 358486 502540 358542
rect 502476 358482 502540 358486
rect 502476 358462 502540 358466
rect 502476 358406 502480 358462
rect 502480 358406 502536 358462
rect 502536 358406 502540 358462
rect 502476 358402 502540 358406
rect 502476 358382 502540 358386
rect 502476 358326 502480 358382
rect 502480 358326 502536 358382
rect 502536 358326 502540 358382
rect 502476 358322 502540 358326
rect 502476 358302 502540 358306
rect 502476 358246 502480 358302
rect 502480 358246 502536 358302
rect 502536 358246 502540 358302
rect 502476 358242 502540 358246
rect 502476 358222 502540 358226
rect 502476 358166 502480 358222
rect 502480 358166 502536 358222
rect 502536 358166 502540 358222
rect 502476 358162 502540 358166
rect 502476 358142 502540 358146
rect 502476 358086 502480 358142
rect 502480 358086 502536 358142
rect 502536 358086 502540 358142
rect 502476 358082 502540 358086
rect 502476 358062 502540 358066
rect 502476 358006 502480 358062
rect 502480 358006 502536 358062
rect 502536 358006 502540 358062
rect 502476 358002 502540 358006
rect 502476 357982 502540 357986
rect 502476 357926 502480 357982
rect 502480 357926 502536 357982
rect 502536 357926 502540 357982
rect 502476 357922 502540 357926
rect 502476 357902 502540 357906
rect 502476 357846 502480 357902
rect 502480 357846 502536 357902
rect 502536 357846 502540 357902
rect 502476 357842 502540 357846
rect 502476 357822 502540 357826
rect 502476 357766 502480 357822
rect 502480 357766 502536 357822
rect 502536 357766 502540 357822
rect 502476 357762 502540 357766
rect 502476 357742 502540 357746
rect 502476 357686 502480 357742
rect 502480 357686 502536 357742
rect 502536 357686 502540 357742
rect 502476 357682 502540 357686
rect 502476 357662 502540 357666
rect 502476 357606 502480 357662
rect 502480 357606 502536 357662
rect 502536 357606 502540 357662
rect 502476 357602 502540 357606
rect 502476 357582 502540 357586
rect 502476 357526 502480 357582
rect 502480 357526 502536 357582
rect 502536 357526 502540 357582
rect 502476 357522 502540 357526
rect 502476 357502 502540 357506
rect 502476 357446 502480 357502
rect 502480 357446 502536 357502
rect 502536 357446 502540 357502
rect 502476 357442 502540 357446
rect 506236 359022 506300 359026
rect 506236 358966 506240 359022
rect 506240 358966 506296 359022
rect 506296 358966 506300 359022
rect 506236 358962 506300 358966
rect 506236 358942 506300 358946
rect 506236 358886 506240 358942
rect 506240 358886 506296 358942
rect 506296 358886 506300 358942
rect 506236 358882 506300 358886
rect 506236 358862 506300 358866
rect 506236 358806 506240 358862
rect 506240 358806 506296 358862
rect 506296 358806 506300 358862
rect 506236 358802 506300 358806
rect 506236 358782 506300 358786
rect 506236 358726 506240 358782
rect 506240 358726 506296 358782
rect 506296 358726 506300 358782
rect 506236 358722 506300 358726
rect 506236 358702 506300 358706
rect 506236 358646 506240 358702
rect 506240 358646 506296 358702
rect 506296 358646 506300 358702
rect 506236 358642 506300 358646
rect 506236 358622 506300 358626
rect 506236 358566 506240 358622
rect 506240 358566 506296 358622
rect 506296 358566 506300 358622
rect 506236 358562 506300 358566
rect 506236 358542 506300 358546
rect 506236 358486 506240 358542
rect 506240 358486 506296 358542
rect 506296 358486 506300 358542
rect 506236 358482 506300 358486
rect 506236 358462 506300 358466
rect 506236 358406 506240 358462
rect 506240 358406 506296 358462
rect 506296 358406 506300 358462
rect 506236 358402 506300 358406
rect 506236 358382 506300 358386
rect 506236 358326 506240 358382
rect 506240 358326 506296 358382
rect 506296 358326 506300 358382
rect 506236 358322 506300 358326
rect 506236 358302 506300 358306
rect 506236 358246 506240 358302
rect 506240 358246 506296 358302
rect 506296 358246 506300 358302
rect 506236 358242 506300 358246
rect 506236 358222 506300 358226
rect 506236 358166 506240 358222
rect 506240 358166 506296 358222
rect 506296 358166 506300 358222
rect 506236 358162 506300 358166
rect 506236 358142 506300 358146
rect 506236 358086 506240 358142
rect 506240 358086 506296 358142
rect 506296 358086 506300 358142
rect 506236 358082 506300 358086
rect 506236 358062 506300 358066
rect 506236 358006 506240 358062
rect 506240 358006 506296 358062
rect 506296 358006 506300 358062
rect 506236 358002 506300 358006
rect 506236 357982 506300 357986
rect 506236 357926 506240 357982
rect 506240 357926 506296 357982
rect 506296 357926 506300 357982
rect 506236 357922 506300 357926
rect 506236 357902 506300 357906
rect 506236 357846 506240 357902
rect 506240 357846 506296 357902
rect 506296 357846 506300 357902
rect 506236 357842 506300 357846
rect 506236 357822 506300 357826
rect 506236 357766 506240 357822
rect 506240 357766 506296 357822
rect 506296 357766 506300 357822
rect 506236 357762 506300 357766
rect 506236 357742 506300 357746
rect 506236 357686 506240 357742
rect 506240 357686 506296 357742
rect 506296 357686 506300 357742
rect 506236 357682 506300 357686
rect 506236 357662 506300 357666
rect 506236 357606 506240 357662
rect 506240 357606 506296 357662
rect 506296 357606 506300 357662
rect 506236 357602 506300 357606
rect 506236 357582 506300 357586
rect 506236 357526 506240 357582
rect 506240 357526 506296 357582
rect 506296 357526 506300 357582
rect 506236 357522 506300 357526
rect 506236 357502 506300 357506
rect 506236 357446 506240 357502
rect 506240 357446 506296 357502
rect 506296 357446 506300 357502
rect 506236 357442 506300 357446
rect 509996 359022 510060 359026
rect 509996 358966 510000 359022
rect 510000 358966 510056 359022
rect 510056 358966 510060 359022
rect 509996 358962 510060 358966
rect 509996 358942 510060 358946
rect 509996 358886 510000 358942
rect 510000 358886 510056 358942
rect 510056 358886 510060 358942
rect 509996 358882 510060 358886
rect 509996 358862 510060 358866
rect 509996 358806 510000 358862
rect 510000 358806 510056 358862
rect 510056 358806 510060 358862
rect 509996 358802 510060 358806
rect 509996 358782 510060 358786
rect 509996 358726 510000 358782
rect 510000 358726 510056 358782
rect 510056 358726 510060 358782
rect 509996 358722 510060 358726
rect 509996 358702 510060 358706
rect 509996 358646 510000 358702
rect 510000 358646 510056 358702
rect 510056 358646 510060 358702
rect 509996 358642 510060 358646
rect 509996 358622 510060 358626
rect 509996 358566 510000 358622
rect 510000 358566 510056 358622
rect 510056 358566 510060 358622
rect 509996 358562 510060 358566
rect 509996 358542 510060 358546
rect 509996 358486 510000 358542
rect 510000 358486 510056 358542
rect 510056 358486 510060 358542
rect 509996 358482 510060 358486
rect 509996 358462 510060 358466
rect 509996 358406 510000 358462
rect 510000 358406 510056 358462
rect 510056 358406 510060 358462
rect 509996 358402 510060 358406
rect 509996 358382 510060 358386
rect 509996 358326 510000 358382
rect 510000 358326 510056 358382
rect 510056 358326 510060 358382
rect 509996 358322 510060 358326
rect 509996 358302 510060 358306
rect 509996 358246 510000 358302
rect 510000 358246 510056 358302
rect 510056 358246 510060 358302
rect 509996 358242 510060 358246
rect 509996 358222 510060 358226
rect 509996 358166 510000 358222
rect 510000 358166 510056 358222
rect 510056 358166 510060 358222
rect 509996 358162 510060 358166
rect 509996 358142 510060 358146
rect 509996 358086 510000 358142
rect 510000 358086 510056 358142
rect 510056 358086 510060 358142
rect 509996 358082 510060 358086
rect 509996 358062 510060 358066
rect 509996 358006 510000 358062
rect 510000 358006 510056 358062
rect 510056 358006 510060 358062
rect 509996 358002 510060 358006
rect 509996 357982 510060 357986
rect 509996 357926 510000 357982
rect 510000 357926 510056 357982
rect 510056 357926 510060 357982
rect 509996 357922 510060 357926
rect 509996 357902 510060 357906
rect 509996 357846 510000 357902
rect 510000 357846 510056 357902
rect 510056 357846 510060 357902
rect 509996 357842 510060 357846
rect 509996 357822 510060 357826
rect 509996 357766 510000 357822
rect 510000 357766 510056 357822
rect 510056 357766 510060 357822
rect 509996 357762 510060 357766
rect 509996 357742 510060 357746
rect 509996 357686 510000 357742
rect 510000 357686 510056 357742
rect 510056 357686 510060 357742
rect 509996 357682 510060 357686
rect 509996 357662 510060 357666
rect 509996 357606 510000 357662
rect 510000 357606 510056 357662
rect 510056 357606 510060 357662
rect 509996 357602 510060 357606
rect 509996 357582 510060 357586
rect 509996 357526 510000 357582
rect 510000 357526 510056 357582
rect 510056 357526 510060 357582
rect 509996 357522 510060 357526
rect 509996 357502 510060 357506
rect 509996 357446 510000 357502
rect 510000 357446 510056 357502
rect 510056 357446 510060 357502
rect 509996 357442 510060 357446
rect 513756 359022 513820 359026
rect 513756 358966 513760 359022
rect 513760 358966 513816 359022
rect 513816 358966 513820 359022
rect 513756 358962 513820 358966
rect 513756 358942 513820 358946
rect 513756 358886 513760 358942
rect 513760 358886 513816 358942
rect 513816 358886 513820 358942
rect 513756 358882 513820 358886
rect 513756 358862 513820 358866
rect 513756 358806 513760 358862
rect 513760 358806 513816 358862
rect 513816 358806 513820 358862
rect 513756 358802 513820 358806
rect 513756 358782 513820 358786
rect 513756 358726 513760 358782
rect 513760 358726 513816 358782
rect 513816 358726 513820 358782
rect 513756 358722 513820 358726
rect 513756 358702 513820 358706
rect 513756 358646 513760 358702
rect 513760 358646 513816 358702
rect 513816 358646 513820 358702
rect 513756 358642 513820 358646
rect 513756 358622 513820 358626
rect 513756 358566 513760 358622
rect 513760 358566 513816 358622
rect 513816 358566 513820 358622
rect 513756 358562 513820 358566
rect 513756 358542 513820 358546
rect 513756 358486 513760 358542
rect 513760 358486 513816 358542
rect 513816 358486 513820 358542
rect 513756 358482 513820 358486
rect 513756 358462 513820 358466
rect 513756 358406 513760 358462
rect 513760 358406 513816 358462
rect 513816 358406 513820 358462
rect 513756 358402 513820 358406
rect 513756 358382 513820 358386
rect 513756 358326 513760 358382
rect 513760 358326 513816 358382
rect 513816 358326 513820 358382
rect 513756 358322 513820 358326
rect 513756 358302 513820 358306
rect 513756 358246 513760 358302
rect 513760 358246 513816 358302
rect 513816 358246 513820 358302
rect 513756 358242 513820 358246
rect 513756 358222 513820 358226
rect 513756 358166 513760 358222
rect 513760 358166 513816 358222
rect 513816 358166 513820 358222
rect 513756 358162 513820 358166
rect 513756 358142 513820 358146
rect 513756 358086 513760 358142
rect 513760 358086 513816 358142
rect 513816 358086 513820 358142
rect 513756 358082 513820 358086
rect 513756 358062 513820 358066
rect 513756 358006 513760 358062
rect 513760 358006 513816 358062
rect 513816 358006 513820 358062
rect 513756 358002 513820 358006
rect 513756 357982 513820 357986
rect 513756 357926 513760 357982
rect 513760 357926 513816 357982
rect 513816 357926 513820 357982
rect 513756 357922 513820 357926
rect 513756 357902 513820 357906
rect 513756 357846 513760 357902
rect 513760 357846 513816 357902
rect 513816 357846 513820 357902
rect 513756 357842 513820 357846
rect 513756 357822 513820 357826
rect 513756 357766 513760 357822
rect 513760 357766 513816 357822
rect 513816 357766 513820 357822
rect 513756 357762 513820 357766
rect 513756 357742 513820 357746
rect 513756 357686 513760 357742
rect 513760 357686 513816 357742
rect 513816 357686 513820 357742
rect 513756 357682 513820 357686
rect 513756 357662 513820 357666
rect 513756 357606 513760 357662
rect 513760 357606 513816 357662
rect 513816 357606 513820 357662
rect 513756 357602 513820 357606
rect 513756 357582 513820 357586
rect 513756 357526 513760 357582
rect 513760 357526 513816 357582
rect 513816 357526 513820 357582
rect 513756 357522 513820 357526
rect 513756 357502 513820 357506
rect 513756 357446 513760 357502
rect 513760 357446 513816 357502
rect 513816 357446 513820 357502
rect 513756 357442 513820 357446
rect 517516 359022 517580 359026
rect 517516 358966 517520 359022
rect 517520 358966 517576 359022
rect 517576 358966 517580 359022
rect 517516 358962 517580 358966
rect 517516 358942 517580 358946
rect 517516 358886 517520 358942
rect 517520 358886 517576 358942
rect 517576 358886 517580 358942
rect 517516 358882 517580 358886
rect 517516 358862 517580 358866
rect 517516 358806 517520 358862
rect 517520 358806 517576 358862
rect 517576 358806 517580 358862
rect 517516 358802 517580 358806
rect 517516 358782 517580 358786
rect 517516 358726 517520 358782
rect 517520 358726 517576 358782
rect 517576 358726 517580 358782
rect 517516 358722 517580 358726
rect 517516 358702 517580 358706
rect 517516 358646 517520 358702
rect 517520 358646 517576 358702
rect 517576 358646 517580 358702
rect 517516 358642 517580 358646
rect 517516 358622 517580 358626
rect 517516 358566 517520 358622
rect 517520 358566 517576 358622
rect 517576 358566 517580 358622
rect 517516 358562 517580 358566
rect 517516 358542 517580 358546
rect 517516 358486 517520 358542
rect 517520 358486 517576 358542
rect 517576 358486 517580 358542
rect 517516 358482 517580 358486
rect 517516 358462 517580 358466
rect 517516 358406 517520 358462
rect 517520 358406 517576 358462
rect 517576 358406 517580 358462
rect 517516 358402 517580 358406
rect 517516 358382 517580 358386
rect 517516 358326 517520 358382
rect 517520 358326 517576 358382
rect 517576 358326 517580 358382
rect 517516 358322 517580 358326
rect 517516 358302 517580 358306
rect 517516 358246 517520 358302
rect 517520 358246 517576 358302
rect 517576 358246 517580 358302
rect 517516 358242 517580 358246
rect 517516 358222 517580 358226
rect 517516 358166 517520 358222
rect 517520 358166 517576 358222
rect 517576 358166 517580 358222
rect 517516 358162 517580 358166
rect 517516 358142 517580 358146
rect 517516 358086 517520 358142
rect 517520 358086 517576 358142
rect 517576 358086 517580 358142
rect 517516 358082 517580 358086
rect 517516 358062 517580 358066
rect 517516 358006 517520 358062
rect 517520 358006 517576 358062
rect 517576 358006 517580 358062
rect 517516 358002 517580 358006
rect 517516 357982 517580 357986
rect 517516 357926 517520 357982
rect 517520 357926 517576 357982
rect 517576 357926 517580 357982
rect 517516 357922 517580 357926
rect 517516 357902 517580 357906
rect 517516 357846 517520 357902
rect 517520 357846 517576 357902
rect 517576 357846 517580 357902
rect 517516 357842 517580 357846
rect 517516 357822 517580 357826
rect 517516 357766 517520 357822
rect 517520 357766 517576 357822
rect 517576 357766 517580 357822
rect 517516 357762 517580 357766
rect 517516 357742 517580 357746
rect 517516 357686 517520 357742
rect 517520 357686 517576 357742
rect 517576 357686 517580 357742
rect 517516 357682 517580 357686
rect 517516 357662 517580 357666
rect 517516 357606 517520 357662
rect 517520 357606 517576 357662
rect 517576 357606 517580 357662
rect 517516 357602 517580 357606
rect 517516 357582 517580 357586
rect 517516 357526 517520 357582
rect 517520 357526 517576 357582
rect 517576 357526 517580 357582
rect 517516 357522 517580 357526
rect 517516 357502 517580 357506
rect 517516 357446 517520 357502
rect 517520 357446 517576 357502
rect 517576 357446 517580 357502
rect 517516 357442 517580 357446
rect 521276 359022 521340 359026
rect 521276 358966 521280 359022
rect 521280 358966 521336 359022
rect 521336 358966 521340 359022
rect 521276 358962 521340 358966
rect 521276 358942 521340 358946
rect 521276 358886 521280 358942
rect 521280 358886 521336 358942
rect 521336 358886 521340 358942
rect 521276 358882 521340 358886
rect 521276 358862 521340 358866
rect 521276 358806 521280 358862
rect 521280 358806 521336 358862
rect 521336 358806 521340 358862
rect 521276 358802 521340 358806
rect 521276 358782 521340 358786
rect 521276 358726 521280 358782
rect 521280 358726 521336 358782
rect 521336 358726 521340 358782
rect 521276 358722 521340 358726
rect 521276 358702 521340 358706
rect 521276 358646 521280 358702
rect 521280 358646 521336 358702
rect 521336 358646 521340 358702
rect 521276 358642 521340 358646
rect 521276 358622 521340 358626
rect 521276 358566 521280 358622
rect 521280 358566 521336 358622
rect 521336 358566 521340 358622
rect 521276 358562 521340 358566
rect 521276 358542 521340 358546
rect 521276 358486 521280 358542
rect 521280 358486 521336 358542
rect 521336 358486 521340 358542
rect 521276 358482 521340 358486
rect 521276 358462 521340 358466
rect 521276 358406 521280 358462
rect 521280 358406 521336 358462
rect 521336 358406 521340 358462
rect 521276 358402 521340 358406
rect 521276 358382 521340 358386
rect 521276 358326 521280 358382
rect 521280 358326 521336 358382
rect 521336 358326 521340 358382
rect 521276 358322 521340 358326
rect 521276 358302 521340 358306
rect 521276 358246 521280 358302
rect 521280 358246 521336 358302
rect 521336 358246 521340 358302
rect 521276 358242 521340 358246
rect 521276 358222 521340 358226
rect 521276 358166 521280 358222
rect 521280 358166 521336 358222
rect 521336 358166 521340 358222
rect 521276 358162 521340 358166
rect 521276 358142 521340 358146
rect 521276 358086 521280 358142
rect 521280 358086 521336 358142
rect 521336 358086 521340 358142
rect 521276 358082 521340 358086
rect 521276 358062 521340 358066
rect 521276 358006 521280 358062
rect 521280 358006 521336 358062
rect 521336 358006 521340 358062
rect 521276 358002 521340 358006
rect 521276 357982 521340 357986
rect 521276 357926 521280 357982
rect 521280 357926 521336 357982
rect 521336 357926 521340 357982
rect 521276 357922 521340 357926
rect 521276 357902 521340 357906
rect 521276 357846 521280 357902
rect 521280 357846 521336 357902
rect 521336 357846 521340 357902
rect 521276 357842 521340 357846
rect 521276 357822 521340 357826
rect 521276 357766 521280 357822
rect 521280 357766 521336 357822
rect 521336 357766 521340 357822
rect 521276 357762 521340 357766
rect 521276 357742 521340 357746
rect 521276 357686 521280 357742
rect 521280 357686 521336 357742
rect 521336 357686 521340 357742
rect 521276 357682 521340 357686
rect 521276 357662 521340 357666
rect 521276 357606 521280 357662
rect 521280 357606 521336 357662
rect 521336 357606 521340 357662
rect 521276 357602 521340 357606
rect 521276 357582 521340 357586
rect 521276 357526 521280 357582
rect 521280 357526 521336 357582
rect 521336 357526 521340 357582
rect 521276 357522 521340 357526
rect 521276 357502 521340 357506
rect 521276 357446 521280 357502
rect 521280 357446 521336 357502
rect 521336 357446 521340 357502
rect 521276 357442 521340 357446
rect 525036 359022 525100 359026
rect 525036 358966 525040 359022
rect 525040 358966 525096 359022
rect 525096 358966 525100 359022
rect 525036 358962 525100 358966
rect 525036 358942 525100 358946
rect 525036 358886 525040 358942
rect 525040 358886 525096 358942
rect 525096 358886 525100 358942
rect 525036 358882 525100 358886
rect 525036 358862 525100 358866
rect 525036 358806 525040 358862
rect 525040 358806 525096 358862
rect 525096 358806 525100 358862
rect 525036 358802 525100 358806
rect 525036 358782 525100 358786
rect 525036 358726 525040 358782
rect 525040 358726 525096 358782
rect 525096 358726 525100 358782
rect 525036 358722 525100 358726
rect 525036 358702 525100 358706
rect 525036 358646 525040 358702
rect 525040 358646 525096 358702
rect 525096 358646 525100 358702
rect 525036 358642 525100 358646
rect 525036 358622 525100 358626
rect 525036 358566 525040 358622
rect 525040 358566 525096 358622
rect 525096 358566 525100 358622
rect 525036 358562 525100 358566
rect 525036 358542 525100 358546
rect 525036 358486 525040 358542
rect 525040 358486 525096 358542
rect 525096 358486 525100 358542
rect 525036 358482 525100 358486
rect 525036 358462 525100 358466
rect 525036 358406 525040 358462
rect 525040 358406 525096 358462
rect 525096 358406 525100 358462
rect 525036 358402 525100 358406
rect 525036 358382 525100 358386
rect 525036 358326 525040 358382
rect 525040 358326 525096 358382
rect 525096 358326 525100 358382
rect 525036 358322 525100 358326
rect 525036 358302 525100 358306
rect 525036 358246 525040 358302
rect 525040 358246 525096 358302
rect 525096 358246 525100 358302
rect 525036 358242 525100 358246
rect 525036 358222 525100 358226
rect 525036 358166 525040 358222
rect 525040 358166 525096 358222
rect 525096 358166 525100 358222
rect 525036 358162 525100 358166
rect 525036 358142 525100 358146
rect 525036 358086 525040 358142
rect 525040 358086 525096 358142
rect 525096 358086 525100 358142
rect 525036 358082 525100 358086
rect 525036 358062 525100 358066
rect 525036 358006 525040 358062
rect 525040 358006 525096 358062
rect 525096 358006 525100 358062
rect 525036 358002 525100 358006
rect 525036 357982 525100 357986
rect 525036 357926 525040 357982
rect 525040 357926 525096 357982
rect 525096 357926 525100 357982
rect 525036 357922 525100 357926
rect 525036 357902 525100 357906
rect 525036 357846 525040 357902
rect 525040 357846 525096 357902
rect 525096 357846 525100 357902
rect 525036 357842 525100 357846
rect 525036 357822 525100 357826
rect 525036 357766 525040 357822
rect 525040 357766 525096 357822
rect 525096 357766 525100 357822
rect 525036 357762 525100 357766
rect 525036 357742 525100 357746
rect 525036 357686 525040 357742
rect 525040 357686 525096 357742
rect 525096 357686 525100 357742
rect 525036 357682 525100 357686
rect 525036 357662 525100 357666
rect 525036 357606 525040 357662
rect 525040 357606 525096 357662
rect 525096 357606 525100 357662
rect 525036 357602 525100 357606
rect 525036 357582 525100 357586
rect 525036 357526 525040 357582
rect 525040 357526 525096 357582
rect 525096 357526 525100 357582
rect 525036 357522 525100 357526
rect 525036 357502 525100 357506
rect 525036 357446 525040 357502
rect 525040 357446 525096 357502
rect 525096 357446 525100 357502
rect 525036 357442 525100 357446
rect 528796 359022 528860 359026
rect 528796 358966 528800 359022
rect 528800 358966 528856 359022
rect 528856 358966 528860 359022
rect 528796 358962 528860 358966
rect 528796 358942 528860 358946
rect 528796 358886 528800 358942
rect 528800 358886 528856 358942
rect 528856 358886 528860 358942
rect 528796 358882 528860 358886
rect 528796 358862 528860 358866
rect 528796 358806 528800 358862
rect 528800 358806 528856 358862
rect 528856 358806 528860 358862
rect 528796 358802 528860 358806
rect 528796 358782 528860 358786
rect 528796 358726 528800 358782
rect 528800 358726 528856 358782
rect 528856 358726 528860 358782
rect 528796 358722 528860 358726
rect 528796 358702 528860 358706
rect 528796 358646 528800 358702
rect 528800 358646 528856 358702
rect 528856 358646 528860 358702
rect 528796 358642 528860 358646
rect 528796 358622 528860 358626
rect 528796 358566 528800 358622
rect 528800 358566 528856 358622
rect 528856 358566 528860 358622
rect 528796 358562 528860 358566
rect 528796 358542 528860 358546
rect 528796 358486 528800 358542
rect 528800 358486 528856 358542
rect 528856 358486 528860 358542
rect 528796 358482 528860 358486
rect 528796 358462 528860 358466
rect 528796 358406 528800 358462
rect 528800 358406 528856 358462
rect 528856 358406 528860 358462
rect 528796 358402 528860 358406
rect 528796 358382 528860 358386
rect 528796 358326 528800 358382
rect 528800 358326 528856 358382
rect 528856 358326 528860 358382
rect 528796 358322 528860 358326
rect 528796 358302 528860 358306
rect 528796 358246 528800 358302
rect 528800 358246 528856 358302
rect 528856 358246 528860 358302
rect 528796 358242 528860 358246
rect 528796 358222 528860 358226
rect 528796 358166 528800 358222
rect 528800 358166 528856 358222
rect 528856 358166 528860 358222
rect 528796 358162 528860 358166
rect 528796 358142 528860 358146
rect 528796 358086 528800 358142
rect 528800 358086 528856 358142
rect 528856 358086 528860 358142
rect 528796 358082 528860 358086
rect 528796 358062 528860 358066
rect 528796 358006 528800 358062
rect 528800 358006 528856 358062
rect 528856 358006 528860 358062
rect 528796 358002 528860 358006
rect 528796 357982 528860 357986
rect 528796 357926 528800 357982
rect 528800 357926 528856 357982
rect 528856 357926 528860 357982
rect 528796 357922 528860 357926
rect 528796 357902 528860 357906
rect 528796 357846 528800 357902
rect 528800 357846 528856 357902
rect 528856 357846 528860 357902
rect 528796 357842 528860 357846
rect 528796 357822 528860 357826
rect 528796 357766 528800 357822
rect 528800 357766 528856 357822
rect 528856 357766 528860 357822
rect 528796 357762 528860 357766
rect 528796 357742 528860 357746
rect 528796 357686 528800 357742
rect 528800 357686 528856 357742
rect 528856 357686 528860 357742
rect 528796 357682 528860 357686
rect 528796 357662 528860 357666
rect 528796 357606 528800 357662
rect 528800 357606 528856 357662
rect 528856 357606 528860 357662
rect 528796 357602 528860 357606
rect 528796 357582 528860 357586
rect 528796 357526 528800 357582
rect 528800 357526 528856 357582
rect 528856 357526 528860 357582
rect 528796 357522 528860 357526
rect 528796 357502 528860 357506
rect 528796 357446 528800 357502
rect 528800 357446 528856 357502
rect 528856 357446 528860 357502
rect 528796 357442 528860 357446
rect 532556 359022 532620 359026
rect 532556 358966 532560 359022
rect 532560 358966 532616 359022
rect 532616 358966 532620 359022
rect 532556 358962 532620 358966
rect 532556 358942 532620 358946
rect 532556 358886 532560 358942
rect 532560 358886 532616 358942
rect 532616 358886 532620 358942
rect 532556 358882 532620 358886
rect 532556 358862 532620 358866
rect 532556 358806 532560 358862
rect 532560 358806 532616 358862
rect 532616 358806 532620 358862
rect 532556 358802 532620 358806
rect 532556 358782 532620 358786
rect 532556 358726 532560 358782
rect 532560 358726 532616 358782
rect 532616 358726 532620 358782
rect 532556 358722 532620 358726
rect 532556 358702 532620 358706
rect 532556 358646 532560 358702
rect 532560 358646 532616 358702
rect 532616 358646 532620 358702
rect 532556 358642 532620 358646
rect 532556 358622 532620 358626
rect 532556 358566 532560 358622
rect 532560 358566 532616 358622
rect 532616 358566 532620 358622
rect 532556 358562 532620 358566
rect 532556 358542 532620 358546
rect 532556 358486 532560 358542
rect 532560 358486 532616 358542
rect 532616 358486 532620 358542
rect 532556 358482 532620 358486
rect 532556 358462 532620 358466
rect 532556 358406 532560 358462
rect 532560 358406 532616 358462
rect 532616 358406 532620 358462
rect 532556 358402 532620 358406
rect 532556 358382 532620 358386
rect 532556 358326 532560 358382
rect 532560 358326 532616 358382
rect 532616 358326 532620 358382
rect 532556 358322 532620 358326
rect 532556 358302 532620 358306
rect 532556 358246 532560 358302
rect 532560 358246 532616 358302
rect 532616 358246 532620 358302
rect 532556 358242 532620 358246
rect 532556 358222 532620 358226
rect 532556 358166 532560 358222
rect 532560 358166 532616 358222
rect 532616 358166 532620 358222
rect 532556 358162 532620 358166
rect 532556 358142 532620 358146
rect 532556 358086 532560 358142
rect 532560 358086 532616 358142
rect 532616 358086 532620 358142
rect 532556 358082 532620 358086
rect 532556 358062 532620 358066
rect 532556 358006 532560 358062
rect 532560 358006 532616 358062
rect 532616 358006 532620 358062
rect 532556 358002 532620 358006
rect 532556 357982 532620 357986
rect 532556 357926 532560 357982
rect 532560 357926 532616 357982
rect 532616 357926 532620 357982
rect 532556 357922 532620 357926
rect 532556 357902 532620 357906
rect 532556 357846 532560 357902
rect 532560 357846 532616 357902
rect 532616 357846 532620 357902
rect 532556 357842 532620 357846
rect 532556 357822 532620 357826
rect 532556 357766 532560 357822
rect 532560 357766 532616 357822
rect 532616 357766 532620 357822
rect 532556 357762 532620 357766
rect 532556 357742 532620 357746
rect 532556 357686 532560 357742
rect 532560 357686 532616 357742
rect 532616 357686 532620 357742
rect 532556 357682 532620 357686
rect 532556 357662 532620 357666
rect 532556 357606 532560 357662
rect 532560 357606 532616 357662
rect 532616 357606 532620 357662
rect 532556 357602 532620 357606
rect 532556 357582 532620 357586
rect 532556 357526 532560 357582
rect 532560 357526 532616 357582
rect 532616 357526 532620 357582
rect 532556 357522 532620 357526
rect 532556 357502 532620 357506
rect 532556 357446 532560 357502
rect 532560 357446 532616 357502
rect 532616 357446 532620 357502
rect 532556 357442 532620 357446
rect 536316 359022 536380 359026
rect 536316 358966 536320 359022
rect 536320 358966 536376 359022
rect 536376 358966 536380 359022
rect 536316 358962 536380 358966
rect 536316 358942 536380 358946
rect 536316 358886 536320 358942
rect 536320 358886 536376 358942
rect 536376 358886 536380 358942
rect 536316 358882 536380 358886
rect 536316 358862 536380 358866
rect 536316 358806 536320 358862
rect 536320 358806 536376 358862
rect 536376 358806 536380 358862
rect 536316 358802 536380 358806
rect 536316 358782 536380 358786
rect 536316 358726 536320 358782
rect 536320 358726 536376 358782
rect 536376 358726 536380 358782
rect 536316 358722 536380 358726
rect 536316 358702 536380 358706
rect 536316 358646 536320 358702
rect 536320 358646 536376 358702
rect 536376 358646 536380 358702
rect 536316 358642 536380 358646
rect 536316 358622 536380 358626
rect 536316 358566 536320 358622
rect 536320 358566 536376 358622
rect 536376 358566 536380 358622
rect 536316 358562 536380 358566
rect 536316 358542 536380 358546
rect 536316 358486 536320 358542
rect 536320 358486 536376 358542
rect 536376 358486 536380 358542
rect 536316 358482 536380 358486
rect 536316 358462 536380 358466
rect 536316 358406 536320 358462
rect 536320 358406 536376 358462
rect 536376 358406 536380 358462
rect 536316 358402 536380 358406
rect 536316 358382 536380 358386
rect 536316 358326 536320 358382
rect 536320 358326 536376 358382
rect 536376 358326 536380 358382
rect 536316 358322 536380 358326
rect 536316 358302 536380 358306
rect 536316 358246 536320 358302
rect 536320 358246 536376 358302
rect 536376 358246 536380 358302
rect 536316 358242 536380 358246
rect 536316 358222 536380 358226
rect 536316 358166 536320 358222
rect 536320 358166 536376 358222
rect 536376 358166 536380 358222
rect 536316 358162 536380 358166
rect 536316 358142 536380 358146
rect 536316 358086 536320 358142
rect 536320 358086 536376 358142
rect 536376 358086 536380 358142
rect 536316 358082 536380 358086
rect 536316 358062 536380 358066
rect 536316 358006 536320 358062
rect 536320 358006 536376 358062
rect 536376 358006 536380 358062
rect 536316 358002 536380 358006
rect 536316 357982 536380 357986
rect 536316 357926 536320 357982
rect 536320 357926 536376 357982
rect 536376 357926 536380 357982
rect 536316 357922 536380 357926
rect 536316 357902 536380 357906
rect 536316 357846 536320 357902
rect 536320 357846 536376 357902
rect 536376 357846 536380 357902
rect 536316 357842 536380 357846
rect 559712 357844 559920 358052
rect 536316 357822 536380 357826
rect 536316 357766 536320 357822
rect 536320 357766 536376 357822
rect 536376 357766 536380 357822
rect 536316 357762 536380 357766
rect 536316 357742 536380 357746
rect 536316 357686 536320 357742
rect 536320 357686 536376 357742
rect 536376 357686 536380 357742
rect 536316 357682 536380 357686
rect 536316 357662 536380 357666
rect 536316 357606 536320 357662
rect 536320 357606 536376 357662
rect 536376 357606 536380 357662
rect 536316 357602 536380 357606
rect 573540 357594 573878 357920
rect 536316 357582 536380 357586
rect 536316 357526 536320 357582
rect 536320 357526 536376 357582
rect 536376 357526 536380 357582
rect 536316 357522 536380 357526
rect 536316 357502 536380 357506
rect 536316 357446 536320 357502
rect 536320 357446 536376 357502
rect 536376 357446 536380 357502
rect 536316 357442 536380 357446
rect 559652 311536 559860 311744
rect 573492 311420 573834 311700
<< mimcap >>
rect 493438 408889 493838 408937
rect 493438 408585 493486 408889
rect 493790 408585 493838 408889
rect 493438 408537 493838 408585
rect 494138 408889 494538 408937
rect 494138 408585 494186 408889
rect 494490 408585 494538 408889
rect 494138 408537 494538 408585
rect 497198 408889 497598 408937
rect 497198 408585 497246 408889
rect 497550 408585 497598 408889
rect 497198 408537 497598 408585
rect 497898 408889 498298 408937
rect 497898 408585 497946 408889
rect 498250 408585 498298 408889
rect 497898 408537 498298 408585
rect 500958 408497 501358 408545
rect 493438 408170 493838 408218
rect 493438 407866 493486 408170
rect 493790 407866 493838 408170
rect 493438 407818 493838 407866
rect 494138 408170 494538 408218
rect 494138 407866 494186 408170
rect 494490 407866 494538 408170
rect 494138 407818 494538 407866
rect 497198 408170 497598 408218
rect 497198 407866 497246 408170
rect 497550 407866 497598 408170
rect 497198 407818 497598 407866
rect 497898 408170 498298 408218
rect 497898 407866 497946 408170
rect 498250 407866 498298 408170
rect 500958 408193 501006 408497
rect 501310 408193 501358 408497
rect 500958 408145 501358 408193
rect 501658 408497 502058 408545
rect 501658 408193 501706 408497
rect 502010 408193 502058 408497
rect 501658 408145 502058 408193
rect 497898 407818 498298 407866
rect 500958 407778 501358 407826
rect 493438 407451 493838 407499
rect 493438 407147 493486 407451
rect 493790 407147 493838 407451
rect 493438 407099 493838 407147
rect 494138 407451 494538 407499
rect 494138 407147 494186 407451
rect 494490 407147 494538 407451
rect 494138 407099 494538 407147
rect 497198 407451 497598 407499
rect 497198 407147 497246 407451
rect 497550 407147 497598 407451
rect 497198 407099 497598 407147
rect 497898 407451 498298 407499
rect 497898 407147 497946 407451
rect 498250 407147 498298 407451
rect 500958 407474 501006 407778
rect 501310 407474 501358 407778
rect 500958 407426 501358 407474
rect 501658 407778 502058 407826
rect 501658 407474 501706 407778
rect 502010 407474 502058 407778
rect 501658 407426 502058 407474
rect 497898 407099 498298 407147
rect 500958 407059 501358 407107
rect 493438 406732 493838 406780
rect 493438 406428 493486 406732
rect 493790 406428 493838 406732
rect 493438 406380 493838 406428
rect 494138 406732 494538 406780
rect 494138 406428 494186 406732
rect 494490 406428 494538 406732
rect 494138 406380 494538 406428
rect 497198 406732 497598 406780
rect 497198 406428 497246 406732
rect 497550 406428 497598 406732
rect 497198 406380 497598 406428
rect 497898 406732 498298 406780
rect 497898 406428 497946 406732
rect 498250 406428 498298 406732
rect 500958 406755 501006 407059
rect 501310 406755 501358 407059
rect 500958 406707 501358 406755
rect 501658 407059 502058 407107
rect 501658 406755 501706 407059
rect 502010 406755 502058 407059
rect 501658 406707 502058 406755
rect 497898 406380 498298 406428
rect 500958 406340 501358 406388
rect 493438 406013 493838 406061
rect 493438 405709 493486 406013
rect 493790 405709 493838 406013
rect 493438 405661 493838 405709
rect 494138 406013 494538 406061
rect 494138 405709 494186 406013
rect 494490 405709 494538 406013
rect 494138 405661 494538 405709
rect 497198 406013 497598 406061
rect 497198 405709 497246 406013
rect 497550 405709 497598 406013
rect 497198 405661 497598 405709
rect 497898 406013 498298 406061
rect 497898 405709 497946 406013
rect 498250 405709 498298 406013
rect 500958 406036 501006 406340
rect 501310 406036 501358 406340
rect 500958 405988 501358 406036
rect 501658 406340 502058 406388
rect 501658 406036 501706 406340
rect 502010 406036 502058 406340
rect 501658 405988 502058 406036
rect 497898 405661 498298 405709
rect 500958 405621 501358 405669
rect 493438 405294 493838 405342
rect 493438 404990 493486 405294
rect 493790 404990 493838 405294
rect 493438 404942 493838 404990
rect 494138 405294 494538 405342
rect 494138 404990 494186 405294
rect 494490 404990 494538 405294
rect 494138 404942 494538 404990
rect 497198 405294 497598 405342
rect 497198 404990 497246 405294
rect 497550 404990 497598 405294
rect 497198 404942 497598 404990
rect 497898 405294 498298 405342
rect 497898 404990 497946 405294
rect 498250 404990 498298 405294
rect 500958 405317 501006 405621
rect 501310 405317 501358 405621
rect 500958 405269 501358 405317
rect 501658 405621 502058 405669
rect 501658 405317 501706 405621
rect 502010 405317 502058 405621
rect 501658 405269 502058 405317
rect 497898 404942 498298 404990
rect 500958 404902 501358 404950
rect 493438 404575 493838 404623
rect 493438 404271 493486 404575
rect 493790 404271 493838 404575
rect 493438 404223 493838 404271
rect 494138 404575 494538 404623
rect 494138 404271 494186 404575
rect 494490 404271 494538 404575
rect 494138 404223 494538 404271
rect 497198 404575 497598 404623
rect 497198 404271 497246 404575
rect 497550 404271 497598 404575
rect 497198 404223 497598 404271
rect 497898 404575 498298 404623
rect 497898 404271 497946 404575
rect 498250 404271 498298 404575
rect 500958 404598 501006 404902
rect 501310 404598 501358 404902
rect 500958 404550 501358 404598
rect 501658 404902 502058 404950
rect 501658 404598 501706 404902
rect 502010 404598 502058 404902
rect 501658 404550 502058 404598
rect 497898 404223 498298 404271
rect 500958 404183 501358 404231
rect 493438 403856 493838 403904
rect 493438 403552 493486 403856
rect 493790 403552 493838 403856
rect 493438 403504 493838 403552
rect 494138 403856 494538 403904
rect 494138 403552 494186 403856
rect 494490 403552 494538 403856
rect 494138 403504 494538 403552
rect 497198 403856 497598 403904
rect 497198 403552 497246 403856
rect 497550 403552 497598 403856
rect 497198 403504 497598 403552
rect 497898 403856 498298 403904
rect 497898 403552 497946 403856
rect 498250 403552 498298 403856
rect 500958 403879 501006 404183
rect 501310 403879 501358 404183
rect 500958 403831 501358 403879
rect 501658 404183 502058 404231
rect 501658 403879 501706 404183
rect 502010 403879 502058 404183
rect 501658 403831 502058 403879
rect 497898 403504 498298 403552
rect 500958 403464 501358 403512
rect 493438 403137 493838 403185
rect 493438 402833 493486 403137
rect 493790 402833 493838 403137
rect 493438 402785 493838 402833
rect 494138 403137 494538 403185
rect 494138 402833 494186 403137
rect 494490 402833 494538 403137
rect 494138 402785 494538 402833
rect 497198 403137 497598 403185
rect 497198 402833 497246 403137
rect 497550 402833 497598 403137
rect 497198 402785 497598 402833
rect 497898 403137 498298 403185
rect 497898 402833 497946 403137
rect 498250 402833 498298 403137
rect 500958 403160 501006 403464
rect 501310 403160 501358 403464
rect 500958 403112 501358 403160
rect 501658 403464 502058 403512
rect 501658 403160 501706 403464
rect 502010 403160 502058 403464
rect 501658 403112 502058 403160
rect 497898 402785 498298 402833
rect 500958 402745 501358 402793
rect 493438 402418 493838 402466
rect 493438 402114 493486 402418
rect 493790 402114 493838 402418
rect 493438 402066 493838 402114
rect 494138 402418 494538 402466
rect 494138 402114 494186 402418
rect 494490 402114 494538 402418
rect 494138 402066 494538 402114
rect 497198 402418 497598 402466
rect 497198 402114 497246 402418
rect 497550 402114 497598 402418
rect 497198 402066 497598 402114
rect 497898 402418 498298 402466
rect 497898 402114 497946 402418
rect 498250 402114 498298 402418
rect 500958 402441 501006 402745
rect 501310 402441 501358 402745
rect 500958 402393 501358 402441
rect 501658 402745 502058 402793
rect 501658 402441 501706 402745
rect 502010 402441 502058 402745
rect 501658 402393 502058 402441
rect 497898 402066 498298 402114
rect 500958 402026 501358 402074
rect 500958 401722 501006 402026
rect 501310 401722 501358 402026
rect 500958 401674 501358 401722
rect 501658 402026 502058 402074
rect 501658 401722 501706 402026
rect 502010 401722 502058 402026
rect 501658 401674 502058 401722
rect 493438 401441 493838 401489
rect 493438 401137 493486 401441
rect 493790 401137 493838 401441
rect 493438 401089 493838 401137
rect 494138 401441 494538 401489
rect 494138 401137 494186 401441
rect 494490 401137 494538 401441
rect 494138 401089 494538 401137
rect 493438 400722 493838 400770
rect 493438 400418 493486 400722
rect 493790 400418 493838 400722
rect 493438 400370 493838 400418
rect 494138 400722 494538 400770
rect 494138 400418 494186 400722
rect 494490 400418 494538 400722
rect 494138 400370 494538 400418
rect 493438 400003 493838 400051
rect 493438 399699 493486 400003
rect 493790 399699 493838 400003
rect 493438 399651 493838 399699
rect 494138 400003 494538 400051
rect 494138 399699 494186 400003
rect 494490 399699 494538 400003
rect 494138 399651 494538 399699
rect 500958 399677 501358 399725
rect 500958 399373 501006 399677
rect 501310 399373 501358 399677
rect 493438 399284 493838 399332
rect 493438 398980 493486 399284
rect 493790 398980 493838 399284
rect 493438 398932 493838 398980
rect 494138 399284 494538 399332
rect 500958 399325 501358 399373
rect 501658 399677 502058 399725
rect 501658 399373 501706 399677
rect 502010 399373 502058 399677
rect 501658 399325 502058 399373
rect 494138 398980 494186 399284
rect 494490 398980 494538 399284
rect 494138 398932 494538 398980
rect 500958 398958 501358 399006
rect 500958 398654 501006 398958
rect 501310 398654 501358 398958
rect 493438 398565 493838 398613
rect 493438 398261 493486 398565
rect 493790 398261 493838 398565
rect 493438 398213 493838 398261
rect 494138 398565 494538 398613
rect 500958 398606 501358 398654
rect 501658 398958 502058 399006
rect 501658 398654 501706 398958
rect 502010 398654 502058 398958
rect 501658 398606 502058 398654
rect 494138 398261 494186 398565
rect 494490 398261 494538 398565
rect 494138 398213 494538 398261
rect 500958 398239 501358 398287
rect 500958 397935 501006 398239
rect 501310 397935 501358 398239
rect 493438 397846 493838 397894
rect 493438 397542 493486 397846
rect 493790 397542 493838 397846
rect 493438 397494 493838 397542
rect 494138 397846 494538 397894
rect 500958 397887 501358 397935
rect 501658 398239 502058 398287
rect 501658 397935 501706 398239
rect 502010 397935 502058 398239
rect 501658 397887 502058 397935
rect 494138 397542 494186 397846
rect 494490 397542 494538 397846
rect 494138 397494 494538 397542
rect 500958 397520 501358 397568
rect 500958 397216 501006 397520
rect 501310 397216 501358 397520
rect 493438 397127 493838 397175
rect 493438 396823 493486 397127
rect 493790 396823 493838 397127
rect 493438 396775 493838 396823
rect 494138 397127 494538 397175
rect 500958 397168 501358 397216
rect 501658 397520 502058 397568
rect 501658 397216 501706 397520
rect 502010 397216 502058 397520
rect 501658 397168 502058 397216
rect 494138 396823 494186 397127
rect 494490 396823 494538 397127
rect 494138 396775 494538 396823
rect 500958 396801 501358 396849
rect 500958 396497 501006 396801
rect 501310 396497 501358 396801
rect 493438 396408 493838 396456
rect 493438 396104 493486 396408
rect 493790 396104 493838 396408
rect 493438 396056 493838 396104
rect 494138 396408 494538 396456
rect 500958 396449 501358 396497
rect 501658 396801 502058 396849
rect 501658 396497 501706 396801
rect 502010 396497 502058 396801
rect 501658 396449 502058 396497
rect 494138 396104 494186 396408
rect 494490 396104 494538 396408
rect 494138 396056 494538 396104
rect 500958 396082 501358 396130
rect 500958 395778 501006 396082
rect 501310 395778 501358 396082
rect 493438 395689 493838 395737
rect 493438 395385 493486 395689
rect 493790 395385 493838 395689
rect 493438 395337 493838 395385
rect 494138 395689 494538 395737
rect 500958 395730 501358 395778
rect 501658 396082 502058 396130
rect 501658 395778 501706 396082
rect 502010 395778 502058 396082
rect 501658 395730 502058 395778
rect 494138 395385 494186 395689
rect 494490 395385 494538 395689
rect 494138 395337 494538 395385
rect 500958 395363 501358 395411
rect 500958 395059 501006 395363
rect 501310 395059 501358 395363
rect 493438 394970 493838 395018
rect 493438 394666 493486 394970
rect 493790 394666 493838 394970
rect 493438 394618 493838 394666
rect 494138 394970 494538 395018
rect 500958 395011 501358 395059
rect 501658 395363 502058 395411
rect 501658 395059 501706 395363
rect 502010 395059 502058 395363
rect 501658 395011 502058 395059
rect 494138 394666 494186 394970
rect 494490 394666 494538 394970
rect 494138 394618 494538 394666
rect 500958 394644 501358 394692
rect 500958 394340 501006 394644
rect 501310 394340 501358 394644
rect 500958 394292 501358 394340
rect 501658 394644 502058 394692
rect 501658 394340 501706 394644
rect 502010 394340 502058 394644
rect 501658 394292 502058 394340
rect 500958 393925 501358 393973
rect 500958 393621 501006 393925
rect 501310 393621 501358 393925
rect 500958 393573 501358 393621
rect 501658 393925 502058 393973
rect 501658 393621 501706 393925
rect 502010 393621 502058 393925
rect 501658 393573 502058 393621
rect 500958 393206 501358 393254
rect 500958 392902 501006 393206
rect 501310 392902 501358 393206
rect 500958 392854 501358 392902
rect 501658 393206 502058 393254
rect 501658 392902 501706 393206
rect 502010 392902 502058 393206
rect 501658 392854 502058 392902
rect 508478 388603 508878 388651
rect 508478 388299 508526 388603
rect 508830 388299 508878 388603
rect 508478 388251 508878 388299
rect 509178 388603 509578 388651
rect 509178 388299 509226 388603
rect 509530 388299 509578 388603
rect 509178 388251 509578 388299
rect 508478 387884 508878 387932
rect 508478 387580 508526 387884
rect 508830 387580 508878 387884
rect 508478 387532 508878 387580
rect 509178 387884 509578 387932
rect 509178 387580 509226 387884
rect 509530 387580 509578 387884
rect 509178 387532 509578 387580
rect 508478 387165 508878 387213
rect 508478 386861 508526 387165
rect 508830 386861 508878 387165
rect 508478 386813 508878 386861
rect 509178 387165 509578 387213
rect 509178 386861 509226 387165
rect 509530 386861 509578 387165
rect 509178 386813 509578 386861
rect 508478 386446 508878 386494
rect 508478 386142 508526 386446
rect 508830 386142 508878 386446
rect 508478 386094 508878 386142
rect 509178 386446 509578 386494
rect 509178 386142 509226 386446
rect 509530 386142 509578 386446
rect 509178 386094 509578 386142
rect 508478 385727 508878 385775
rect 508478 385423 508526 385727
rect 508830 385423 508878 385727
rect 508478 385375 508878 385423
rect 509178 385727 509578 385775
rect 509178 385423 509226 385727
rect 509530 385423 509578 385727
rect 509178 385375 509578 385423
rect 508478 385008 508878 385056
rect 504718 384879 505118 384927
rect 504718 384575 504766 384879
rect 505070 384575 505118 384879
rect 504718 384527 505118 384575
rect 505418 384879 505818 384927
rect 505418 384575 505466 384879
rect 505770 384575 505818 384879
rect 508478 384704 508526 385008
rect 508830 384704 508878 385008
rect 508478 384656 508878 384704
rect 509178 385008 509578 385056
rect 509178 384704 509226 385008
rect 509530 384704 509578 385008
rect 509178 384656 509578 384704
rect 512238 384879 512638 384927
rect 505418 384527 505818 384575
rect 512238 384575 512286 384879
rect 512590 384575 512638 384879
rect 512238 384527 512638 384575
rect 512938 384879 513338 384927
rect 512938 384575 512986 384879
rect 513290 384575 513338 384879
rect 512938 384527 513338 384575
rect 515998 384879 516398 384927
rect 515998 384575 516046 384879
rect 516350 384575 516398 384879
rect 515998 384527 516398 384575
rect 516698 384879 517098 384927
rect 516698 384575 516746 384879
rect 517050 384575 517098 384879
rect 516698 384527 517098 384575
rect 508478 384289 508878 384337
rect 504718 384160 505118 384208
rect 504718 383856 504766 384160
rect 505070 383856 505118 384160
rect 504718 383808 505118 383856
rect 505418 384160 505818 384208
rect 505418 383856 505466 384160
rect 505770 383856 505818 384160
rect 508478 383985 508526 384289
rect 508830 383985 508878 384289
rect 508478 383937 508878 383985
rect 509178 384289 509578 384337
rect 509178 383985 509226 384289
rect 509530 383985 509578 384289
rect 509178 383937 509578 383985
rect 512238 384160 512638 384208
rect 505418 383808 505818 383856
rect 512238 383856 512286 384160
rect 512590 383856 512638 384160
rect 512238 383808 512638 383856
rect 512938 384160 513338 384208
rect 512938 383856 512986 384160
rect 513290 383856 513338 384160
rect 512938 383808 513338 383856
rect 515998 384160 516398 384208
rect 515998 383856 516046 384160
rect 516350 383856 516398 384160
rect 515998 383808 516398 383856
rect 516698 384160 517098 384208
rect 516698 383856 516746 384160
rect 517050 383856 517098 384160
rect 516698 383808 517098 383856
rect 508478 383570 508878 383618
rect 504718 383441 505118 383489
rect 504718 383137 504766 383441
rect 505070 383137 505118 383441
rect 504718 383089 505118 383137
rect 505418 383441 505818 383489
rect 505418 383137 505466 383441
rect 505770 383137 505818 383441
rect 508478 383266 508526 383570
rect 508830 383266 508878 383570
rect 508478 383218 508878 383266
rect 509178 383570 509578 383618
rect 509178 383266 509226 383570
rect 509530 383266 509578 383570
rect 509178 383218 509578 383266
rect 512238 383441 512638 383489
rect 505418 383089 505818 383137
rect 512238 383137 512286 383441
rect 512590 383137 512638 383441
rect 512238 383089 512638 383137
rect 512938 383441 513338 383489
rect 512938 383137 512986 383441
rect 513290 383137 513338 383441
rect 512938 383089 513338 383137
rect 515998 383441 516398 383489
rect 515998 383137 516046 383441
rect 516350 383137 516398 383441
rect 515998 383089 516398 383137
rect 516698 383441 517098 383489
rect 516698 383137 516746 383441
rect 517050 383137 517098 383441
rect 516698 383089 517098 383137
rect 508478 382851 508878 382899
rect 504718 382722 505118 382770
rect 504718 382418 504766 382722
rect 505070 382418 505118 382722
rect 504718 382370 505118 382418
rect 505418 382722 505818 382770
rect 505418 382418 505466 382722
rect 505770 382418 505818 382722
rect 508478 382547 508526 382851
rect 508830 382547 508878 382851
rect 508478 382499 508878 382547
rect 509178 382851 509578 382899
rect 509178 382547 509226 382851
rect 509530 382547 509578 382851
rect 509178 382499 509578 382547
rect 512238 382722 512638 382770
rect 505418 382370 505818 382418
rect 512238 382418 512286 382722
rect 512590 382418 512638 382722
rect 512238 382370 512638 382418
rect 512938 382722 513338 382770
rect 512938 382418 512986 382722
rect 513290 382418 513338 382722
rect 512938 382370 513338 382418
rect 515998 382722 516398 382770
rect 515998 382418 516046 382722
rect 516350 382418 516398 382722
rect 515998 382370 516398 382418
rect 516698 382722 517098 382770
rect 516698 382418 516746 382722
rect 517050 382418 517098 382722
rect 516698 382370 517098 382418
rect 508478 382132 508878 382180
rect 504718 382003 505118 382051
rect 504718 381699 504766 382003
rect 505070 381699 505118 382003
rect 504718 381651 505118 381699
rect 505418 382003 505818 382051
rect 505418 381699 505466 382003
rect 505770 381699 505818 382003
rect 508478 381828 508526 382132
rect 508830 381828 508878 382132
rect 508478 381780 508878 381828
rect 509178 382132 509578 382180
rect 509178 381828 509226 382132
rect 509530 381828 509578 382132
rect 509178 381780 509578 381828
rect 512238 382003 512638 382051
rect 505418 381651 505818 381699
rect 512238 381699 512286 382003
rect 512590 381699 512638 382003
rect 512238 381651 512638 381699
rect 512938 382003 513338 382051
rect 512938 381699 512986 382003
rect 513290 381699 513338 382003
rect 512938 381651 513338 381699
rect 515998 382003 516398 382051
rect 515998 381699 516046 382003
rect 516350 381699 516398 382003
rect 515998 381651 516398 381699
rect 516698 382003 517098 382051
rect 516698 381699 516746 382003
rect 517050 381699 517098 382003
rect 516698 381651 517098 381699
rect 504718 381284 505118 381332
rect 504718 380980 504766 381284
rect 505070 380980 505118 381284
rect 504718 380932 505118 380980
rect 505418 381284 505818 381332
rect 505418 380980 505466 381284
rect 505770 380980 505818 381284
rect 512238 381284 512638 381332
rect 505418 380932 505818 380980
rect 508478 381155 508878 381203
rect 508478 380851 508526 381155
rect 508830 380851 508878 381155
rect 508478 380803 508878 380851
rect 509178 381155 509578 381203
rect 509178 380851 509226 381155
rect 509530 380851 509578 381155
rect 512238 380980 512286 381284
rect 512590 380980 512638 381284
rect 512238 380932 512638 380980
rect 512938 381284 513338 381332
rect 512938 380980 512986 381284
rect 513290 380980 513338 381284
rect 512938 380932 513338 380980
rect 515998 381284 516398 381332
rect 515998 380980 516046 381284
rect 516350 380980 516398 381284
rect 515998 380932 516398 380980
rect 516698 381284 517098 381332
rect 516698 380980 516746 381284
rect 517050 380980 517098 381284
rect 516698 380932 517098 380980
rect 509178 380803 509578 380851
rect 504718 380565 505118 380613
rect 504718 380261 504766 380565
rect 505070 380261 505118 380565
rect 504718 380213 505118 380261
rect 505418 380565 505818 380613
rect 505418 380261 505466 380565
rect 505770 380261 505818 380565
rect 512238 380565 512638 380613
rect 505418 380213 505818 380261
rect 508478 380436 508878 380484
rect 508478 380132 508526 380436
rect 508830 380132 508878 380436
rect 508478 380084 508878 380132
rect 509178 380436 509578 380484
rect 509178 380132 509226 380436
rect 509530 380132 509578 380436
rect 512238 380261 512286 380565
rect 512590 380261 512638 380565
rect 512238 380213 512638 380261
rect 512938 380565 513338 380613
rect 512938 380261 512986 380565
rect 513290 380261 513338 380565
rect 512938 380213 513338 380261
rect 515998 380565 516398 380613
rect 515998 380261 516046 380565
rect 516350 380261 516398 380565
rect 515998 380213 516398 380261
rect 516698 380565 517098 380613
rect 516698 380261 516746 380565
rect 517050 380261 517098 380565
rect 516698 380213 517098 380261
rect 509178 380084 509578 380132
rect 504718 379846 505118 379894
rect 504718 379542 504766 379846
rect 505070 379542 505118 379846
rect 504718 379494 505118 379542
rect 505418 379846 505818 379894
rect 505418 379542 505466 379846
rect 505770 379542 505818 379846
rect 512238 379846 512638 379894
rect 505418 379494 505818 379542
rect 508478 379717 508878 379765
rect 508478 379413 508526 379717
rect 508830 379413 508878 379717
rect 508478 379365 508878 379413
rect 509178 379717 509578 379765
rect 509178 379413 509226 379717
rect 509530 379413 509578 379717
rect 512238 379542 512286 379846
rect 512590 379542 512638 379846
rect 512238 379494 512638 379542
rect 512938 379846 513338 379894
rect 512938 379542 512986 379846
rect 513290 379542 513338 379846
rect 512938 379494 513338 379542
rect 515998 379846 516398 379894
rect 515998 379542 516046 379846
rect 516350 379542 516398 379846
rect 515998 379494 516398 379542
rect 516698 379846 517098 379894
rect 516698 379542 516746 379846
rect 517050 379542 517098 379846
rect 516698 379494 517098 379542
rect 509178 379365 509578 379413
rect 504718 379127 505118 379175
rect 504718 378823 504766 379127
rect 505070 378823 505118 379127
rect 504718 378775 505118 378823
rect 505418 379127 505818 379175
rect 505418 378823 505466 379127
rect 505770 378823 505818 379127
rect 512238 379127 512638 379175
rect 505418 378775 505818 378823
rect 508478 378998 508878 379046
rect 508478 378694 508526 378998
rect 508830 378694 508878 378998
rect 508478 378646 508878 378694
rect 509178 378998 509578 379046
rect 509178 378694 509226 378998
rect 509530 378694 509578 378998
rect 512238 378823 512286 379127
rect 512590 378823 512638 379127
rect 512238 378775 512638 378823
rect 512938 379127 513338 379175
rect 512938 378823 512986 379127
rect 513290 378823 513338 379127
rect 512938 378775 513338 378823
rect 515998 379127 516398 379175
rect 515998 378823 516046 379127
rect 516350 378823 516398 379127
rect 515998 378775 516398 378823
rect 516698 379127 517098 379175
rect 516698 378823 516746 379127
rect 517050 378823 517098 379127
rect 516698 378775 517098 378823
rect 509178 378646 509578 378694
rect 504718 378408 505118 378456
rect 504718 378104 504766 378408
rect 505070 378104 505118 378408
rect 504718 378056 505118 378104
rect 505418 378408 505818 378456
rect 505418 378104 505466 378408
rect 505770 378104 505818 378408
rect 512238 378408 512638 378456
rect 505418 378056 505818 378104
rect 508478 378279 508878 378327
rect 508478 377975 508526 378279
rect 508830 377975 508878 378279
rect 508478 377927 508878 377975
rect 509178 378279 509578 378327
rect 509178 377975 509226 378279
rect 509530 377975 509578 378279
rect 512238 378104 512286 378408
rect 512590 378104 512638 378408
rect 512238 378056 512638 378104
rect 512938 378408 513338 378456
rect 512938 378104 512986 378408
rect 513290 378104 513338 378408
rect 512938 378056 513338 378104
rect 515998 378408 516398 378456
rect 515998 378104 516046 378408
rect 516350 378104 516398 378408
rect 515998 378056 516398 378104
rect 516698 378408 517098 378456
rect 516698 378104 516746 378408
rect 517050 378104 517098 378408
rect 516698 378056 517098 378104
rect 509178 377927 509578 377975
rect 508478 377560 508878 377608
rect 508478 377256 508526 377560
rect 508830 377256 508878 377560
rect 508478 377208 508878 377256
rect 509178 377560 509578 377608
rect 509178 377256 509226 377560
rect 509530 377256 509578 377560
rect 509178 377208 509578 377256
rect 508478 376841 508878 376889
rect 508478 376537 508526 376841
rect 508830 376537 508878 376841
rect 508478 376489 508878 376537
rect 509178 376841 509578 376889
rect 509178 376537 509226 376841
rect 509530 376537 509578 376841
rect 509178 376489 509578 376537
rect 508478 376122 508878 376170
rect 508478 375818 508526 376122
rect 508830 375818 508878 376122
rect 508478 375770 508878 375818
rect 509178 376122 509578 376170
rect 509178 375818 509226 376122
rect 509530 375818 509578 376122
rect 509178 375770 509578 375818
rect 508478 375403 508878 375451
rect 508478 375099 508526 375403
rect 508830 375099 508878 375403
rect 508478 375051 508878 375099
rect 509178 375403 509578 375451
rect 509178 375099 509226 375403
rect 509530 375099 509578 375403
rect 509178 375051 509578 375099
rect 508478 374684 508878 374732
rect 508478 374380 508526 374684
rect 508830 374380 508878 374684
rect 508478 374332 508878 374380
rect 509178 374684 509578 374732
rect 509178 374380 509226 374684
rect 509530 374380 509578 374684
rect 509178 374332 509578 374380
<< mimcapcontact >>
rect 493486 408585 493790 408889
rect 494186 408585 494490 408889
rect 497246 408585 497550 408889
rect 497946 408585 498250 408889
rect 493486 407866 493790 408170
rect 494186 407866 494490 408170
rect 497246 407866 497550 408170
rect 497946 407866 498250 408170
rect 501006 408193 501310 408497
rect 501706 408193 502010 408497
rect 493486 407147 493790 407451
rect 494186 407147 494490 407451
rect 497246 407147 497550 407451
rect 497946 407147 498250 407451
rect 501006 407474 501310 407778
rect 501706 407474 502010 407778
rect 493486 406428 493790 406732
rect 494186 406428 494490 406732
rect 497246 406428 497550 406732
rect 497946 406428 498250 406732
rect 501006 406755 501310 407059
rect 501706 406755 502010 407059
rect 493486 405709 493790 406013
rect 494186 405709 494490 406013
rect 497246 405709 497550 406013
rect 497946 405709 498250 406013
rect 501006 406036 501310 406340
rect 501706 406036 502010 406340
rect 493486 404990 493790 405294
rect 494186 404990 494490 405294
rect 497246 404990 497550 405294
rect 497946 404990 498250 405294
rect 501006 405317 501310 405621
rect 501706 405317 502010 405621
rect 493486 404271 493790 404575
rect 494186 404271 494490 404575
rect 497246 404271 497550 404575
rect 497946 404271 498250 404575
rect 501006 404598 501310 404902
rect 501706 404598 502010 404902
rect 493486 403552 493790 403856
rect 494186 403552 494490 403856
rect 497246 403552 497550 403856
rect 497946 403552 498250 403856
rect 501006 403879 501310 404183
rect 501706 403879 502010 404183
rect 493486 402833 493790 403137
rect 494186 402833 494490 403137
rect 497246 402833 497550 403137
rect 497946 402833 498250 403137
rect 501006 403160 501310 403464
rect 501706 403160 502010 403464
rect 493486 402114 493790 402418
rect 494186 402114 494490 402418
rect 497246 402114 497550 402418
rect 497946 402114 498250 402418
rect 501006 402441 501310 402745
rect 501706 402441 502010 402745
rect 501006 401722 501310 402026
rect 501706 401722 502010 402026
rect 493486 401137 493790 401441
rect 494186 401137 494490 401441
rect 493486 400418 493790 400722
rect 494186 400418 494490 400722
rect 493486 399699 493790 400003
rect 494186 399699 494490 400003
rect 501006 399373 501310 399677
rect 493486 398980 493790 399284
rect 501706 399373 502010 399677
rect 494186 398980 494490 399284
rect 501006 398654 501310 398958
rect 493486 398261 493790 398565
rect 501706 398654 502010 398958
rect 494186 398261 494490 398565
rect 501006 397935 501310 398239
rect 493486 397542 493790 397846
rect 501706 397935 502010 398239
rect 494186 397542 494490 397846
rect 501006 397216 501310 397520
rect 493486 396823 493790 397127
rect 501706 397216 502010 397520
rect 494186 396823 494490 397127
rect 501006 396497 501310 396801
rect 493486 396104 493790 396408
rect 501706 396497 502010 396801
rect 494186 396104 494490 396408
rect 501006 395778 501310 396082
rect 493486 395385 493790 395689
rect 501706 395778 502010 396082
rect 494186 395385 494490 395689
rect 501006 395059 501310 395363
rect 493486 394666 493790 394970
rect 501706 395059 502010 395363
rect 494186 394666 494490 394970
rect 501006 394340 501310 394644
rect 501706 394340 502010 394644
rect 501006 393621 501310 393925
rect 501706 393621 502010 393925
rect 501006 392902 501310 393206
rect 501706 392902 502010 393206
rect 508526 388299 508830 388603
rect 509226 388299 509530 388603
rect 508526 387580 508830 387884
rect 509226 387580 509530 387884
rect 508526 386861 508830 387165
rect 509226 386861 509530 387165
rect 508526 386142 508830 386446
rect 509226 386142 509530 386446
rect 508526 385423 508830 385727
rect 509226 385423 509530 385727
rect 504766 384575 505070 384879
rect 505466 384575 505770 384879
rect 508526 384704 508830 385008
rect 509226 384704 509530 385008
rect 512286 384575 512590 384879
rect 512986 384575 513290 384879
rect 516046 384575 516350 384879
rect 516746 384575 517050 384879
rect 504766 383856 505070 384160
rect 505466 383856 505770 384160
rect 508526 383985 508830 384289
rect 509226 383985 509530 384289
rect 512286 383856 512590 384160
rect 512986 383856 513290 384160
rect 516046 383856 516350 384160
rect 516746 383856 517050 384160
rect 504766 383137 505070 383441
rect 505466 383137 505770 383441
rect 508526 383266 508830 383570
rect 509226 383266 509530 383570
rect 512286 383137 512590 383441
rect 512986 383137 513290 383441
rect 516046 383137 516350 383441
rect 516746 383137 517050 383441
rect 504766 382418 505070 382722
rect 505466 382418 505770 382722
rect 508526 382547 508830 382851
rect 509226 382547 509530 382851
rect 512286 382418 512590 382722
rect 512986 382418 513290 382722
rect 516046 382418 516350 382722
rect 516746 382418 517050 382722
rect 504766 381699 505070 382003
rect 505466 381699 505770 382003
rect 508526 381828 508830 382132
rect 509226 381828 509530 382132
rect 512286 381699 512590 382003
rect 512986 381699 513290 382003
rect 516046 381699 516350 382003
rect 516746 381699 517050 382003
rect 504766 380980 505070 381284
rect 505466 380980 505770 381284
rect 508526 380851 508830 381155
rect 509226 380851 509530 381155
rect 512286 380980 512590 381284
rect 512986 380980 513290 381284
rect 516046 380980 516350 381284
rect 516746 380980 517050 381284
rect 504766 380261 505070 380565
rect 505466 380261 505770 380565
rect 508526 380132 508830 380436
rect 509226 380132 509530 380436
rect 512286 380261 512590 380565
rect 512986 380261 513290 380565
rect 516046 380261 516350 380565
rect 516746 380261 517050 380565
rect 504766 379542 505070 379846
rect 505466 379542 505770 379846
rect 508526 379413 508830 379717
rect 509226 379413 509530 379717
rect 512286 379542 512590 379846
rect 512986 379542 513290 379846
rect 516046 379542 516350 379846
rect 516746 379542 517050 379846
rect 504766 378823 505070 379127
rect 505466 378823 505770 379127
rect 508526 378694 508830 378998
rect 509226 378694 509530 378998
rect 512286 378823 512590 379127
rect 512986 378823 513290 379127
rect 516046 378823 516350 379127
rect 516746 378823 517050 379127
rect 504766 378104 505070 378408
rect 505466 378104 505770 378408
rect 508526 377975 508830 378279
rect 509226 377975 509530 378279
rect 512286 378104 512590 378408
rect 512986 378104 513290 378408
rect 516046 378104 516350 378408
rect 516746 378104 517050 378408
rect 508526 377256 508830 377560
rect 509226 377256 509530 377560
rect 508526 376537 508830 376841
rect 509226 376537 509530 376841
rect 508526 375818 508830 376122
rect 509226 375818 509530 376122
rect 508526 375099 508830 375403
rect 509226 375099 509530 375403
rect 508526 374380 508830 374684
rect 509226 374380 509530 374684
<< metal4 >>
rect 502376 697378 560022 697790
rect 502376 689882 510704 697378
rect 515202 697354 560022 697378
rect 515202 689882 520704 697354
rect 502376 689858 520704 689882
rect 525202 689858 560022 697354
rect 502376 689742 560022 689858
rect 551974 492536 560022 689742
rect 567305 644324 573723 644325
rect 567305 640080 567306 644324
rect 573722 640080 573723 644324
rect 567305 640079 573723 640080
rect 567305 634256 573723 634257
rect 567305 630012 567306 634256
rect 573722 630012 573723 634256
rect 567305 630011 573723 630012
rect 551974 492324 559802 492536
rect 560012 492324 560022 492536
rect 551974 414054 560022 492324
rect 573563 492160 573875 492161
rect 573563 491888 573564 492160
rect 573874 491888 573875 492160
rect 573563 491887 573875 491888
rect 485484 414030 560022 414054
rect 485484 413996 491196 414030
rect 485484 412480 486390 413996
rect 487906 413966 491196 413996
rect 491260 413966 494956 414030
rect 495020 413966 498716 414030
rect 498780 413966 502476 414030
rect 502540 413966 506236 414030
rect 506300 413966 509996 414030
rect 510060 413966 513756 414030
rect 513820 413966 517516 414030
rect 517580 413966 521276 414030
rect 521340 413966 525036 414030
rect 525100 413966 528796 414030
rect 528860 413966 532556 414030
rect 532620 413966 536316 414030
rect 536380 413996 560022 414030
rect 536380 413966 539670 413996
rect 487906 413950 539670 413966
rect 487906 413886 491196 413950
rect 491260 413886 494956 413950
rect 495020 413886 498716 413950
rect 498780 413886 502476 413950
rect 502540 413886 506236 413950
rect 506300 413886 509996 413950
rect 510060 413886 513756 413950
rect 513820 413886 517516 413950
rect 517580 413886 521276 413950
rect 521340 413886 525036 413950
rect 525100 413886 528796 413950
rect 528860 413886 532556 413950
rect 532620 413886 536316 413950
rect 536380 413886 539670 413950
rect 487906 413870 539670 413886
rect 487906 413806 491196 413870
rect 491260 413806 494956 413870
rect 495020 413806 498716 413870
rect 498780 413806 502476 413870
rect 502540 413806 506236 413870
rect 506300 413806 509996 413870
rect 510060 413806 513756 413870
rect 513820 413806 517516 413870
rect 517580 413806 521276 413870
rect 521340 413806 525036 413870
rect 525100 413806 528796 413870
rect 528860 413806 532556 413870
rect 532620 413806 536316 413870
rect 536380 413806 539670 413870
rect 487906 413790 539670 413806
rect 487906 413726 491196 413790
rect 491260 413726 494956 413790
rect 495020 413726 498716 413790
rect 498780 413726 502476 413790
rect 502540 413726 506236 413790
rect 506300 413726 509996 413790
rect 510060 413726 513756 413790
rect 513820 413726 517516 413790
rect 517580 413726 521276 413790
rect 521340 413726 525036 413790
rect 525100 413726 528796 413790
rect 528860 413726 532556 413790
rect 532620 413726 536316 413790
rect 536380 413726 539670 413790
rect 487906 413710 539670 413726
rect 487906 413646 491196 413710
rect 491260 413646 494956 413710
rect 495020 413646 498716 413710
rect 498780 413646 502476 413710
rect 502540 413646 506236 413710
rect 506300 413646 509996 413710
rect 510060 413646 513756 413710
rect 513820 413646 517516 413710
rect 517580 413646 521276 413710
rect 521340 413646 525036 413710
rect 525100 413646 528796 413710
rect 528860 413646 532556 413710
rect 532620 413646 536316 413710
rect 536380 413646 539670 413710
rect 487906 413630 539670 413646
rect 487906 413566 491196 413630
rect 491260 413566 494956 413630
rect 495020 413566 498716 413630
rect 498780 413566 502476 413630
rect 502540 413566 506236 413630
rect 506300 413566 509996 413630
rect 510060 413566 513756 413630
rect 513820 413566 517516 413630
rect 517580 413566 521276 413630
rect 521340 413566 525036 413630
rect 525100 413566 528796 413630
rect 528860 413566 532556 413630
rect 532620 413566 536316 413630
rect 536380 413566 539670 413630
rect 487906 413550 539670 413566
rect 487906 413486 491196 413550
rect 491260 413486 494956 413550
rect 495020 413486 498716 413550
rect 498780 413486 502476 413550
rect 502540 413486 506236 413550
rect 506300 413486 509996 413550
rect 510060 413486 513756 413550
rect 513820 413486 517516 413550
rect 517580 413486 521276 413550
rect 521340 413486 525036 413550
rect 525100 413486 528796 413550
rect 528860 413486 532556 413550
rect 532620 413486 536316 413550
rect 536380 413486 539670 413550
rect 487906 413470 539670 413486
rect 487906 413406 491196 413470
rect 491260 413406 494956 413470
rect 495020 413406 498716 413470
rect 498780 413406 502476 413470
rect 502540 413406 506236 413470
rect 506300 413406 509996 413470
rect 510060 413406 513756 413470
rect 513820 413406 517516 413470
rect 517580 413406 521276 413470
rect 521340 413406 525036 413470
rect 525100 413406 528796 413470
rect 528860 413406 532556 413470
rect 532620 413406 536316 413470
rect 536380 413406 539670 413470
rect 487906 413390 539670 413406
rect 487906 413326 491196 413390
rect 491260 413326 494956 413390
rect 495020 413326 498716 413390
rect 498780 413326 502476 413390
rect 502540 413326 506236 413390
rect 506300 413326 509996 413390
rect 510060 413326 513756 413390
rect 513820 413326 517516 413390
rect 517580 413326 521276 413390
rect 521340 413326 525036 413390
rect 525100 413326 528796 413390
rect 528860 413326 532556 413390
rect 532620 413326 536316 413390
rect 536380 413326 539670 413390
rect 487906 413310 539670 413326
rect 487906 413246 491196 413310
rect 491260 413246 494956 413310
rect 495020 413246 498716 413310
rect 498780 413246 502476 413310
rect 502540 413246 506236 413310
rect 506300 413246 509996 413310
rect 510060 413246 513756 413310
rect 513820 413246 517516 413310
rect 517580 413246 521276 413310
rect 521340 413246 525036 413310
rect 525100 413246 528796 413310
rect 528860 413246 532556 413310
rect 532620 413246 536316 413310
rect 536380 413246 539670 413310
rect 487906 413230 539670 413246
rect 487906 413166 491196 413230
rect 491260 413166 494956 413230
rect 495020 413166 498716 413230
rect 498780 413166 502476 413230
rect 502540 413166 506236 413230
rect 506300 413166 509996 413230
rect 510060 413166 513756 413230
rect 513820 413166 517516 413230
rect 517580 413166 521276 413230
rect 521340 413166 525036 413230
rect 525100 413166 528796 413230
rect 528860 413166 532556 413230
rect 532620 413166 536316 413230
rect 536380 413166 539670 413230
rect 487906 413150 539670 413166
rect 487906 413086 491196 413150
rect 491260 413086 494956 413150
rect 495020 413086 498716 413150
rect 498780 413086 502476 413150
rect 502540 413086 506236 413150
rect 506300 413086 509996 413150
rect 510060 413086 513756 413150
rect 513820 413086 517516 413150
rect 517580 413086 521276 413150
rect 521340 413086 525036 413150
rect 525100 413086 528796 413150
rect 528860 413086 532556 413150
rect 532620 413086 536316 413150
rect 536380 413086 539670 413150
rect 487906 413070 539670 413086
rect 487906 413006 491196 413070
rect 491260 413006 494956 413070
rect 495020 413006 498716 413070
rect 498780 413006 502476 413070
rect 502540 413006 506236 413070
rect 506300 413006 509996 413070
rect 510060 413006 513756 413070
rect 513820 413006 517516 413070
rect 517580 413006 521276 413070
rect 521340 413006 525036 413070
rect 525100 413006 528796 413070
rect 528860 413006 532556 413070
rect 532620 413006 536316 413070
rect 536380 413006 539670 413070
rect 487906 412990 539670 413006
rect 487906 412926 491196 412990
rect 491260 412926 494956 412990
rect 495020 412926 498716 412990
rect 498780 412926 502476 412990
rect 502540 412926 506236 412990
rect 506300 412926 509996 412990
rect 510060 412926 513756 412990
rect 513820 412926 517516 412990
rect 517580 412926 521276 412990
rect 521340 412926 525036 412990
rect 525100 412926 528796 412990
rect 528860 412926 532556 412990
rect 532620 412926 536316 412990
rect 536380 412926 539670 412990
rect 487906 412910 539670 412926
rect 487906 412846 491196 412910
rect 491260 412846 494956 412910
rect 495020 412846 498716 412910
rect 498780 412846 502476 412910
rect 502540 412846 506236 412910
rect 506300 412846 509996 412910
rect 510060 412846 513756 412910
rect 513820 412846 517516 412910
rect 517580 412846 521276 412910
rect 521340 412846 525036 412910
rect 525100 412846 528796 412910
rect 528860 412846 532556 412910
rect 532620 412846 536316 412910
rect 536380 412846 539670 412910
rect 487906 412830 539670 412846
rect 487906 412766 491196 412830
rect 491260 412766 494956 412830
rect 495020 412766 498716 412830
rect 498780 412766 502476 412830
rect 502540 412766 506236 412830
rect 506300 412766 509996 412830
rect 510060 412766 513756 412830
rect 513820 412766 517516 412830
rect 517580 412766 521276 412830
rect 521340 412766 525036 412830
rect 525100 412766 528796 412830
rect 528860 412766 532556 412830
rect 532620 412766 536316 412830
rect 536380 412766 539670 412830
rect 487906 412750 539670 412766
rect 487906 412686 491196 412750
rect 491260 412686 494956 412750
rect 495020 412686 498716 412750
rect 498780 412686 502476 412750
rect 502540 412686 506236 412750
rect 506300 412686 509996 412750
rect 510060 412686 513756 412750
rect 513820 412686 517516 412750
rect 517580 412686 521276 412750
rect 521340 412686 525036 412750
rect 525100 412686 528796 412750
rect 528860 412686 532556 412750
rect 532620 412686 536316 412750
rect 536380 412686 539670 412750
rect 487906 412670 539670 412686
rect 487906 412606 491196 412670
rect 491260 412606 494956 412670
rect 495020 412606 498716 412670
rect 498780 412606 502476 412670
rect 502540 412606 506236 412670
rect 506300 412606 509996 412670
rect 510060 412606 513756 412670
rect 513820 412606 517516 412670
rect 517580 412606 521276 412670
rect 521340 412606 525036 412670
rect 525100 412606 528796 412670
rect 528860 412606 532556 412670
rect 532620 412606 536316 412670
rect 536380 412606 539670 412670
rect 487906 412590 539670 412606
rect 487906 412526 491196 412590
rect 491260 412526 494956 412590
rect 495020 412526 498716 412590
rect 498780 412526 502476 412590
rect 502540 412526 506236 412590
rect 506300 412526 509996 412590
rect 510060 412526 513756 412590
rect 513820 412526 517516 412590
rect 517580 412526 521276 412590
rect 521340 412526 525036 412590
rect 525100 412526 528796 412590
rect 528860 412526 532556 412590
rect 532620 412526 536316 412590
rect 536380 412526 539670 412590
rect 487906 412510 539670 412526
rect 487906 412480 491196 412510
rect 485484 412446 491196 412480
rect 491260 412446 494956 412510
rect 495020 412446 498716 412510
rect 498780 412446 502476 412510
rect 502540 412446 506236 412510
rect 506300 412446 509996 412510
rect 510060 412446 513756 412510
rect 513820 412446 517516 412510
rect 517580 412446 521276 412510
rect 521340 412446 525036 412510
rect 525100 412446 528796 412510
rect 528860 412446 532556 412510
rect 532620 412446 536316 412510
rect 536380 412480 539670 412510
rect 541186 412480 560022 413996
rect 536380 412446 560022 412480
rect 485484 412422 560022 412446
rect 485484 411582 542060 411606
rect 485484 411548 493076 411582
rect 485484 410032 488838 411548
rect 490354 411518 493076 411548
rect 493140 411518 496836 411582
rect 496900 411518 500596 411582
rect 500660 411518 504356 411582
rect 504420 411518 508116 411582
rect 508180 411518 511876 411582
rect 511940 411518 515636 411582
rect 515700 411518 519396 411582
rect 519460 411518 523156 411582
rect 523220 411518 526916 411582
rect 526980 411518 530676 411582
rect 530740 411518 534436 411582
rect 534500 411548 542060 411582
rect 534500 411518 537222 411548
rect 490354 411502 537222 411518
rect 490354 411438 493076 411502
rect 493140 411438 496836 411502
rect 496900 411438 500596 411502
rect 500660 411438 504356 411502
rect 504420 411438 508116 411502
rect 508180 411438 511876 411502
rect 511940 411438 515636 411502
rect 515700 411438 519396 411502
rect 519460 411438 523156 411502
rect 523220 411438 526916 411502
rect 526980 411438 530676 411502
rect 530740 411438 534436 411502
rect 534500 411438 537222 411502
rect 490354 411422 537222 411438
rect 490354 411358 493076 411422
rect 493140 411358 496836 411422
rect 496900 411358 500596 411422
rect 500660 411358 504356 411422
rect 504420 411358 508116 411422
rect 508180 411358 511876 411422
rect 511940 411358 515636 411422
rect 515700 411358 519396 411422
rect 519460 411358 523156 411422
rect 523220 411358 526916 411422
rect 526980 411358 530676 411422
rect 530740 411358 534436 411422
rect 534500 411358 537222 411422
rect 490354 411342 537222 411358
rect 490354 411278 493076 411342
rect 493140 411278 496836 411342
rect 496900 411278 500596 411342
rect 500660 411278 504356 411342
rect 504420 411278 508116 411342
rect 508180 411278 511876 411342
rect 511940 411278 515636 411342
rect 515700 411278 519396 411342
rect 519460 411278 523156 411342
rect 523220 411278 526916 411342
rect 526980 411278 530676 411342
rect 530740 411278 534436 411342
rect 534500 411278 537222 411342
rect 490354 411262 537222 411278
rect 490354 411198 493076 411262
rect 493140 411198 496836 411262
rect 496900 411198 500596 411262
rect 500660 411198 504356 411262
rect 504420 411198 508116 411262
rect 508180 411198 511876 411262
rect 511940 411198 515636 411262
rect 515700 411198 519396 411262
rect 519460 411198 523156 411262
rect 523220 411198 526916 411262
rect 526980 411198 530676 411262
rect 530740 411198 534436 411262
rect 534500 411198 537222 411262
rect 490354 411182 537222 411198
rect 490354 411118 493076 411182
rect 493140 411118 496836 411182
rect 496900 411118 500596 411182
rect 500660 411118 504356 411182
rect 504420 411118 508116 411182
rect 508180 411118 511876 411182
rect 511940 411118 515636 411182
rect 515700 411118 519396 411182
rect 519460 411118 523156 411182
rect 523220 411118 526916 411182
rect 526980 411118 530676 411182
rect 530740 411118 534436 411182
rect 534500 411118 537222 411182
rect 490354 411102 537222 411118
rect 490354 411038 493076 411102
rect 493140 411038 496836 411102
rect 496900 411038 500596 411102
rect 500660 411038 504356 411102
rect 504420 411038 508116 411102
rect 508180 411038 511876 411102
rect 511940 411038 515636 411102
rect 515700 411038 519396 411102
rect 519460 411038 523156 411102
rect 523220 411038 526916 411102
rect 526980 411038 530676 411102
rect 530740 411038 534436 411102
rect 534500 411038 537222 411102
rect 490354 411022 537222 411038
rect 490354 410958 493076 411022
rect 493140 410958 496836 411022
rect 496900 410958 500596 411022
rect 500660 410958 504356 411022
rect 504420 410958 508116 411022
rect 508180 410958 511876 411022
rect 511940 410958 515636 411022
rect 515700 410958 519396 411022
rect 519460 410958 523156 411022
rect 523220 410958 526916 411022
rect 526980 410958 530676 411022
rect 530740 410958 534436 411022
rect 534500 410958 537222 411022
rect 490354 410942 537222 410958
rect 490354 410878 493076 410942
rect 493140 410878 496836 410942
rect 496900 410878 500596 410942
rect 500660 410878 504356 410942
rect 504420 410878 508116 410942
rect 508180 410878 511876 410942
rect 511940 410878 515636 410942
rect 515700 410878 519396 410942
rect 519460 410878 523156 410942
rect 523220 410878 526916 410942
rect 526980 410878 530676 410942
rect 530740 410878 534436 410942
rect 534500 410878 537222 410942
rect 490354 410862 537222 410878
rect 490354 410798 493076 410862
rect 493140 410798 496836 410862
rect 496900 410798 500596 410862
rect 500660 410798 504356 410862
rect 504420 410798 508116 410862
rect 508180 410798 511876 410862
rect 511940 410798 515636 410862
rect 515700 410798 519396 410862
rect 519460 410798 523156 410862
rect 523220 410798 526916 410862
rect 526980 410798 530676 410862
rect 530740 410798 534436 410862
rect 534500 410798 537222 410862
rect 490354 410782 537222 410798
rect 490354 410718 493076 410782
rect 493140 410718 496836 410782
rect 496900 410718 500596 410782
rect 500660 410718 504356 410782
rect 504420 410718 508116 410782
rect 508180 410718 511876 410782
rect 511940 410718 515636 410782
rect 515700 410718 519396 410782
rect 519460 410718 523156 410782
rect 523220 410718 526916 410782
rect 526980 410718 530676 410782
rect 530740 410718 534436 410782
rect 534500 410718 537222 410782
rect 490354 410702 537222 410718
rect 490354 410638 493076 410702
rect 493140 410638 496836 410702
rect 496900 410638 500596 410702
rect 500660 410638 504356 410702
rect 504420 410638 508116 410702
rect 508180 410638 511876 410702
rect 511940 410638 515636 410702
rect 515700 410638 519396 410702
rect 519460 410638 523156 410702
rect 523220 410638 526916 410702
rect 526980 410638 530676 410702
rect 530740 410638 534436 410702
rect 534500 410638 537222 410702
rect 490354 410622 537222 410638
rect 490354 410558 493076 410622
rect 493140 410558 496836 410622
rect 496900 410558 500596 410622
rect 500660 410558 504356 410622
rect 504420 410558 508116 410622
rect 508180 410558 511876 410622
rect 511940 410558 515636 410622
rect 515700 410558 519396 410622
rect 519460 410558 523156 410622
rect 523220 410558 526916 410622
rect 526980 410558 530676 410622
rect 530740 410558 534436 410622
rect 534500 410558 537222 410622
rect 490354 410542 537222 410558
rect 490354 410478 493076 410542
rect 493140 410478 496836 410542
rect 496900 410478 500596 410542
rect 500660 410478 504356 410542
rect 504420 410478 508116 410542
rect 508180 410478 511876 410542
rect 511940 410478 515636 410542
rect 515700 410478 519396 410542
rect 519460 410478 523156 410542
rect 523220 410478 526916 410542
rect 526980 410478 530676 410542
rect 530740 410478 534436 410542
rect 534500 410478 537222 410542
rect 490354 410462 537222 410478
rect 490354 410398 493076 410462
rect 493140 410398 496836 410462
rect 496900 410398 500596 410462
rect 500660 410398 504356 410462
rect 504420 410398 508116 410462
rect 508180 410398 511876 410462
rect 511940 410398 515636 410462
rect 515700 410398 519396 410462
rect 519460 410398 523156 410462
rect 523220 410398 526916 410462
rect 526980 410398 530676 410462
rect 530740 410398 534436 410462
rect 534500 410398 537222 410462
rect 490354 410382 537222 410398
rect 490354 410318 493076 410382
rect 493140 410318 496836 410382
rect 496900 410318 500596 410382
rect 500660 410318 504356 410382
rect 504420 410318 508116 410382
rect 508180 410318 511876 410382
rect 511940 410318 515636 410382
rect 515700 410318 519396 410382
rect 519460 410318 523156 410382
rect 523220 410318 526916 410382
rect 526980 410318 530676 410382
rect 530740 410318 534436 410382
rect 534500 410318 537222 410382
rect 490354 410302 537222 410318
rect 490354 410238 493076 410302
rect 493140 410238 496836 410302
rect 496900 410238 500596 410302
rect 500660 410238 504356 410302
rect 504420 410238 508116 410302
rect 508180 410238 511876 410302
rect 511940 410238 515636 410302
rect 515700 410238 519396 410302
rect 519460 410238 523156 410302
rect 523220 410238 526916 410302
rect 526980 410238 530676 410302
rect 530740 410238 534436 410302
rect 534500 410238 537222 410302
rect 490354 410222 537222 410238
rect 490354 410158 493076 410222
rect 493140 410158 496836 410222
rect 496900 410158 500596 410222
rect 500660 410158 504356 410222
rect 504420 410158 508116 410222
rect 508180 410158 511876 410222
rect 511940 410158 515636 410222
rect 515700 410158 519396 410222
rect 519460 410158 523156 410222
rect 523220 410158 526916 410222
rect 526980 410158 530676 410222
rect 530740 410158 534436 410222
rect 534500 410158 537222 410222
rect 490354 410142 537222 410158
rect 490354 410078 493076 410142
rect 493140 410078 496836 410142
rect 496900 410078 500596 410142
rect 500660 410078 504356 410142
rect 504420 410078 508116 410142
rect 508180 410078 511876 410142
rect 511940 410078 515636 410142
rect 515700 410078 519396 410142
rect 519460 410078 523156 410142
rect 523220 410078 526916 410142
rect 526980 410078 530676 410142
rect 530740 410078 534436 410142
rect 534500 410078 537222 410142
rect 490354 410062 537222 410078
rect 490354 410032 493076 410062
rect 485484 409998 493076 410032
rect 493140 409998 496836 410062
rect 496900 409998 500596 410062
rect 500660 409998 504356 410062
rect 504420 409998 508116 410062
rect 508180 409998 511876 410062
rect 511940 409998 515636 410062
rect 515700 409998 519396 410062
rect 519460 409998 523156 410062
rect 523220 409998 526916 410062
rect 526980 409998 530676 410062
rect 530740 409998 534436 410062
rect 534500 410032 537222 410062
rect 538738 410032 542060 411548
rect 534500 409998 542060 410032
rect 485484 409974 542060 409998
rect 493096 409220 496816 409280
rect 493096 408418 493156 409220
rect 494738 409008 494858 409036
rect 494738 408944 494766 409008
rect 494830 408944 494858 409008
rect 494738 408928 494858 408944
rect 494738 408898 494766 408928
rect 493458 408889 494766 408898
rect 493458 408585 493486 408889
rect 493790 408585 494186 408889
rect 494490 408864 494766 408889
rect 494830 408864 494858 408928
rect 494490 408585 494858 408864
rect 493458 408578 494858 408585
rect 493477 408576 493799 408578
rect 494177 408576 494499 408578
rect 493350 408422 493926 408438
rect 493350 408418 493366 408422
rect 493096 408358 493366 408418
rect 493430 408358 493446 408422
rect 493510 408358 493526 408422
rect 493590 408358 493606 408422
rect 493670 408358 493686 408422
rect 493750 408358 493766 408422
rect 493830 408358 493846 408422
rect 493910 408358 493926 408422
rect 493350 408342 493926 408358
rect 494050 408422 494626 408438
rect 494050 408358 494066 408422
rect 494130 408358 494146 408422
rect 494210 408358 494226 408422
rect 494290 408358 494306 408422
rect 494370 408358 494386 408422
rect 494450 408358 494466 408422
rect 494530 408358 494546 408422
rect 494610 408358 494626 408422
rect 494050 408342 494626 408358
rect 493477 408178 493799 408179
rect 494177 408178 494499 408179
rect 494738 408178 494858 408578
rect 496756 408418 496816 409220
rect 498498 409008 498618 409036
rect 498498 408944 498526 409008
rect 498590 408944 498618 409008
rect 498498 408928 498618 408944
rect 498498 408898 498526 408928
rect 497218 408889 498526 408898
rect 497218 408585 497246 408889
rect 497550 408585 497946 408889
rect 498250 408864 498526 408889
rect 498590 408864 498618 408928
rect 498250 408585 498618 408864
rect 497218 408578 498618 408585
rect 497237 408576 497559 408578
rect 497937 408576 498259 408578
rect 497110 408422 497686 408438
rect 497110 408418 497126 408422
rect 496756 408358 497126 408418
rect 497190 408358 497206 408422
rect 497270 408358 497286 408422
rect 497350 408358 497366 408422
rect 497430 408358 497446 408422
rect 497510 408358 497526 408422
rect 497590 408358 497606 408422
rect 497670 408358 497686 408422
rect 497110 408342 497686 408358
rect 497810 408422 498386 408438
rect 497810 408358 497826 408422
rect 497890 408358 497906 408422
rect 497970 408358 497986 408422
rect 498050 408358 498066 408422
rect 498130 408358 498146 408422
rect 498210 408358 498226 408422
rect 498290 408358 498306 408422
rect 498370 408358 498386 408422
rect 497810 408342 498386 408358
rect 498498 408314 498618 408578
rect 502258 408616 502378 408644
rect 502258 408552 502286 408616
rect 502350 408552 502378 408616
rect 502258 408536 502378 408552
rect 502258 408506 502286 408536
rect 500978 408497 502286 408506
rect 500978 408314 501006 408497
rect 498498 408254 501006 408314
rect 497237 408178 497559 408179
rect 497937 408178 498259 408179
rect 498498 408178 498618 408254
rect 500978 408193 501006 408254
rect 501310 408193 501706 408497
rect 502010 408472 502286 408497
rect 502350 408472 502378 408536
rect 502010 408193 502378 408472
rect 500978 408186 502378 408193
rect 500997 408184 501319 408186
rect 501697 408184 502019 408186
rect 493458 408170 494858 408178
rect 493458 407866 493486 408170
rect 493790 407866 494186 408170
rect 494490 407866 494858 408170
rect 493458 407858 494858 407866
rect 497218 408170 498618 408178
rect 497218 407866 497246 408170
rect 497550 407866 497946 408170
rect 498250 407866 498618 408170
rect 500657 408040 500723 408041
rect 500657 407976 500658 408040
rect 500722 408038 500723 408040
rect 500870 408038 501446 408046
rect 500722 408030 501446 408038
rect 500722 407978 500886 408030
rect 500722 407976 500723 407978
rect 500657 407975 500723 407976
rect 500870 407966 500886 407978
rect 500950 407966 500966 408030
rect 501030 407966 501046 408030
rect 501110 407966 501126 408030
rect 501190 407966 501206 408030
rect 501270 407966 501286 408030
rect 501350 407966 501366 408030
rect 501430 407966 501446 408030
rect 500870 407950 501446 407966
rect 501570 408030 502146 408046
rect 501570 407966 501586 408030
rect 501650 407966 501666 408030
rect 501730 407966 501746 408030
rect 501810 407966 501826 408030
rect 501890 407966 501906 408030
rect 501970 407966 501986 408030
rect 502050 407966 502066 408030
rect 502130 407966 502146 408030
rect 501570 407950 502146 407966
rect 497218 407858 498618 407866
rect 493477 407857 493799 407858
rect 494177 407857 494499 407858
rect 493350 407703 493926 407719
rect 493350 407639 493366 407703
rect 493430 407639 493446 407703
rect 493510 407639 493526 407703
rect 493590 407639 493606 407703
rect 493670 407639 493686 407703
rect 493750 407639 493766 407703
rect 493830 407639 493846 407703
rect 493910 407639 493926 407703
rect 493350 407623 493926 407639
rect 494050 407703 494626 407719
rect 494050 407639 494066 407703
rect 494130 407639 494146 407703
rect 494210 407639 494226 407703
rect 494290 407639 494306 407703
rect 494370 407639 494386 407703
rect 494450 407639 494466 407703
rect 494530 407639 494546 407703
rect 494610 407639 494626 407703
rect 494050 407623 494626 407639
rect 493477 407458 493799 407460
rect 494177 407458 494499 407460
rect 494738 407458 494858 407858
rect 497237 407857 497559 407858
rect 497937 407857 498259 407858
rect 497110 407703 497686 407719
rect 497110 407639 497126 407703
rect 497190 407639 497206 407703
rect 497270 407639 497286 407703
rect 497350 407639 497366 407703
rect 497430 407639 497446 407703
rect 497510 407639 497526 407703
rect 497590 407639 497606 407703
rect 497670 407639 497686 407703
rect 497110 407623 497686 407639
rect 497810 407703 498386 407719
rect 497810 407639 497826 407703
rect 497890 407639 497906 407703
rect 497970 407639 497986 407703
rect 498050 407639 498066 407703
rect 498130 407639 498146 407703
rect 498210 407639 498226 407703
rect 498290 407639 498306 407703
rect 498370 407639 498386 407703
rect 497810 407623 498386 407639
rect 497237 407458 497559 407460
rect 497937 407458 498259 407460
rect 498498 407458 498618 407858
rect 500997 407786 501319 407787
rect 501697 407786 502019 407787
rect 502258 407786 502378 408186
rect 500978 407778 502378 407786
rect 500978 407474 501006 407778
rect 501310 407474 501706 407778
rect 502010 407474 502378 407778
rect 500978 407466 502378 407474
rect 500997 407465 501319 407466
rect 501697 407465 502019 407466
rect 493458 407451 494858 407458
rect 493458 407147 493486 407451
rect 493790 407147 494186 407451
rect 494490 407147 494858 407451
rect 493458 407138 494858 407147
rect 497218 407451 498618 407458
rect 497218 407147 497246 407451
rect 497550 407147 497946 407451
rect 498250 407147 498618 407451
rect 500870 407311 501446 407327
rect 500870 407247 500886 407311
rect 500950 407247 500966 407311
rect 501030 407247 501046 407311
rect 501110 407247 501126 407311
rect 501190 407247 501206 407311
rect 501270 407247 501286 407311
rect 501350 407247 501366 407311
rect 501430 407247 501446 407311
rect 500870 407231 501446 407247
rect 501570 407311 502146 407327
rect 501570 407247 501586 407311
rect 501650 407247 501666 407311
rect 501730 407247 501746 407311
rect 501810 407247 501826 407311
rect 501890 407247 501906 407311
rect 501970 407247 501986 407311
rect 502050 407247 502066 407311
rect 502130 407247 502146 407311
rect 501570 407231 502146 407247
rect 497218 407138 498618 407147
rect 493350 406984 493926 407000
rect 493350 406920 493366 406984
rect 493430 406920 493446 406984
rect 493510 406920 493526 406984
rect 493590 406920 493606 406984
rect 493670 406920 493686 406984
rect 493750 406920 493766 406984
rect 493830 406920 493846 406984
rect 493910 406920 493926 406984
rect 493350 406904 493926 406920
rect 494050 406984 494626 407000
rect 494050 406920 494066 406984
rect 494130 406920 494146 406984
rect 494210 406920 494226 406984
rect 494290 406920 494306 406984
rect 494370 406920 494386 406984
rect 494450 406920 494466 406984
rect 494530 406920 494546 406984
rect 494610 406920 494626 406984
rect 494050 406904 494626 406920
rect 493477 406738 493799 406741
rect 494177 406738 494499 406741
rect 494738 406738 494858 407138
rect 497110 406984 497686 407000
rect 497110 406920 497126 406984
rect 497190 406920 497206 406984
rect 497270 406920 497286 406984
rect 497350 406920 497366 406984
rect 497430 406920 497446 406984
rect 497510 406920 497526 406984
rect 497590 406920 497606 406984
rect 497670 406920 497686 406984
rect 497110 406904 497686 406920
rect 497810 406984 498386 407000
rect 497810 406920 497826 406984
rect 497890 406920 497906 406984
rect 497970 406920 497986 406984
rect 498050 406920 498066 406984
rect 498130 406920 498146 406984
rect 498210 406920 498226 406984
rect 498290 406920 498306 406984
rect 498370 406920 498386 406984
rect 497810 406904 498386 406920
rect 497237 406738 497559 406741
rect 497937 406738 498259 406741
rect 498498 406738 498618 407138
rect 500997 407066 501319 407068
rect 501697 407066 502019 407068
rect 502258 407066 502378 407466
rect 500978 407059 502378 407066
rect 500978 406755 501006 407059
rect 501310 406755 501706 407059
rect 502010 406755 502378 407059
rect 500978 406746 502378 406755
rect 493458 406732 494858 406738
rect 493458 406428 493486 406732
rect 493790 406428 494186 406732
rect 494490 406428 494858 406732
rect 493458 406418 494858 406428
rect 497218 406732 498618 406738
rect 497218 406428 497246 406732
rect 497550 406428 497946 406732
rect 498250 406658 498618 406732
rect 498705 406660 498771 406661
rect 498705 406658 498706 406660
rect 498250 406598 498706 406658
rect 498250 406428 498618 406598
rect 498705 406596 498706 406598
rect 498770 406596 498771 406660
rect 498705 406595 498771 406596
rect 500870 406592 501446 406608
rect 500870 406528 500886 406592
rect 500950 406528 500966 406592
rect 501030 406528 501046 406592
rect 501110 406528 501126 406592
rect 501190 406528 501206 406592
rect 501270 406528 501286 406592
rect 501350 406528 501366 406592
rect 501430 406528 501446 406592
rect 500870 406512 501446 406528
rect 501570 406592 502146 406608
rect 501570 406528 501586 406592
rect 501650 406528 501666 406592
rect 501730 406528 501746 406592
rect 501810 406528 501826 406592
rect 501890 406528 501906 406592
rect 501970 406528 501986 406592
rect 502050 406528 502066 406592
rect 502130 406528 502146 406592
rect 501570 406512 502146 406528
rect 497218 406418 498618 406428
rect 493350 406265 493926 406281
rect 493350 406201 493366 406265
rect 493430 406201 493446 406265
rect 493510 406201 493526 406265
rect 493590 406201 493606 406265
rect 493670 406201 493686 406265
rect 493750 406201 493766 406265
rect 493830 406201 493846 406265
rect 493910 406201 493926 406265
rect 493350 406185 493926 406201
rect 494050 406265 494626 406281
rect 494050 406201 494066 406265
rect 494130 406201 494146 406265
rect 494210 406201 494226 406265
rect 494290 406201 494306 406265
rect 494370 406201 494386 406265
rect 494450 406201 494466 406265
rect 494530 406201 494546 406265
rect 494610 406201 494626 406265
rect 494050 406185 494626 406201
rect 493477 406018 493799 406022
rect 494177 406018 494499 406022
rect 494738 406018 494858 406418
rect 497110 406265 497686 406281
rect 497110 406201 497126 406265
rect 497190 406201 497206 406265
rect 497270 406201 497286 406265
rect 497350 406201 497366 406265
rect 497430 406201 497446 406265
rect 497510 406201 497526 406265
rect 497590 406201 497606 406265
rect 497670 406201 497686 406265
rect 497110 406185 497686 406201
rect 497810 406265 498386 406281
rect 497810 406201 497826 406265
rect 497890 406201 497906 406265
rect 497970 406201 497986 406265
rect 498050 406201 498066 406265
rect 498130 406201 498146 406265
rect 498210 406201 498226 406265
rect 498290 406201 498306 406265
rect 498370 406201 498386 406265
rect 497810 406185 498386 406201
rect 497237 406018 497559 406022
rect 497937 406018 498259 406022
rect 498498 406018 498618 406418
rect 500997 406346 501319 406349
rect 501697 406346 502019 406349
rect 502258 406346 502378 406746
rect 500978 406340 502378 406346
rect 500978 406036 501006 406340
rect 501310 406036 501706 406340
rect 502010 406036 502378 406340
rect 500978 406026 502378 406036
rect 493458 406013 494858 406018
rect 493458 405709 493486 406013
rect 493790 405709 494186 406013
rect 494490 405709 494858 406013
rect 493458 405698 494858 405709
rect 497218 406013 498618 406018
rect 497218 405709 497246 406013
rect 497550 405709 497946 406013
rect 498250 405709 498618 406013
rect 500870 405873 501446 405889
rect 500870 405809 500886 405873
rect 500950 405809 500966 405873
rect 501030 405809 501046 405873
rect 501110 405809 501126 405873
rect 501190 405809 501206 405873
rect 501270 405809 501286 405873
rect 501350 405809 501366 405873
rect 501430 405809 501446 405873
rect 500870 405793 501446 405809
rect 501570 405873 502146 405889
rect 501570 405809 501586 405873
rect 501650 405809 501666 405873
rect 501730 405809 501746 405873
rect 501810 405809 501826 405873
rect 501890 405809 501906 405873
rect 501970 405809 501986 405873
rect 502050 405809 502066 405873
rect 502130 405809 502146 405873
rect 501570 405793 502146 405809
rect 497218 405698 498618 405709
rect 493350 405546 493926 405562
rect 493350 405482 493366 405546
rect 493430 405482 493446 405546
rect 493510 405482 493526 405546
rect 493590 405482 493606 405546
rect 493670 405482 493686 405546
rect 493750 405482 493766 405546
rect 493830 405482 493846 405546
rect 493910 405482 493926 405546
rect 493350 405466 493926 405482
rect 494050 405546 494626 405562
rect 494050 405482 494066 405546
rect 494130 405482 494146 405546
rect 494210 405482 494226 405546
rect 494290 405482 494306 405546
rect 494370 405482 494386 405546
rect 494450 405482 494466 405546
rect 494530 405482 494546 405546
rect 494610 405482 494626 405546
rect 494050 405466 494626 405482
rect 493477 405298 493799 405303
rect 494177 405298 494499 405303
rect 494738 405298 494858 405698
rect 497110 405546 497686 405562
rect 497110 405482 497126 405546
rect 497190 405482 497206 405546
rect 497270 405482 497286 405546
rect 497350 405482 497366 405546
rect 497430 405482 497446 405546
rect 497510 405482 497526 405546
rect 497590 405482 497606 405546
rect 497670 405482 497686 405546
rect 497110 405466 497686 405482
rect 497810 405546 498386 405562
rect 497810 405482 497826 405546
rect 497890 405482 497906 405546
rect 497970 405482 497986 405546
rect 498050 405482 498066 405546
rect 498130 405482 498146 405546
rect 498210 405482 498226 405546
rect 498290 405482 498306 405546
rect 498370 405482 498386 405546
rect 497810 405466 498386 405482
rect 497237 405298 497559 405303
rect 497937 405298 498259 405303
rect 498498 405298 498618 405698
rect 500997 405626 501319 405630
rect 501697 405626 502019 405630
rect 502258 405626 502378 406026
rect 500978 405621 502378 405626
rect 500978 405317 501006 405621
rect 501310 405317 501706 405621
rect 502010 405317 502378 405621
rect 500978 405306 502378 405317
rect 493458 405294 494858 405298
rect 493458 404990 493486 405294
rect 493790 404990 494186 405294
rect 494490 404990 494858 405294
rect 493458 404978 494858 404990
rect 497218 405294 498618 405298
rect 497218 404990 497246 405294
rect 497550 404990 497946 405294
rect 498250 404990 498618 405294
rect 500870 405154 501446 405170
rect 500870 405090 500886 405154
rect 500950 405090 500966 405154
rect 501030 405090 501046 405154
rect 501110 405090 501126 405154
rect 501190 405090 501206 405154
rect 501270 405090 501286 405154
rect 501350 405090 501366 405154
rect 501430 405090 501446 405154
rect 500870 405074 501446 405090
rect 501570 405154 502146 405170
rect 501570 405090 501586 405154
rect 501650 405090 501666 405154
rect 501730 405090 501746 405154
rect 501810 405090 501826 405154
rect 501890 405090 501906 405154
rect 501970 405090 501986 405154
rect 502050 405090 502066 405154
rect 502130 405090 502146 405154
rect 501570 405074 502146 405090
rect 497218 404978 498618 404990
rect 493350 404827 493926 404843
rect 493350 404763 493366 404827
rect 493430 404763 493446 404827
rect 493510 404763 493526 404827
rect 493590 404763 493606 404827
rect 493670 404763 493686 404827
rect 493750 404763 493766 404827
rect 493830 404763 493846 404827
rect 493910 404763 493926 404827
rect 493350 404747 493926 404763
rect 494050 404827 494626 404843
rect 494050 404763 494066 404827
rect 494130 404763 494146 404827
rect 494210 404763 494226 404827
rect 494290 404763 494306 404827
rect 494370 404763 494386 404827
rect 494450 404763 494466 404827
rect 494530 404763 494546 404827
rect 494610 404763 494626 404827
rect 494050 404747 494626 404763
rect 493477 404578 493799 404584
rect 494177 404578 494499 404584
rect 494738 404578 494858 404978
rect 497110 404827 497686 404843
rect 497110 404763 497126 404827
rect 497190 404763 497206 404827
rect 497270 404763 497286 404827
rect 497350 404763 497366 404827
rect 497430 404763 497446 404827
rect 497510 404763 497526 404827
rect 497590 404763 497606 404827
rect 497670 404763 497686 404827
rect 497110 404747 497686 404763
rect 497810 404827 498386 404843
rect 497810 404763 497826 404827
rect 497890 404763 497906 404827
rect 497970 404763 497986 404827
rect 498050 404763 498066 404827
rect 498130 404763 498146 404827
rect 498210 404763 498226 404827
rect 498290 404763 498306 404827
rect 498370 404763 498386 404827
rect 497810 404747 498386 404763
rect 497237 404578 497559 404584
rect 497937 404578 498259 404584
rect 498498 404578 498618 404978
rect 500997 404906 501319 404911
rect 501697 404906 502019 404911
rect 502258 404906 502378 405306
rect 500978 404902 502378 404906
rect 500978 404598 501006 404902
rect 501310 404598 501706 404902
rect 502010 404598 502378 404902
rect 500978 404586 502378 404598
rect 493458 404575 494858 404578
rect 493458 404271 493486 404575
rect 493790 404271 494186 404575
rect 494490 404271 494858 404575
rect 493458 404258 494858 404271
rect 497218 404575 498618 404578
rect 497218 404271 497246 404575
rect 497550 404271 497946 404575
rect 498250 404271 498618 404575
rect 500870 404435 501446 404451
rect 500870 404371 500886 404435
rect 500950 404371 500966 404435
rect 501030 404371 501046 404435
rect 501110 404371 501126 404435
rect 501190 404371 501206 404435
rect 501270 404371 501286 404435
rect 501350 404371 501366 404435
rect 501430 404371 501446 404435
rect 500870 404355 501446 404371
rect 501570 404435 502146 404451
rect 501570 404371 501586 404435
rect 501650 404371 501666 404435
rect 501730 404371 501746 404435
rect 501810 404371 501826 404435
rect 501890 404371 501906 404435
rect 501970 404371 501986 404435
rect 502050 404371 502066 404435
rect 502130 404371 502146 404435
rect 501570 404355 502146 404371
rect 497218 404258 498618 404271
rect 493350 404108 493926 404124
rect 493350 404044 493366 404108
rect 493430 404044 493446 404108
rect 493510 404044 493526 404108
rect 493590 404044 493606 404108
rect 493670 404044 493686 404108
rect 493750 404044 493766 404108
rect 493830 404044 493846 404108
rect 493910 404044 493926 404108
rect 493350 404028 493926 404044
rect 494050 404108 494626 404124
rect 494050 404044 494066 404108
rect 494130 404044 494146 404108
rect 494210 404044 494226 404108
rect 494290 404044 494306 404108
rect 494370 404044 494386 404108
rect 494450 404044 494466 404108
rect 494530 404044 494546 404108
rect 494610 404044 494626 404108
rect 494050 404028 494626 404044
rect 493477 403858 493799 403865
rect 494177 403858 494499 403865
rect 494738 403858 494858 404258
rect 497110 404108 497686 404124
rect 497110 404044 497126 404108
rect 497190 404044 497206 404108
rect 497270 404044 497286 404108
rect 497350 404044 497366 404108
rect 497430 404044 497446 404108
rect 497510 404044 497526 404108
rect 497590 404044 497606 404108
rect 497670 404044 497686 404108
rect 497110 404028 497686 404044
rect 497810 404108 498386 404124
rect 497810 404044 497826 404108
rect 497890 404044 497906 404108
rect 497970 404044 497986 404108
rect 498050 404044 498066 404108
rect 498130 404044 498146 404108
rect 498210 404044 498226 404108
rect 498290 404044 498306 404108
rect 498370 404044 498386 404108
rect 497810 404028 498386 404044
rect 497237 403858 497559 403865
rect 497937 403858 498259 403865
rect 498498 403858 498618 404258
rect 500997 404186 501319 404192
rect 501697 404186 502019 404192
rect 502258 404186 502378 404586
rect 500978 404183 502378 404186
rect 500978 403879 501006 404183
rect 501310 403879 501706 404183
rect 502010 403879 502378 404183
rect 500978 403866 502378 403879
rect 493458 403856 494858 403858
rect 493458 403552 493486 403856
rect 493790 403552 494186 403856
rect 494490 403552 494858 403856
rect 493458 403538 494858 403552
rect 497218 403856 498618 403858
rect 497218 403552 497246 403856
rect 497550 403552 497946 403856
rect 498250 403552 498618 403856
rect 500870 403716 501446 403732
rect 500870 403652 500886 403716
rect 500950 403652 500966 403716
rect 501030 403652 501046 403716
rect 501110 403652 501126 403716
rect 501190 403652 501206 403716
rect 501270 403652 501286 403716
rect 501350 403652 501366 403716
rect 501430 403652 501446 403716
rect 500870 403636 501446 403652
rect 501570 403716 502146 403732
rect 501570 403652 501586 403716
rect 501650 403652 501666 403716
rect 501730 403652 501746 403716
rect 501810 403652 501826 403716
rect 501890 403652 501906 403716
rect 501970 403652 501986 403716
rect 502050 403652 502066 403716
rect 502130 403652 502146 403716
rect 501570 403636 502146 403652
rect 497218 403538 498618 403552
rect 493350 403389 493926 403405
rect 493350 403325 493366 403389
rect 493430 403325 493446 403389
rect 493510 403325 493526 403389
rect 493590 403325 493606 403389
rect 493670 403325 493686 403389
rect 493750 403325 493766 403389
rect 493830 403325 493846 403389
rect 493910 403325 493926 403389
rect 493350 403309 493926 403325
rect 494050 403389 494626 403405
rect 494050 403325 494066 403389
rect 494130 403325 494146 403389
rect 494210 403325 494226 403389
rect 494290 403325 494306 403389
rect 494370 403325 494386 403389
rect 494450 403325 494466 403389
rect 494530 403325 494546 403389
rect 494610 403325 494626 403389
rect 494050 403309 494626 403325
rect 493477 403138 493799 403146
rect 494177 403138 494499 403146
rect 494738 403138 494858 403538
rect 497110 403389 497686 403405
rect 497110 403325 497126 403389
rect 497190 403325 497206 403389
rect 497270 403325 497286 403389
rect 497350 403325 497366 403389
rect 497430 403325 497446 403389
rect 497510 403325 497526 403389
rect 497590 403325 497606 403389
rect 497670 403325 497686 403389
rect 497110 403309 497686 403325
rect 497810 403389 498386 403405
rect 497810 403325 497826 403389
rect 497890 403325 497906 403389
rect 497970 403325 497986 403389
rect 498050 403325 498066 403389
rect 498130 403325 498146 403389
rect 498210 403325 498226 403389
rect 498290 403325 498306 403389
rect 498370 403325 498386 403389
rect 497810 403309 498386 403325
rect 497237 403138 497559 403146
rect 497937 403138 498259 403146
rect 498498 403138 498618 403538
rect 500997 403466 501319 403473
rect 501697 403466 502019 403473
rect 502258 403466 502378 403866
rect 500978 403464 502378 403466
rect 500978 403160 501006 403464
rect 501310 403160 501706 403464
rect 502010 403160 502378 403464
rect 500978 403146 502378 403160
rect 493458 403137 494858 403138
rect 493458 402833 493486 403137
rect 493790 402833 494186 403137
rect 494490 402833 494858 403137
rect 493458 402818 494858 402833
rect 497218 403137 498618 403138
rect 497218 402833 497246 403137
rect 497550 402833 497946 403137
rect 498250 402833 498618 403137
rect 500870 402997 501446 403013
rect 500870 402933 500886 402997
rect 500950 402933 500966 402997
rect 501030 402933 501046 402997
rect 501110 402933 501126 402997
rect 501190 402933 501206 402997
rect 501270 402933 501286 402997
rect 501350 402933 501366 402997
rect 501430 402933 501446 402997
rect 500870 402917 501446 402933
rect 501570 402997 502146 403013
rect 501570 402933 501586 402997
rect 501650 402933 501666 402997
rect 501730 402933 501746 402997
rect 501810 402933 501826 402997
rect 501890 402933 501906 402997
rect 501970 402933 501986 402997
rect 502050 402933 502066 402997
rect 502130 402933 502146 402997
rect 501570 402917 502146 402933
rect 497218 402818 498618 402833
rect 493350 402670 493926 402686
rect 493350 402606 493366 402670
rect 493430 402606 493446 402670
rect 493510 402606 493526 402670
rect 493590 402606 493606 402670
rect 493670 402606 493686 402670
rect 493750 402606 493766 402670
rect 493830 402606 493846 402670
rect 493910 402606 493926 402670
rect 493350 402590 493926 402606
rect 494050 402670 494626 402686
rect 494050 402606 494066 402670
rect 494130 402606 494146 402670
rect 494210 402606 494226 402670
rect 494290 402606 494306 402670
rect 494370 402606 494386 402670
rect 494450 402606 494466 402670
rect 494530 402606 494546 402670
rect 494610 402606 494626 402670
rect 494050 402590 494626 402606
rect 493477 402418 493799 402427
rect 494177 402418 494499 402427
rect 494738 402418 494858 402818
rect 497110 402670 497686 402686
rect 497110 402606 497126 402670
rect 497190 402606 497206 402670
rect 497270 402606 497286 402670
rect 497350 402606 497366 402670
rect 497430 402606 497446 402670
rect 497510 402606 497526 402670
rect 497590 402606 497606 402670
rect 497670 402606 497686 402670
rect 497110 402590 497686 402606
rect 497810 402670 498386 402686
rect 497810 402606 497826 402670
rect 497890 402606 497906 402670
rect 497970 402606 497986 402670
rect 498050 402606 498066 402670
rect 498130 402606 498146 402670
rect 498210 402606 498226 402670
rect 498290 402606 498306 402670
rect 498370 402606 498386 402670
rect 497810 402590 498386 402606
rect 497237 402418 497559 402427
rect 497937 402418 498259 402427
rect 498498 402418 498618 402818
rect 500997 402746 501319 402754
rect 501697 402746 502019 402754
rect 502258 402746 502378 403146
rect 500978 402745 502378 402746
rect 500978 402441 501006 402745
rect 501310 402441 501706 402745
rect 502010 402441 502378 402745
rect 500978 402426 502378 402441
rect 493458 402114 493486 402418
rect 493790 402114 494186 402418
rect 494490 402114 494858 402418
rect 493458 402098 494858 402114
rect 497218 402114 497246 402418
rect 497550 402114 497946 402418
rect 498250 402114 498618 402418
rect 500870 402278 501446 402294
rect 500870 402214 500886 402278
rect 500950 402214 500966 402278
rect 501030 402214 501046 402278
rect 501110 402214 501126 402278
rect 501190 402214 501206 402278
rect 501270 402214 501286 402278
rect 501350 402214 501366 402278
rect 501430 402214 501446 402278
rect 500870 402198 501446 402214
rect 501570 402278 502146 402294
rect 501570 402214 501586 402278
rect 501650 402214 501666 402278
rect 501730 402214 501746 402278
rect 501810 402214 501826 402278
rect 501890 402214 501906 402278
rect 501970 402214 501986 402278
rect 502050 402214 502066 402278
rect 502130 402214 502146 402278
rect 501570 402198 502146 402214
rect 497218 402098 498618 402114
rect 493350 401966 493926 401967
rect 493096 401951 493926 401966
rect 493096 401906 493366 401951
rect 493096 400966 493156 401906
rect 493350 401887 493366 401906
rect 493430 401887 493446 401951
rect 493510 401887 493526 401951
rect 493590 401887 493606 401951
rect 493670 401887 493686 401951
rect 493750 401887 493766 401951
rect 493830 401887 493846 401951
rect 493910 401887 493926 401951
rect 493350 401871 493926 401887
rect 494050 401951 494626 401967
rect 494050 401887 494066 401951
rect 494130 401887 494146 401951
rect 494210 401887 494226 401951
rect 494290 401887 494306 401951
rect 494370 401887 494386 401951
rect 494450 401887 494466 401951
rect 494530 401887 494546 401951
rect 494610 401887 494626 401951
rect 494050 401871 494626 401887
rect 494738 401966 494858 402098
rect 494738 401906 495108 401966
rect 494738 401868 494858 401906
rect 494738 401560 494858 401588
rect 494738 401496 494766 401560
rect 494830 401552 494858 401560
rect 495048 401552 495108 401906
rect 497110 401951 497686 401967
rect 497110 401887 497126 401951
rect 497190 401887 497206 401951
rect 497270 401887 497286 401951
rect 497350 401887 497366 401951
rect 497430 401887 497446 401951
rect 497510 401887 497526 401951
rect 497590 401887 497606 401951
rect 497670 401887 497686 401951
rect 497110 401871 497686 401887
rect 497810 401951 498386 401967
rect 497810 401887 497826 401951
rect 497890 401887 497906 401951
rect 497970 401887 497986 401951
rect 498050 401887 498066 401951
rect 498130 401887 498146 401951
rect 498210 401887 498226 401951
rect 498290 401887 498306 401951
rect 498370 401887 498386 401951
rect 497810 401871 498386 401887
rect 498220 401555 498280 401871
rect 498498 401868 498618 402098
rect 500997 402026 501319 402035
rect 501697 402026 502019 402035
rect 502258 402026 502378 402426
rect 500978 401722 501006 402026
rect 501310 401722 501706 402026
rect 502010 401722 502378 402026
rect 500978 401706 502378 401722
rect 500870 401559 501446 401575
rect 494830 401496 495108 401552
rect 494738 401492 495108 401496
rect 498217 401554 498283 401555
rect 494738 401480 494858 401492
rect 498217 401490 498218 401554
rect 498282 401552 498283 401554
rect 500870 401552 500886 401559
rect 498282 401495 500886 401552
rect 500950 401495 500966 401559
rect 501030 401495 501046 401559
rect 501110 401495 501126 401559
rect 501190 401495 501206 401559
rect 501270 401495 501286 401559
rect 501350 401495 501366 401559
rect 501430 401495 501446 401559
rect 498282 401492 501446 401495
rect 498282 401490 498283 401492
rect 498217 401489 498283 401490
rect 494738 401450 494766 401480
rect 493458 401441 494766 401450
rect 493458 401137 493486 401441
rect 493790 401137 494186 401441
rect 494490 401416 494766 401441
rect 494830 401416 494858 401480
rect 500870 401479 501446 401492
rect 501570 401559 502146 401575
rect 501570 401495 501586 401559
rect 501650 401495 501666 401559
rect 501730 401495 501746 401559
rect 501810 401495 501826 401559
rect 501890 401495 501906 401559
rect 501970 401495 501986 401559
rect 502050 401495 502066 401559
rect 502130 401552 502146 401559
rect 502130 401495 502184 401552
rect 501570 401479 502184 401495
rect 494490 401137 494858 401416
rect 502124 401414 502184 401479
rect 502258 401476 502378 401706
rect 551974 403368 560022 412422
rect 551974 403192 559736 403368
rect 559926 403192 560022 403368
rect 504805 401416 504871 401417
rect 504805 401414 504806 401416
rect 502124 401354 504806 401414
rect 504805 401352 504806 401354
rect 504870 401352 504871 401416
rect 504805 401351 504871 401352
rect 493458 401130 494858 401137
rect 493477 401128 493799 401130
rect 494177 401128 494499 401130
rect 493350 400974 493926 400990
rect 493350 400966 493366 400974
rect 493096 400910 493366 400966
rect 493430 400910 493446 400974
rect 493510 400910 493526 400974
rect 493590 400910 493606 400974
rect 493670 400910 493686 400974
rect 493750 400910 493766 400974
rect 493830 400910 493846 400974
rect 493910 400910 493926 400974
rect 493096 400906 493926 400910
rect 493350 400894 493926 400906
rect 494050 400974 494626 400990
rect 494050 400910 494066 400974
rect 494130 400910 494146 400974
rect 494210 400910 494226 400974
rect 494290 400910 494306 400974
rect 494370 400910 494386 400974
rect 494450 400910 494466 400974
rect 494530 400910 494546 400974
rect 494610 400910 494626 400974
rect 494050 400894 494626 400910
rect 493477 400730 493799 400731
rect 494177 400730 494499 400731
rect 494738 400730 494858 401130
rect 493458 400722 494858 400730
rect 493458 400418 493486 400722
rect 493790 400418 494186 400722
rect 494490 400418 494858 400722
rect 493458 400410 494858 400418
rect 493477 400409 493799 400410
rect 494177 400409 494499 400410
rect 493350 400255 493926 400271
rect 493350 400191 493366 400255
rect 493430 400191 493446 400255
rect 493510 400191 493526 400255
rect 493590 400191 493606 400255
rect 493670 400191 493686 400255
rect 493750 400191 493766 400255
rect 493830 400191 493846 400255
rect 493910 400191 493926 400255
rect 493350 400175 493926 400191
rect 494050 400255 494626 400271
rect 494050 400191 494066 400255
rect 494130 400191 494146 400255
rect 494210 400191 494226 400255
rect 494290 400191 494306 400255
rect 494370 400191 494386 400255
rect 494450 400191 494466 400255
rect 494530 400191 494546 400255
rect 494610 400191 494626 400255
rect 494050 400175 494626 400191
rect 493477 400010 493799 400012
rect 494177 400010 494499 400012
rect 494738 400010 494858 400410
rect 493458 400003 494858 400010
rect 493458 399699 493486 400003
rect 493790 399699 494186 400003
rect 494490 399699 494858 400003
rect 493458 399690 494858 399699
rect 493350 399536 493926 399552
rect 493350 399472 493366 399536
rect 493430 399472 493446 399536
rect 493510 399472 493526 399536
rect 493590 399472 493606 399536
rect 493670 399472 493686 399536
rect 493750 399472 493766 399536
rect 493830 399472 493846 399536
rect 493910 399472 493926 399536
rect 493350 399456 493926 399472
rect 494050 399536 494626 399552
rect 494050 399472 494066 399536
rect 494130 399472 494146 399536
rect 494210 399472 494226 399536
rect 494290 399472 494306 399536
rect 494370 399472 494386 399536
rect 494450 399472 494466 399536
rect 494530 399472 494546 399536
rect 494610 399472 494626 399536
rect 494050 399456 494626 399472
rect 493477 399290 493799 399293
rect 494177 399290 494499 399293
rect 494738 399290 494858 399690
rect 502258 399796 502378 399824
rect 502258 399732 502286 399796
rect 502350 399732 502378 399796
rect 502258 399716 502378 399732
rect 502258 399686 502286 399716
rect 500978 399677 502286 399686
rect 500978 399373 501006 399677
rect 501310 399373 501706 399677
rect 502010 399652 502286 399677
rect 502350 399652 502378 399716
rect 502010 399485 502378 399652
rect 502010 399484 502431 399485
rect 502010 399420 502366 399484
rect 502430 399420 502431 399484
rect 502010 399419 502431 399420
rect 502010 399373 502378 399419
rect 500978 399366 502378 399373
rect 500997 399364 501319 399366
rect 501697 399364 502019 399366
rect 493458 399284 494858 399290
rect 493458 398980 493486 399284
rect 493790 398980 494186 399284
rect 494490 398980 494858 399284
rect 500870 399210 501446 399226
rect 500870 399146 500886 399210
rect 500950 399146 500966 399210
rect 501030 399146 501046 399210
rect 501110 399146 501126 399210
rect 501190 399146 501206 399210
rect 501270 399146 501286 399210
rect 501350 399146 501366 399210
rect 501430 399146 501446 399210
rect 500870 399130 501446 399146
rect 501570 399210 502146 399226
rect 501570 399146 501586 399210
rect 501650 399146 501666 399210
rect 501730 399146 501746 399210
rect 501810 399146 501826 399210
rect 501890 399146 501906 399210
rect 501970 399146 501986 399210
rect 502050 399146 502066 399210
rect 502130 399146 502146 399210
rect 501570 399130 502146 399146
rect 493458 398970 494858 398980
rect 493350 398817 493926 398833
rect 493350 398753 493366 398817
rect 493430 398753 493446 398817
rect 493510 398753 493526 398817
rect 493590 398753 493606 398817
rect 493670 398753 493686 398817
rect 493750 398753 493766 398817
rect 493830 398753 493846 398817
rect 493910 398753 493926 398817
rect 493350 398737 493926 398753
rect 494050 398817 494626 398833
rect 494050 398753 494066 398817
rect 494130 398753 494146 398817
rect 494210 398753 494226 398817
rect 494290 398753 494306 398817
rect 494370 398753 494386 398817
rect 494450 398753 494466 398817
rect 494530 398753 494546 398817
rect 494610 398753 494626 398817
rect 494050 398737 494626 398753
rect 493477 398570 493799 398574
rect 494177 398570 494499 398574
rect 494738 398570 494858 398970
rect 500997 398966 501319 398967
rect 501697 398966 502019 398967
rect 502258 398966 502378 399366
rect 500978 398958 502378 398966
rect 500978 398654 501006 398958
rect 501310 398654 501706 398958
rect 502010 398654 502378 398958
rect 500978 398646 502378 398654
rect 500997 398645 501319 398646
rect 501697 398645 502019 398646
rect 493458 398565 494858 398570
rect 493458 398261 493486 398565
rect 493790 398261 494186 398565
rect 494490 398261 494858 398565
rect 500870 398491 501446 398507
rect 500870 398427 500886 398491
rect 500950 398427 500966 398491
rect 501030 398427 501046 398491
rect 501110 398427 501126 398491
rect 501190 398427 501206 398491
rect 501270 398427 501286 398491
rect 501350 398427 501366 398491
rect 501430 398427 501446 398491
rect 500870 398411 501446 398427
rect 501570 398491 502146 398507
rect 501570 398427 501586 398491
rect 501650 398427 501666 398491
rect 501730 398427 501746 398491
rect 501810 398427 501826 398491
rect 501890 398427 501906 398491
rect 501970 398427 501986 398491
rect 502050 398427 502066 398491
rect 502130 398427 502146 398491
rect 501570 398411 502146 398427
rect 493458 398250 494858 398261
rect 493350 398098 493926 398114
rect 493350 398034 493366 398098
rect 493430 398034 493446 398098
rect 493510 398034 493526 398098
rect 493590 398034 493606 398098
rect 493670 398034 493686 398098
rect 493750 398034 493766 398098
rect 493830 398034 493846 398098
rect 493910 398034 493926 398098
rect 493350 398018 493926 398034
rect 494050 398098 494626 398114
rect 494050 398034 494066 398098
rect 494130 398034 494146 398098
rect 494210 398034 494226 398098
rect 494290 398034 494306 398098
rect 494370 398034 494386 398098
rect 494450 398034 494466 398098
rect 494530 398034 494546 398098
rect 494610 398034 494626 398098
rect 494050 398018 494626 398034
rect 493477 397850 493799 397855
rect 494177 397850 494499 397855
rect 494738 397850 494858 398250
rect 500997 398246 501319 398248
rect 501697 398246 502019 398248
rect 502258 398246 502378 398646
rect 500978 398239 502378 398246
rect 500978 397935 501006 398239
rect 501310 397935 501706 398239
rect 502010 397935 502378 398239
rect 500978 397926 502378 397935
rect 493458 397846 494858 397850
rect 493458 397542 493486 397846
rect 493790 397542 494186 397846
rect 494490 397542 494858 397846
rect 500870 397772 501446 397788
rect 500870 397708 500886 397772
rect 500950 397708 500966 397772
rect 501030 397708 501046 397772
rect 501110 397708 501126 397772
rect 501190 397708 501206 397772
rect 501270 397708 501286 397772
rect 501350 397708 501366 397772
rect 501430 397708 501446 397772
rect 500870 397692 501446 397708
rect 501570 397772 502146 397788
rect 501570 397708 501586 397772
rect 501650 397708 501666 397772
rect 501730 397708 501746 397772
rect 501810 397708 501826 397772
rect 501890 397708 501906 397772
rect 501970 397708 501986 397772
rect 502050 397708 502066 397772
rect 502130 397708 502146 397772
rect 501570 397692 502146 397708
rect 493458 397530 494858 397542
rect 493350 397379 493926 397395
rect 493350 397315 493366 397379
rect 493430 397315 493446 397379
rect 493510 397315 493526 397379
rect 493590 397315 493606 397379
rect 493670 397315 493686 397379
rect 493750 397315 493766 397379
rect 493830 397315 493846 397379
rect 493910 397315 493926 397379
rect 493350 397299 493926 397315
rect 494050 397379 494626 397395
rect 494050 397315 494066 397379
rect 494130 397315 494146 397379
rect 494210 397315 494226 397379
rect 494290 397315 494306 397379
rect 494370 397315 494386 397379
rect 494450 397315 494466 397379
rect 494530 397315 494546 397379
rect 494610 397315 494626 397379
rect 494050 397299 494626 397315
rect 494738 397274 494858 397530
rect 500997 397526 501319 397529
rect 501697 397526 502019 397529
rect 502258 397526 502378 397926
rect 500978 397520 502378 397526
rect 494923 397276 494989 397277
rect 494923 397274 494924 397276
rect 494738 397214 494924 397274
rect 493477 397130 493799 397136
rect 494177 397130 494499 397136
rect 494738 397130 494858 397214
rect 494923 397212 494924 397214
rect 494988 397212 494989 397276
rect 494923 397211 494989 397212
rect 500978 397216 501006 397520
rect 501310 397216 501706 397520
rect 502010 397216 502378 397520
rect 500978 397206 502378 397216
rect 493458 397127 494858 397130
rect 493458 396823 493486 397127
rect 493790 396823 494186 397127
rect 494490 396823 494858 397127
rect 500870 397053 501446 397069
rect 500870 396989 500886 397053
rect 500950 396989 500966 397053
rect 501030 396989 501046 397053
rect 501110 396989 501126 397053
rect 501190 396989 501206 397053
rect 501270 396989 501286 397053
rect 501350 396989 501366 397053
rect 501430 396989 501446 397053
rect 500870 396973 501446 396989
rect 501570 397053 502146 397069
rect 501570 396989 501586 397053
rect 501650 396989 501666 397053
rect 501730 396989 501746 397053
rect 501810 396989 501826 397053
rect 501890 396989 501906 397053
rect 501970 396989 501986 397053
rect 502050 396989 502066 397053
rect 502130 396989 502146 397053
rect 501570 396973 502146 396989
rect 493458 396810 494858 396823
rect 493350 396660 493926 396676
rect 493350 396596 493366 396660
rect 493430 396596 493446 396660
rect 493510 396596 493526 396660
rect 493590 396596 493606 396660
rect 493670 396596 493686 396660
rect 493750 396596 493766 396660
rect 493830 396596 493846 396660
rect 493910 396596 493926 396660
rect 493350 396580 493926 396596
rect 494050 396660 494626 396676
rect 494050 396596 494066 396660
rect 494130 396596 494146 396660
rect 494210 396596 494226 396660
rect 494290 396596 494306 396660
rect 494370 396596 494386 396660
rect 494450 396596 494466 396660
rect 494530 396596 494546 396660
rect 494610 396596 494626 396660
rect 494050 396580 494626 396596
rect 493477 396410 493799 396417
rect 494177 396410 494499 396417
rect 494738 396410 494858 396810
rect 500997 396806 501319 396810
rect 501697 396806 502019 396810
rect 502258 396806 502378 397206
rect 500978 396801 502378 396806
rect 500978 396497 501006 396801
rect 501310 396497 501706 396801
rect 502010 396497 502378 396801
rect 500978 396486 502378 396497
rect 493458 396408 494858 396410
rect 493458 396104 493486 396408
rect 493790 396104 494186 396408
rect 494490 396104 494858 396408
rect 500870 396334 501446 396350
rect 500870 396270 500886 396334
rect 500950 396270 500966 396334
rect 501030 396270 501046 396334
rect 501110 396270 501126 396334
rect 501190 396270 501206 396334
rect 501270 396270 501286 396334
rect 501350 396270 501366 396334
rect 501430 396270 501446 396334
rect 500870 396254 501446 396270
rect 501570 396334 502146 396350
rect 501570 396270 501586 396334
rect 501650 396270 501666 396334
rect 501730 396270 501746 396334
rect 501810 396270 501826 396334
rect 501890 396270 501906 396334
rect 501970 396270 501986 396334
rect 502050 396270 502066 396334
rect 502130 396270 502146 396334
rect 501570 396254 502146 396270
rect 493458 396090 494858 396104
rect 493350 395941 493926 395957
rect 493350 395877 493366 395941
rect 493430 395877 493446 395941
rect 493510 395877 493526 395941
rect 493590 395877 493606 395941
rect 493670 395877 493686 395941
rect 493750 395877 493766 395941
rect 493830 395877 493846 395941
rect 493910 395877 493926 395941
rect 493350 395861 493926 395877
rect 494050 395941 494626 395957
rect 494050 395877 494066 395941
rect 494130 395877 494146 395941
rect 494210 395877 494226 395941
rect 494290 395877 494306 395941
rect 494370 395877 494386 395941
rect 494450 395877 494466 395941
rect 494530 395877 494546 395941
rect 494610 395877 494626 395941
rect 494050 395861 494626 395877
rect 493477 395690 493799 395698
rect 494177 395690 494499 395698
rect 494738 395690 494858 396090
rect 500997 396086 501319 396091
rect 501697 396086 502019 396091
rect 502258 396086 502378 396486
rect 500978 396082 502378 396086
rect 500978 395778 501006 396082
rect 501310 395778 501706 396082
rect 502010 395778 502378 396082
rect 500978 395766 502378 395778
rect 493458 395689 494858 395690
rect 493458 395385 493486 395689
rect 493790 395385 494186 395689
rect 494490 395385 494858 395689
rect 500870 395615 501446 395631
rect 500870 395551 500886 395615
rect 500950 395551 500966 395615
rect 501030 395551 501046 395615
rect 501110 395551 501126 395615
rect 501190 395551 501206 395615
rect 501270 395551 501286 395615
rect 501350 395551 501366 395615
rect 501430 395551 501446 395615
rect 500870 395535 501446 395551
rect 501570 395615 502146 395631
rect 501570 395551 501586 395615
rect 501650 395551 501666 395615
rect 501730 395551 501746 395615
rect 501810 395551 501826 395615
rect 501890 395551 501906 395615
rect 501970 395551 501986 395615
rect 502050 395551 502066 395615
rect 502130 395551 502146 395615
rect 501570 395535 502146 395551
rect 493458 395370 494858 395385
rect 493350 395222 493926 395238
rect 493350 395158 493366 395222
rect 493430 395158 493446 395222
rect 493510 395158 493526 395222
rect 493590 395158 493606 395222
rect 493670 395158 493686 395222
rect 493750 395158 493766 395222
rect 493830 395158 493846 395222
rect 493910 395158 493926 395222
rect 493350 395142 493926 395158
rect 494050 395222 494626 395238
rect 494050 395158 494066 395222
rect 494130 395158 494146 395222
rect 494210 395158 494226 395222
rect 494290 395158 494306 395222
rect 494370 395158 494386 395222
rect 494450 395158 494466 395222
rect 494530 395158 494546 395222
rect 494610 395158 494626 395222
rect 494050 395142 494626 395158
rect 493477 394970 493799 394979
rect 494177 394970 494499 394979
rect 494738 394970 494858 395370
rect 500997 395366 501319 395372
rect 501697 395366 502019 395372
rect 502258 395366 502378 395766
rect 500978 395363 502378 395366
rect 500978 395059 501006 395363
rect 501310 395059 501706 395363
rect 502010 395059 502378 395363
rect 500978 395046 502378 395059
rect 493458 394666 493486 394970
rect 493790 394666 494186 394970
rect 494490 394666 494858 394970
rect 500870 394896 501446 394912
rect 500870 394832 500886 394896
rect 500950 394832 500966 394896
rect 501030 394832 501046 394896
rect 501110 394832 501126 394896
rect 501190 394832 501206 394896
rect 501270 394832 501286 394896
rect 501350 394832 501366 394896
rect 501430 394832 501446 394896
rect 500870 394816 501446 394832
rect 501570 394896 502146 394912
rect 501570 394832 501586 394896
rect 501650 394832 501666 394896
rect 501730 394832 501746 394896
rect 501810 394832 501826 394896
rect 501890 394832 501906 394896
rect 501970 394832 501986 394896
rect 502050 394832 502066 394896
rect 502130 394832 502146 394896
rect 501570 394816 502146 394832
rect 493458 394650 494858 394666
rect 493350 394503 493926 394519
rect 493350 394439 493366 394503
rect 493430 394439 493446 394503
rect 493510 394439 493526 394503
rect 493590 394439 493606 394503
rect 493670 394439 493686 394503
rect 493750 394439 493766 394503
rect 493830 394439 493846 394503
rect 493910 394439 493926 394503
rect 493350 394423 493926 394439
rect 494050 394503 494626 394519
rect 494050 394439 494066 394503
rect 494130 394439 494146 394503
rect 494210 394439 494226 394503
rect 494290 394439 494306 394503
rect 494370 394439 494386 394503
rect 494450 394439 494466 394503
rect 494530 394439 494546 394503
rect 494610 394439 494626 394503
rect 494050 394423 494626 394439
rect 494738 394420 494858 394650
rect 500997 394646 501319 394653
rect 501697 394646 502019 394653
rect 502258 394646 502378 395046
rect 500978 394644 502378 394646
rect 500978 394340 501006 394644
rect 501310 394340 501706 394644
rect 502010 394340 502378 394644
rect 500978 394326 502378 394340
rect 500870 394177 501446 394193
rect 500870 394113 500886 394177
rect 500950 394113 500966 394177
rect 501030 394113 501046 394177
rect 501110 394113 501126 394177
rect 501190 394113 501206 394177
rect 501270 394113 501286 394177
rect 501350 394113 501366 394177
rect 501430 394113 501446 394177
rect 500870 394097 501446 394113
rect 501570 394177 502146 394193
rect 501570 394113 501586 394177
rect 501650 394113 501666 394177
rect 501730 394113 501746 394177
rect 501810 394113 501826 394177
rect 501890 394113 501906 394177
rect 501970 394113 501986 394177
rect 502050 394113 502066 394177
rect 502130 394113 502146 394177
rect 501570 394097 502146 394113
rect 500997 393926 501319 393934
rect 501697 393926 502019 393934
rect 502258 393926 502378 394326
rect 500978 393925 502378 393926
rect 500978 393621 501006 393925
rect 501310 393621 501706 393925
rect 502010 393621 502378 393925
rect 500978 393606 502378 393621
rect 500870 393458 501446 393474
rect 500870 393394 500886 393458
rect 500950 393394 500966 393458
rect 501030 393394 501046 393458
rect 501110 393394 501126 393458
rect 501190 393394 501206 393458
rect 501270 393394 501286 393458
rect 501350 393394 501366 393458
rect 501430 393394 501446 393458
rect 500870 393378 501446 393394
rect 501570 393458 502146 393474
rect 501570 393394 501586 393458
rect 501650 393394 501666 393458
rect 501730 393394 501746 393458
rect 501810 393394 501826 393458
rect 501890 393394 501906 393458
rect 501970 393394 501986 393458
rect 502050 393394 502066 393458
rect 502130 393394 502146 393458
rect 501570 393378 502146 393394
rect 500997 393206 501319 393215
rect 501697 393206 502019 393215
rect 502258 393206 502378 393606
rect 500978 392902 501006 393206
rect 501310 392902 501706 393206
rect 502010 392902 502378 393206
rect 500978 392886 502378 392902
rect 500870 392739 501446 392755
rect 500657 392722 500723 392723
rect 500657 392658 500658 392722
rect 500722 392720 500723 392722
rect 500870 392720 500886 392739
rect 500722 392675 500886 392720
rect 500950 392675 500966 392739
rect 501030 392675 501046 392739
rect 501110 392675 501126 392739
rect 501190 392675 501206 392739
rect 501270 392675 501286 392739
rect 501350 392675 501366 392739
rect 501430 392675 501446 392739
rect 500722 392660 501446 392675
rect 500722 392658 500723 392660
rect 500870 392659 501446 392660
rect 501570 392739 502146 392755
rect 501570 392675 501586 392739
rect 501650 392675 501666 392739
rect 501730 392675 501746 392739
rect 501810 392675 501826 392739
rect 501890 392675 501906 392739
rect 501970 392675 501986 392739
rect 502050 392675 502066 392739
rect 502130 392675 502146 392739
rect 501570 392659 502146 392675
rect 500657 392657 500723 392658
rect 502258 392656 502378 392886
rect 509778 388722 509898 388750
rect 509778 388658 509806 388722
rect 509870 388658 509898 388722
rect 509778 388642 509898 388658
rect 509778 388612 509806 388642
rect 508498 388603 509806 388612
rect 508498 388299 508526 388603
rect 508830 388299 509226 388603
rect 509530 388578 509806 388603
rect 509870 388578 509898 388642
rect 509530 388299 509898 388578
rect 508498 388292 509898 388299
rect 508517 388290 508839 388292
rect 509217 388290 509539 388292
rect 508390 388136 508966 388152
rect 508390 388072 508406 388136
rect 508470 388072 508486 388136
rect 508550 388072 508566 388136
rect 508630 388072 508646 388136
rect 508710 388072 508726 388136
rect 508790 388072 508806 388136
rect 508870 388072 508886 388136
rect 508950 388072 508966 388136
rect 508390 388056 508966 388072
rect 509090 388136 509666 388152
rect 509090 388072 509106 388136
rect 509170 388072 509186 388136
rect 509250 388072 509266 388136
rect 509330 388072 509346 388136
rect 509410 388072 509426 388136
rect 509490 388072 509506 388136
rect 509570 388072 509586 388136
rect 509650 388072 509666 388136
rect 509090 388056 509666 388072
rect 508517 387892 508839 387893
rect 509217 387892 509539 387893
rect 509778 387892 509898 388292
rect 508498 387884 509898 387892
rect 508498 387580 508526 387884
rect 508830 387580 509226 387884
rect 509530 387580 509898 387884
rect 508498 387572 509898 387580
rect 508517 387571 508839 387572
rect 509217 387571 509539 387572
rect 508390 387417 508966 387433
rect 508390 387353 508406 387417
rect 508470 387353 508486 387417
rect 508550 387353 508566 387417
rect 508630 387353 508646 387417
rect 508710 387353 508726 387417
rect 508790 387353 508806 387417
rect 508870 387353 508886 387417
rect 508950 387353 508966 387417
rect 508390 387337 508966 387353
rect 509090 387417 509666 387433
rect 509090 387353 509106 387417
rect 509170 387353 509186 387417
rect 509250 387353 509266 387417
rect 509330 387353 509346 387417
rect 509410 387353 509426 387417
rect 509490 387353 509506 387417
rect 509570 387353 509586 387417
rect 509650 387353 509666 387417
rect 509090 387337 509666 387353
rect 508517 387172 508839 387174
rect 509217 387172 509539 387174
rect 509778 387172 509898 387572
rect 508498 387165 509898 387172
rect 508498 386861 508526 387165
rect 508830 386861 509226 387165
rect 509530 386861 509898 387165
rect 508498 386852 509898 386861
rect 508390 386698 508966 386714
rect 508390 386634 508406 386698
rect 508470 386634 508486 386698
rect 508550 386634 508566 386698
rect 508630 386634 508646 386698
rect 508710 386634 508726 386698
rect 508790 386634 508806 386698
rect 508870 386634 508886 386698
rect 508950 386634 508966 386698
rect 508390 386618 508966 386634
rect 509090 386698 509666 386714
rect 509090 386634 509106 386698
rect 509170 386634 509186 386698
rect 509250 386634 509266 386698
rect 509330 386634 509346 386698
rect 509410 386634 509426 386698
rect 509490 386634 509506 386698
rect 509570 386634 509586 386698
rect 509650 386634 509666 386698
rect 509090 386618 509666 386634
rect 508517 386452 508839 386455
rect 509217 386452 509539 386455
rect 509778 386452 509898 386852
rect 508498 386446 509898 386452
rect 508498 386142 508526 386446
rect 508830 386142 509226 386446
rect 509530 386142 509898 386446
rect 508498 386132 509898 386142
rect 508390 385979 508966 385995
rect 508390 385915 508406 385979
rect 508470 385915 508486 385979
rect 508550 385915 508566 385979
rect 508630 385915 508646 385979
rect 508710 385915 508726 385979
rect 508790 385915 508806 385979
rect 508870 385915 508886 385979
rect 508950 385915 508966 385979
rect 508390 385899 508966 385915
rect 509090 385979 509666 385995
rect 509090 385915 509106 385979
rect 509170 385915 509186 385979
rect 509250 385915 509266 385979
rect 509330 385915 509346 385979
rect 509410 385915 509426 385979
rect 509490 385915 509506 385979
rect 509570 385915 509586 385979
rect 509650 385915 509666 385979
rect 509090 385899 509666 385915
rect 508517 385732 508839 385736
rect 509217 385732 509539 385736
rect 509778 385732 509898 386132
rect 508498 385727 509898 385732
rect 508498 385423 508526 385727
rect 508830 385423 509226 385727
rect 509530 385423 509898 385727
rect 508498 385412 509898 385423
rect 505049 385270 505115 385271
rect 505049 385206 505050 385270
rect 505114 385206 505115 385270
rect 505049 385205 505115 385206
rect 508390 385260 508966 385276
rect 505052 384888 505112 385205
rect 508390 385196 508406 385260
rect 508470 385196 508486 385260
rect 508550 385196 508566 385260
rect 508630 385196 508646 385260
rect 508710 385196 508726 385260
rect 508790 385196 508806 385260
rect 508870 385196 508886 385260
rect 508950 385196 508966 385260
rect 508390 385180 508966 385196
rect 509090 385260 509666 385276
rect 509090 385196 509106 385260
rect 509170 385196 509186 385260
rect 509250 385196 509266 385260
rect 509330 385196 509346 385260
rect 509410 385196 509426 385260
rect 509490 385196 509506 385260
rect 509570 385196 509586 385260
rect 509650 385196 509666 385260
rect 509090 385180 509666 385196
rect 506018 384998 506138 385026
rect 508517 385012 508839 385017
rect 509217 385012 509539 385017
rect 509778 385012 509898 385412
rect 516273 385270 516339 385271
rect 516273 385206 516274 385270
rect 516338 385206 516339 385270
rect 516273 385205 516339 385206
rect 506018 384934 506046 384998
rect 506110 384934 506138 384998
rect 506018 384918 506138 384934
rect 506018 384888 506046 384918
rect 504738 384879 506046 384888
rect 504738 384575 504766 384879
rect 505070 384575 505466 384879
rect 505770 384854 506046 384879
rect 506110 384854 506138 384918
rect 505770 384575 506138 384854
rect 508498 385008 509898 385012
rect 508498 384704 508526 385008
rect 508830 384704 509226 385008
rect 509530 384704 509898 385008
rect 513538 384998 513658 385026
rect 513538 384934 513566 384998
rect 513630 384934 513658 384998
rect 513538 384918 513658 384934
rect 513538 384888 513566 384918
rect 508498 384692 509898 384704
rect 504738 384568 506138 384575
rect 504757 384566 505079 384568
rect 505457 384566 505779 384568
rect 504630 384412 505206 384428
rect 504630 384348 504646 384412
rect 504710 384348 504726 384412
rect 504790 384348 504806 384412
rect 504870 384348 504886 384412
rect 504950 384348 504966 384412
rect 505030 384348 505046 384412
rect 505110 384348 505126 384412
rect 505190 384348 505206 384412
rect 504630 384332 505206 384348
rect 505330 384412 505906 384428
rect 505330 384348 505346 384412
rect 505410 384348 505426 384412
rect 505490 384348 505506 384412
rect 505570 384348 505586 384412
rect 505650 384348 505666 384412
rect 505730 384348 505746 384412
rect 505810 384348 505826 384412
rect 505890 384348 505906 384412
rect 505330 384332 505906 384348
rect 504757 384168 505079 384169
rect 505457 384168 505779 384169
rect 506018 384168 506138 384568
rect 508390 384541 508966 384557
rect 508390 384477 508406 384541
rect 508470 384477 508486 384541
rect 508550 384477 508566 384541
rect 508630 384477 508646 384541
rect 508710 384477 508726 384541
rect 508790 384477 508806 384541
rect 508870 384477 508886 384541
rect 508950 384477 508966 384541
rect 508390 384461 508966 384477
rect 509090 384541 509666 384557
rect 509090 384477 509106 384541
rect 509170 384477 509186 384541
rect 509250 384477 509266 384541
rect 509330 384477 509346 384541
rect 509410 384477 509426 384541
rect 509490 384477 509506 384541
rect 509570 384477 509586 384541
rect 509650 384477 509666 384541
rect 509090 384461 509666 384477
rect 508517 384292 508839 384298
rect 509217 384292 509539 384298
rect 509778 384292 509898 384692
rect 512258 384879 513566 384888
rect 512258 384575 512286 384879
rect 512590 384575 512986 384879
rect 513290 384854 513566 384879
rect 513630 384854 513658 384918
rect 516276 384888 516336 385205
rect 517298 384998 517418 385026
rect 517298 384934 517326 384998
rect 517390 384934 517418 384998
rect 517298 384918 517418 384934
rect 517298 384888 517326 384918
rect 513290 384575 513658 384854
rect 512258 384568 513658 384575
rect 516018 384879 517326 384888
rect 516018 384575 516046 384879
rect 516350 384575 516746 384879
rect 517050 384854 517326 384879
rect 517390 384854 517418 384918
rect 517050 384575 517418 384854
rect 516018 384568 517418 384575
rect 512277 384566 512599 384568
rect 512977 384566 513299 384568
rect 512150 384412 512726 384428
rect 512150 384348 512166 384412
rect 512230 384348 512246 384412
rect 512310 384348 512326 384412
rect 512390 384348 512406 384412
rect 512470 384348 512486 384412
rect 512550 384348 512566 384412
rect 512630 384348 512646 384412
rect 512710 384348 512726 384412
rect 512150 384332 512726 384348
rect 512850 384412 513426 384428
rect 512850 384348 512866 384412
rect 512930 384348 512946 384412
rect 513010 384348 513026 384412
rect 513090 384348 513106 384412
rect 513170 384348 513186 384412
rect 513250 384348 513266 384412
rect 513330 384348 513346 384412
rect 513410 384348 513426 384412
rect 512850 384332 513426 384348
rect 504738 384160 506138 384168
rect 504738 383856 504766 384160
rect 505070 383856 505466 384160
rect 505770 383856 506138 384160
rect 508498 384289 509898 384292
rect 508498 383985 508526 384289
rect 508830 383985 509226 384289
rect 509530 383985 509898 384289
rect 512277 384168 512599 384169
rect 512977 384168 513299 384169
rect 513538 384168 513658 384568
rect 516037 384566 516359 384568
rect 516737 384566 517059 384568
rect 515910 384412 516486 384428
rect 515910 384348 515926 384412
rect 515990 384348 516006 384412
rect 516070 384348 516086 384412
rect 516150 384348 516166 384412
rect 516230 384348 516246 384412
rect 516310 384348 516326 384412
rect 516390 384348 516406 384412
rect 516470 384348 516486 384412
rect 515910 384332 516486 384348
rect 516610 384412 517186 384428
rect 516610 384348 516626 384412
rect 516690 384348 516706 384412
rect 516770 384348 516786 384412
rect 516850 384348 516866 384412
rect 516930 384348 516946 384412
rect 517010 384348 517026 384412
rect 517090 384348 517106 384412
rect 517170 384348 517186 384412
rect 516610 384332 517186 384348
rect 516037 384168 516359 384169
rect 516737 384168 517059 384169
rect 517298 384168 517418 384568
rect 508498 383972 509898 383985
rect 504738 383848 506138 383856
rect 504757 383847 505079 383848
rect 505457 383847 505779 383848
rect 504630 383693 505206 383709
rect 504630 383629 504646 383693
rect 504710 383629 504726 383693
rect 504790 383629 504806 383693
rect 504870 383629 504886 383693
rect 504950 383629 504966 383693
rect 505030 383629 505046 383693
rect 505110 383629 505126 383693
rect 505190 383629 505206 383693
rect 504630 383613 505206 383629
rect 505330 383693 505906 383709
rect 505330 383629 505346 383693
rect 505410 383629 505426 383693
rect 505490 383629 505506 383693
rect 505570 383629 505586 383693
rect 505650 383629 505666 383693
rect 505730 383629 505746 383693
rect 505810 383629 505826 383693
rect 505890 383629 505906 383693
rect 505330 383613 505906 383629
rect 504757 383448 505079 383450
rect 505457 383448 505779 383450
rect 506018 383448 506138 383848
rect 508390 383822 508966 383838
rect 508390 383758 508406 383822
rect 508470 383758 508486 383822
rect 508550 383758 508566 383822
rect 508630 383758 508646 383822
rect 508710 383758 508726 383822
rect 508790 383758 508806 383822
rect 508870 383758 508886 383822
rect 508950 383758 508966 383822
rect 508390 383742 508966 383758
rect 509090 383822 509666 383838
rect 509090 383758 509106 383822
rect 509170 383758 509186 383822
rect 509250 383758 509266 383822
rect 509330 383758 509346 383822
rect 509410 383758 509426 383822
rect 509490 383758 509506 383822
rect 509570 383758 509586 383822
rect 509650 383758 509666 383822
rect 509090 383742 509666 383758
rect 508517 383572 508839 383579
rect 509217 383572 509539 383579
rect 509778 383572 509898 383972
rect 512258 384160 513658 384168
rect 512258 383856 512286 384160
rect 512590 383856 512986 384160
rect 513290 383856 513658 384160
rect 512258 383848 513658 383856
rect 516018 384160 517418 384168
rect 516018 383856 516046 384160
rect 516350 383856 516746 384160
rect 517050 383856 517418 384160
rect 516018 383848 517418 383856
rect 512277 383847 512599 383848
rect 512977 383847 513299 383848
rect 512150 383693 512726 383709
rect 512150 383629 512166 383693
rect 512230 383629 512246 383693
rect 512310 383629 512326 383693
rect 512390 383629 512406 383693
rect 512470 383629 512486 383693
rect 512550 383629 512566 383693
rect 512630 383629 512646 383693
rect 512710 383629 512726 383693
rect 512150 383613 512726 383629
rect 512850 383693 513426 383709
rect 512850 383629 512866 383693
rect 512930 383629 512946 383693
rect 513010 383629 513026 383693
rect 513090 383629 513106 383693
rect 513170 383629 513186 383693
rect 513250 383629 513266 383693
rect 513330 383629 513346 383693
rect 513410 383629 513426 383693
rect 512850 383613 513426 383629
rect 504738 383441 506138 383448
rect 504738 383137 504766 383441
rect 505070 383137 505466 383441
rect 505770 383137 506138 383441
rect 508498 383570 509898 383572
rect 508498 383266 508526 383570
rect 508830 383266 509226 383570
rect 509530 383266 509898 383570
rect 512277 383448 512599 383450
rect 512977 383448 513299 383450
rect 513538 383448 513658 383848
rect 516037 383847 516359 383848
rect 516737 383847 517059 383848
rect 515910 383693 516486 383709
rect 515910 383629 515926 383693
rect 515990 383629 516006 383693
rect 516070 383629 516086 383693
rect 516150 383629 516166 383693
rect 516230 383629 516246 383693
rect 516310 383629 516326 383693
rect 516390 383629 516406 383693
rect 516470 383629 516486 383693
rect 515910 383613 516486 383629
rect 516610 383693 517186 383709
rect 516610 383629 516626 383693
rect 516690 383629 516706 383693
rect 516770 383629 516786 383693
rect 516850 383629 516866 383693
rect 516930 383629 516946 383693
rect 517010 383629 517026 383693
rect 517090 383629 517106 383693
rect 517170 383629 517186 383693
rect 516610 383613 517186 383629
rect 516037 383448 516359 383450
rect 516737 383448 517059 383450
rect 517298 383448 517418 383848
rect 508498 383252 509898 383266
rect 504738 383128 506138 383137
rect 504630 382974 505206 382990
rect 504630 382910 504646 382974
rect 504710 382910 504726 382974
rect 504790 382910 504806 382974
rect 504870 382910 504886 382974
rect 504950 382910 504966 382974
rect 505030 382910 505046 382974
rect 505110 382910 505126 382974
rect 505190 382910 505206 382974
rect 504630 382894 505206 382910
rect 505330 382974 505906 382990
rect 505330 382910 505346 382974
rect 505410 382910 505426 382974
rect 505490 382910 505506 382974
rect 505570 382910 505586 382974
rect 505650 382910 505666 382974
rect 505730 382910 505746 382974
rect 505810 382910 505826 382974
rect 505890 382910 505906 382974
rect 505330 382894 505906 382910
rect 504757 382728 505079 382731
rect 505457 382728 505779 382731
rect 506018 382728 506138 383128
rect 508390 383103 508966 383119
rect 508390 383039 508406 383103
rect 508470 383039 508486 383103
rect 508550 383039 508566 383103
rect 508630 383039 508646 383103
rect 508710 383039 508726 383103
rect 508790 383039 508806 383103
rect 508870 383039 508886 383103
rect 508950 383039 508966 383103
rect 508390 383023 508966 383039
rect 509090 383103 509666 383119
rect 509090 383039 509106 383103
rect 509170 383039 509186 383103
rect 509250 383039 509266 383103
rect 509330 383039 509346 383103
rect 509410 383039 509426 383103
rect 509490 383039 509506 383103
rect 509570 383039 509586 383103
rect 509650 383039 509666 383103
rect 509090 383023 509666 383039
rect 508517 382852 508839 382860
rect 509217 382852 509539 382860
rect 509778 382852 509898 383252
rect 512258 383441 513658 383448
rect 512258 383137 512286 383441
rect 512590 383137 512986 383441
rect 513290 383336 513658 383441
rect 516018 383441 517418 383448
rect 516018 383336 516046 383441
rect 513290 383276 516046 383336
rect 513290 383137 513658 383276
rect 512258 383128 513658 383137
rect 516018 383137 516046 383276
rect 516350 383137 516746 383441
rect 517050 383137 517418 383441
rect 516018 383128 517418 383137
rect 512150 382974 512726 382990
rect 512150 382910 512166 382974
rect 512230 382910 512246 382974
rect 512310 382910 512326 382974
rect 512390 382910 512406 382974
rect 512470 382910 512486 382974
rect 512550 382910 512566 382974
rect 512630 382910 512646 382974
rect 512710 382910 512726 382974
rect 512150 382894 512726 382910
rect 512850 382974 513426 382990
rect 512850 382910 512866 382974
rect 512930 382910 512946 382974
rect 513010 382910 513026 382974
rect 513090 382910 513106 382974
rect 513170 382910 513186 382974
rect 513250 382910 513266 382974
rect 513330 382910 513346 382974
rect 513410 382910 513426 382974
rect 512850 382894 513426 382910
rect 504738 382722 506138 382728
rect 504738 382418 504766 382722
rect 505070 382418 505466 382722
rect 505770 382418 506138 382722
rect 508498 382851 509898 382852
rect 508498 382547 508526 382851
rect 508830 382547 509226 382851
rect 509530 382547 509898 382851
rect 512277 382728 512599 382731
rect 512977 382728 513299 382731
rect 513538 382728 513658 383128
rect 515910 382974 516486 382990
rect 515910 382910 515926 382974
rect 515990 382910 516006 382974
rect 516070 382910 516086 382974
rect 516150 382910 516166 382974
rect 516230 382910 516246 382974
rect 516310 382910 516326 382974
rect 516390 382910 516406 382974
rect 516470 382910 516486 382974
rect 515910 382894 516486 382910
rect 516610 382974 517186 382990
rect 516610 382910 516626 382974
rect 516690 382910 516706 382974
rect 516770 382910 516786 382974
rect 516850 382910 516866 382974
rect 516930 382910 516946 382974
rect 517010 382910 517026 382974
rect 517090 382910 517106 382974
rect 517170 382910 517186 382974
rect 516610 382894 517186 382910
rect 516037 382728 516359 382731
rect 516737 382728 517059 382731
rect 517298 382728 517418 383128
rect 508498 382532 509898 382547
rect 504738 382408 506138 382418
rect 504630 382255 505206 382271
rect 504630 382191 504646 382255
rect 504710 382191 504726 382255
rect 504790 382191 504806 382255
rect 504870 382191 504886 382255
rect 504950 382191 504966 382255
rect 505030 382191 505046 382255
rect 505110 382191 505126 382255
rect 505190 382191 505206 382255
rect 504630 382175 505206 382191
rect 505330 382255 505906 382271
rect 505330 382191 505346 382255
rect 505410 382191 505426 382255
rect 505490 382191 505506 382255
rect 505570 382191 505586 382255
rect 505650 382191 505666 382255
rect 505730 382191 505746 382255
rect 505810 382191 505826 382255
rect 505890 382191 505906 382255
rect 505330 382175 505906 382191
rect 504757 382008 505079 382012
rect 505457 382008 505779 382012
rect 506018 382008 506138 382408
rect 508390 382384 508966 382400
rect 508390 382320 508406 382384
rect 508470 382320 508486 382384
rect 508550 382320 508566 382384
rect 508630 382320 508646 382384
rect 508710 382320 508726 382384
rect 508790 382320 508806 382384
rect 508870 382320 508886 382384
rect 508950 382320 508966 382384
rect 508390 382304 508966 382320
rect 509090 382384 509666 382400
rect 509090 382320 509106 382384
rect 509170 382320 509186 382384
rect 509250 382320 509266 382384
rect 509330 382320 509346 382384
rect 509410 382320 509426 382384
rect 509490 382320 509506 382384
rect 509570 382320 509586 382384
rect 509650 382320 509666 382384
rect 509090 382304 509666 382320
rect 508517 382132 508839 382141
rect 509217 382132 509539 382141
rect 509778 382132 509898 382532
rect 512258 382722 513658 382728
rect 512258 382418 512286 382722
rect 512590 382418 512986 382722
rect 513290 382418 513658 382722
rect 512258 382408 513658 382418
rect 516018 382722 517418 382728
rect 516018 382418 516046 382722
rect 516350 382418 516746 382722
rect 517050 382418 517418 382722
rect 516018 382408 517418 382418
rect 512150 382255 512726 382271
rect 512150 382191 512166 382255
rect 512230 382191 512246 382255
rect 512310 382191 512326 382255
rect 512390 382191 512406 382255
rect 512470 382191 512486 382255
rect 512550 382191 512566 382255
rect 512630 382191 512646 382255
rect 512710 382191 512726 382255
rect 512150 382175 512726 382191
rect 512850 382255 513426 382271
rect 512850 382191 512866 382255
rect 512930 382191 512946 382255
rect 513010 382191 513026 382255
rect 513090 382191 513106 382255
rect 513170 382191 513186 382255
rect 513250 382191 513266 382255
rect 513330 382191 513346 382255
rect 513410 382191 513426 382255
rect 512850 382175 513426 382191
rect 504738 382003 506138 382008
rect 504738 381699 504766 382003
rect 505070 381699 505466 382003
rect 505770 381956 506138 382003
rect 508498 381956 508526 382132
rect 505770 381896 508526 381956
rect 505770 381699 506138 381896
rect 508498 381828 508526 381896
rect 508830 381828 509226 382132
rect 509530 381828 509898 382132
rect 512277 382008 512599 382012
rect 512977 382008 513299 382012
rect 513538 382008 513658 382408
rect 515910 382255 516486 382271
rect 515910 382191 515926 382255
rect 515990 382191 516006 382255
rect 516070 382191 516086 382255
rect 516150 382191 516166 382255
rect 516230 382191 516246 382255
rect 516310 382191 516326 382255
rect 516390 382191 516406 382255
rect 516470 382191 516486 382255
rect 515910 382175 516486 382191
rect 516610 382255 517186 382271
rect 516610 382191 516626 382255
rect 516690 382191 516706 382255
rect 516770 382191 516786 382255
rect 516850 382191 516866 382255
rect 516930 382191 516946 382255
rect 517010 382191 517026 382255
rect 517090 382191 517106 382255
rect 517170 382191 517186 382255
rect 516610 382175 517186 382191
rect 516037 382008 516359 382012
rect 516737 382008 517059 382012
rect 517298 382008 517418 382408
rect 508498 381812 509898 381828
rect 504738 381688 506138 381699
rect 504439 381544 504505 381545
rect 504439 381480 504440 381544
rect 504504 381542 504505 381544
rect 504630 381542 505206 381552
rect 504504 381536 505206 381542
rect 504504 381482 504646 381536
rect 504504 381480 504505 381482
rect 504439 381479 504505 381480
rect 504630 381472 504646 381482
rect 504710 381472 504726 381536
rect 504790 381472 504806 381536
rect 504870 381472 504886 381536
rect 504950 381472 504966 381536
rect 505030 381472 505046 381536
rect 505110 381472 505126 381536
rect 505190 381472 505206 381536
rect 504630 381456 505206 381472
rect 505330 381536 505906 381552
rect 505330 381472 505346 381536
rect 505410 381472 505426 381536
rect 505490 381472 505506 381536
rect 505570 381472 505586 381536
rect 505650 381472 505666 381536
rect 505730 381472 505746 381536
rect 505810 381472 505826 381536
rect 505890 381472 505906 381536
rect 505330 381456 505906 381472
rect 504757 381288 505079 381293
rect 505457 381288 505779 381293
rect 506018 381288 506138 381688
rect 508221 381682 508287 381683
rect 508221 381618 508222 381682
rect 508286 381680 508287 381682
rect 508390 381680 508966 381681
rect 508286 381665 508966 381680
rect 508286 381620 508406 381665
rect 508286 381618 508287 381620
rect 508221 381617 508287 381618
rect 508390 381601 508406 381620
rect 508470 381601 508486 381665
rect 508550 381601 508566 381665
rect 508630 381601 508646 381665
rect 508710 381601 508726 381665
rect 508790 381601 508806 381665
rect 508870 381601 508886 381665
rect 508950 381601 508966 381665
rect 508390 381585 508966 381601
rect 509090 381665 509666 381681
rect 509090 381601 509106 381665
rect 509170 381601 509186 381665
rect 509250 381601 509266 381665
rect 509330 381601 509346 381665
rect 509410 381601 509426 381665
rect 509490 381601 509506 381665
rect 509570 381601 509586 381665
rect 509650 381601 509666 381665
rect 509090 381585 509666 381601
rect 509778 381582 509898 381812
rect 512258 382003 513658 382008
rect 512258 381699 512286 382003
rect 512590 381699 512986 382003
rect 513290 381699 513658 382003
rect 512258 381688 513658 381699
rect 516018 382003 517418 382008
rect 516018 381699 516046 382003
rect 516350 381699 516746 382003
rect 517050 381699 517418 382003
rect 516018 381688 517418 381699
rect 509810 381302 509870 381582
rect 511881 381544 511947 381545
rect 511881 381480 511882 381544
rect 511946 381542 511947 381544
rect 512150 381542 512726 381552
rect 511946 381536 512726 381542
rect 511946 381482 512166 381536
rect 511946 381480 511947 381482
rect 511881 381479 511947 381480
rect 512150 381472 512166 381482
rect 512230 381472 512246 381536
rect 512310 381472 512326 381536
rect 512390 381472 512406 381536
rect 512470 381472 512486 381536
rect 512550 381472 512566 381536
rect 512630 381472 512646 381536
rect 512710 381472 512726 381536
rect 512150 381456 512726 381472
rect 512850 381536 513426 381552
rect 512850 381472 512866 381536
rect 512930 381472 512946 381536
rect 513010 381472 513026 381536
rect 513090 381472 513106 381536
rect 513170 381472 513186 381536
rect 513250 381472 513266 381536
rect 513330 381472 513346 381536
rect 513410 381472 513426 381536
rect 512850 381456 513426 381472
rect 504738 381284 506138 381288
rect 504738 380980 504766 381284
rect 505070 380980 505466 381284
rect 505770 380980 506138 381284
rect 509778 381274 509898 381302
rect 512277 381288 512599 381293
rect 512977 381288 513299 381293
rect 513538 381288 513658 381688
rect 515663 381544 515729 381545
rect 515663 381480 515664 381544
rect 515728 381542 515729 381544
rect 515910 381542 516486 381552
rect 515728 381536 516486 381542
rect 515728 381482 515926 381536
rect 515728 381480 515729 381482
rect 515663 381479 515729 381480
rect 515910 381472 515926 381482
rect 515990 381472 516006 381536
rect 516070 381472 516086 381536
rect 516150 381472 516166 381536
rect 516230 381472 516246 381536
rect 516310 381472 516326 381536
rect 516390 381472 516406 381536
rect 516470 381472 516486 381536
rect 515910 381456 516486 381472
rect 516610 381536 517186 381552
rect 516610 381472 516626 381536
rect 516690 381472 516706 381536
rect 516770 381472 516786 381536
rect 516850 381472 516866 381536
rect 516930 381472 516946 381536
rect 517010 381472 517026 381536
rect 517090 381472 517106 381536
rect 517170 381472 517186 381536
rect 516610 381456 517186 381472
rect 516037 381288 516359 381293
rect 516737 381288 517059 381293
rect 517298 381288 517418 381688
rect 509778 381210 509806 381274
rect 509870 381210 509898 381274
rect 509778 381194 509898 381210
rect 509778 381164 509806 381194
rect 504738 380968 506138 380980
rect 504630 380817 505206 380833
rect 504630 380753 504646 380817
rect 504710 380753 504726 380817
rect 504790 380753 504806 380817
rect 504870 380753 504886 380817
rect 504950 380753 504966 380817
rect 505030 380753 505046 380817
rect 505110 380753 505126 380817
rect 505190 380753 505206 380817
rect 504630 380737 505206 380753
rect 505330 380817 505906 380833
rect 505330 380753 505346 380817
rect 505410 380753 505426 380817
rect 505490 380753 505506 380817
rect 505570 380753 505586 380817
rect 505650 380753 505666 380817
rect 505730 380753 505746 380817
rect 505810 380753 505826 380817
rect 505890 380753 505906 380817
rect 505330 380737 505906 380753
rect 504757 380568 505079 380574
rect 505457 380568 505779 380574
rect 506018 380568 506138 380968
rect 508498 381155 509806 381164
rect 508221 380854 508287 380855
rect 508221 380790 508222 380854
rect 508286 380790 508287 380854
rect 508498 380851 508526 381155
rect 508830 380851 509226 381155
rect 509530 381130 509806 381155
rect 509870 381130 509898 381194
rect 509530 381128 509898 381130
rect 512258 381284 513658 381288
rect 512258 381128 512286 381284
rect 509530 381068 512286 381128
rect 509530 380851 509898 381068
rect 512258 380980 512286 381068
rect 512590 380980 512986 381284
rect 513290 380980 513658 381284
rect 512258 380968 513658 380980
rect 516018 381284 517418 381288
rect 516018 380980 516046 381284
rect 516350 380980 516746 381284
rect 517050 380980 517418 381284
rect 516018 380968 517418 380980
rect 508498 380844 509898 380851
rect 508517 380842 508839 380844
rect 509217 380842 509539 380844
rect 508221 380789 508287 380790
rect 508224 380680 508284 380789
rect 508390 380688 508966 380704
rect 508390 380680 508406 380688
rect 508224 380624 508406 380680
rect 508470 380624 508486 380688
rect 508550 380624 508566 380688
rect 508630 380624 508646 380688
rect 508710 380624 508726 380688
rect 508790 380624 508806 380688
rect 508870 380624 508886 380688
rect 508950 380624 508966 380688
rect 508224 380620 508966 380624
rect 508390 380608 508966 380620
rect 509090 380688 509666 380704
rect 509090 380624 509106 380688
rect 509170 380624 509186 380688
rect 509250 380624 509266 380688
rect 509330 380624 509346 380688
rect 509410 380624 509426 380688
rect 509490 380624 509506 380688
rect 509570 380624 509586 380688
rect 509650 380624 509666 380688
rect 509090 380608 509666 380624
rect 504738 380565 506138 380568
rect 504738 380261 504766 380565
rect 505070 380261 505466 380565
rect 505770 380261 506138 380565
rect 508517 380444 508839 380445
rect 509217 380444 509539 380445
rect 509778 380444 509898 380844
rect 512150 380817 512726 380833
rect 512150 380753 512166 380817
rect 512230 380753 512246 380817
rect 512310 380753 512326 380817
rect 512390 380753 512406 380817
rect 512470 380753 512486 380817
rect 512550 380753 512566 380817
rect 512630 380753 512646 380817
rect 512710 380753 512726 380817
rect 512150 380737 512726 380753
rect 512850 380817 513426 380833
rect 512850 380753 512866 380817
rect 512930 380753 512946 380817
rect 513010 380753 513026 380817
rect 513090 380753 513106 380817
rect 513170 380753 513186 380817
rect 513250 380753 513266 380817
rect 513330 380753 513346 380817
rect 513410 380753 513426 380817
rect 512850 380737 513426 380753
rect 512277 380568 512599 380574
rect 512977 380568 513299 380574
rect 513538 380568 513658 380968
rect 515910 380817 516486 380833
rect 515910 380753 515926 380817
rect 515990 380753 516006 380817
rect 516070 380753 516086 380817
rect 516150 380753 516166 380817
rect 516230 380753 516246 380817
rect 516310 380753 516326 380817
rect 516390 380753 516406 380817
rect 516470 380753 516486 380817
rect 515910 380737 516486 380753
rect 516610 380817 517186 380833
rect 516610 380753 516626 380817
rect 516690 380753 516706 380817
rect 516770 380753 516786 380817
rect 516850 380753 516866 380817
rect 516930 380753 516946 380817
rect 517010 380753 517026 380817
rect 517090 380753 517106 380817
rect 517170 380753 517186 380817
rect 516610 380737 517186 380753
rect 516037 380568 516359 380574
rect 516737 380568 517059 380574
rect 517298 380568 517418 380968
rect 504738 380248 506138 380261
rect 504630 380098 505206 380114
rect 504630 380034 504646 380098
rect 504710 380034 504726 380098
rect 504790 380034 504806 380098
rect 504870 380034 504886 380098
rect 504950 380034 504966 380098
rect 505030 380034 505046 380098
rect 505110 380034 505126 380098
rect 505190 380034 505206 380098
rect 504630 380018 505206 380034
rect 505330 380098 505906 380114
rect 505330 380034 505346 380098
rect 505410 380034 505426 380098
rect 505490 380034 505506 380098
rect 505570 380034 505586 380098
rect 505650 380034 505666 380098
rect 505730 380034 505746 380098
rect 505810 380034 505826 380098
rect 505890 380034 505906 380098
rect 505330 380018 505906 380034
rect 504757 379848 505079 379855
rect 505457 379848 505779 379855
rect 506018 379848 506138 380248
rect 508498 380436 509898 380444
rect 508498 380132 508526 380436
rect 508830 380132 509226 380436
rect 509530 380132 509898 380436
rect 512258 380565 513658 380568
rect 512258 380261 512286 380565
rect 512590 380261 512986 380565
rect 513290 380261 513658 380565
rect 512258 380248 513658 380261
rect 516018 380565 517418 380568
rect 516018 380261 516046 380565
rect 516350 380261 516746 380565
rect 517050 380261 517418 380565
rect 516018 380248 517418 380261
rect 508498 380124 509898 380132
rect 508517 380123 508839 380124
rect 509217 380123 509539 380124
rect 508390 379969 508966 379985
rect 508390 379905 508406 379969
rect 508470 379905 508486 379969
rect 508550 379905 508566 379969
rect 508630 379905 508646 379969
rect 508710 379905 508726 379969
rect 508790 379905 508806 379969
rect 508870 379905 508886 379969
rect 508950 379905 508966 379969
rect 508390 379889 508966 379905
rect 509090 379969 509666 379985
rect 509090 379905 509106 379969
rect 509170 379905 509186 379969
rect 509250 379905 509266 379969
rect 509330 379905 509346 379969
rect 509410 379905 509426 379969
rect 509490 379905 509506 379969
rect 509570 379905 509586 379969
rect 509650 379905 509666 379969
rect 509090 379889 509666 379905
rect 504738 379846 506138 379848
rect 504738 379542 504766 379846
rect 505070 379542 505466 379846
rect 505770 379542 506138 379846
rect 508517 379724 508839 379726
rect 509217 379724 509539 379726
rect 509778 379724 509898 380124
rect 512150 380098 512726 380114
rect 512150 380034 512166 380098
rect 512230 380034 512246 380098
rect 512310 380034 512326 380098
rect 512390 380034 512406 380098
rect 512470 380034 512486 380098
rect 512550 380034 512566 380098
rect 512630 380034 512646 380098
rect 512710 380034 512726 380098
rect 512150 380018 512726 380034
rect 512850 380098 513426 380114
rect 512850 380034 512866 380098
rect 512930 380034 512946 380098
rect 513010 380034 513026 380098
rect 513090 380034 513106 380098
rect 513170 380034 513186 380098
rect 513250 380034 513266 380098
rect 513330 380034 513346 380098
rect 513410 380034 513426 380098
rect 512850 380018 513426 380034
rect 512277 379848 512599 379855
rect 512977 379848 513299 379855
rect 513538 379848 513658 380248
rect 515910 380098 516486 380114
rect 515910 380034 515926 380098
rect 515990 380034 516006 380098
rect 516070 380034 516086 380098
rect 516150 380034 516166 380098
rect 516230 380034 516246 380098
rect 516310 380034 516326 380098
rect 516390 380034 516406 380098
rect 516470 380034 516486 380098
rect 515910 380018 516486 380034
rect 516610 380098 517186 380114
rect 516610 380034 516626 380098
rect 516690 380034 516706 380098
rect 516770 380034 516786 380098
rect 516850 380034 516866 380098
rect 516930 380034 516946 380098
rect 517010 380034 517026 380098
rect 517090 380034 517106 380098
rect 517170 380034 517186 380098
rect 516610 380018 517186 380034
rect 516037 379848 516359 379855
rect 516737 379848 517059 379855
rect 517298 379848 517418 380248
rect 504738 379528 506138 379542
rect 504630 379379 505206 379395
rect 504630 379315 504646 379379
rect 504710 379315 504726 379379
rect 504790 379315 504806 379379
rect 504870 379315 504886 379379
rect 504950 379315 504966 379379
rect 505030 379315 505046 379379
rect 505110 379315 505126 379379
rect 505190 379315 505206 379379
rect 504630 379299 505206 379315
rect 505330 379379 505906 379395
rect 505330 379315 505346 379379
rect 505410 379315 505426 379379
rect 505490 379315 505506 379379
rect 505570 379315 505586 379379
rect 505650 379315 505666 379379
rect 505730 379315 505746 379379
rect 505810 379315 505826 379379
rect 505890 379315 505906 379379
rect 505330 379299 505906 379315
rect 504757 379128 505079 379136
rect 505457 379128 505779 379136
rect 506018 379128 506138 379528
rect 508498 379717 509898 379724
rect 508498 379413 508526 379717
rect 508830 379413 509226 379717
rect 509530 379413 509898 379717
rect 512258 379846 513658 379848
rect 512258 379542 512286 379846
rect 512590 379542 512986 379846
rect 513290 379542 513658 379846
rect 512258 379528 513658 379542
rect 516018 379846 517418 379848
rect 516018 379542 516046 379846
rect 516350 379542 516746 379846
rect 517050 379542 517418 379846
rect 516018 379528 517418 379542
rect 508498 379404 509898 379413
rect 508390 379250 508966 379266
rect 508390 379186 508406 379250
rect 508470 379186 508486 379250
rect 508550 379186 508566 379250
rect 508630 379186 508646 379250
rect 508710 379186 508726 379250
rect 508790 379186 508806 379250
rect 508870 379186 508886 379250
rect 508950 379186 508966 379250
rect 508390 379170 508966 379186
rect 509090 379250 509666 379266
rect 509090 379186 509106 379250
rect 509170 379186 509186 379250
rect 509250 379186 509266 379250
rect 509330 379186 509346 379250
rect 509410 379186 509426 379250
rect 509490 379186 509506 379250
rect 509570 379186 509586 379250
rect 509650 379186 509666 379250
rect 509090 379170 509666 379186
rect 504738 379127 506138 379128
rect 504738 378823 504766 379127
rect 505070 378823 505466 379127
rect 505770 378823 506138 379127
rect 508517 379004 508839 379007
rect 509217 379004 509539 379007
rect 509778 379004 509898 379404
rect 512150 379379 512726 379395
rect 512150 379315 512166 379379
rect 512230 379315 512246 379379
rect 512310 379315 512326 379379
rect 512390 379315 512406 379379
rect 512470 379315 512486 379379
rect 512550 379315 512566 379379
rect 512630 379315 512646 379379
rect 512710 379315 512726 379379
rect 512150 379299 512726 379315
rect 512850 379379 513426 379395
rect 512850 379315 512866 379379
rect 512930 379315 512946 379379
rect 513010 379315 513026 379379
rect 513090 379315 513106 379379
rect 513170 379315 513186 379379
rect 513250 379315 513266 379379
rect 513330 379315 513346 379379
rect 513410 379315 513426 379379
rect 512850 379299 513426 379315
rect 512277 379128 512599 379136
rect 512977 379128 513299 379136
rect 513538 379128 513658 379528
rect 515910 379379 516486 379395
rect 515910 379315 515926 379379
rect 515990 379315 516006 379379
rect 516070 379315 516086 379379
rect 516150 379315 516166 379379
rect 516230 379315 516246 379379
rect 516310 379315 516326 379379
rect 516390 379315 516406 379379
rect 516470 379315 516486 379379
rect 515910 379299 516486 379315
rect 516610 379379 517186 379395
rect 516610 379315 516626 379379
rect 516690 379315 516706 379379
rect 516770 379315 516786 379379
rect 516850 379315 516866 379379
rect 516930 379315 516946 379379
rect 517010 379315 517026 379379
rect 517090 379315 517106 379379
rect 517170 379315 517186 379379
rect 516610 379299 517186 379315
rect 516037 379128 516359 379136
rect 516737 379128 517059 379136
rect 517298 379128 517418 379528
rect 504738 378808 506138 378823
rect 504630 378660 505206 378676
rect 504630 378596 504646 378660
rect 504710 378596 504726 378660
rect 504790 378596 504806 378660
rect 504870 378596 504886 378660
rect 504950 378596 504966 378660
rect 505030 378596 505046 378660
rect 505110 378596 505126 378660
rect 505190 378596 505206 378660
rect 504630 378580 505206 378596
rect 505330 378660 505906 378676
rect 505330 378596 505346 378660
rect 505410 378596 505426 378660
rect 505490 378596 505506 378660
rect 505570 378596 505586 378660
rect 505650 378596 505666 378660
rect 505730 378596 505746 378660
rect 505810 378596 505826 378660
rect 505890 378596 505906 378660
rect 505330 378580 505906 378596
rect 504757 378408 505079 378417
rect 505457 378408 505779 378417
rect 506018 378408 506138 378808
rect 508498 378998 509898 379004
rect 508498 378694 508526 378998
rect 508830 378694 509226 378998
rect 509530 378694 509898 378998
rect 512258 379127 513658 379128
rect 512258 378823 512286 379127
rect 512590 378823 512986 379127
rect 513290 378823 513658 379127
rect 512258 378808 513658 378823
rect 516018 379127 517418 379128
rect 516018 378823 516046 379127
rect 516350 378823 516746 379127
rect 517050 378823 517418 379127
rect 516018 378808 517418 378823
rect 508498 378684 509898 378694
rect 508390 378531 508966 378547
rect 508390 378467 508406 378531
rect 508470 378467 508486 378531
rect 508550 378467 508566 378531
rect 508630 378467 508646 378531
rect 508710 378467 508726 378531
rect 508790 378467 508806 378531
rect 508870 378467 508886 378531
rect 508950 378467 508966 378531
rect 508390 378451 508966 378467
rect 509090 378531 509666 378547
rect 509090 378467 509106 378531
rect 509170 378467 509186 378531
rect 509250 378467 509266 378531
rect 509330 378467 509346 378531
rect 509410 378467 509426 378531
rect 509490 378467 509506 378531
rect 509570 378467 509586 378531
rect 509650 378467 509666 378531
rect 509090 378451 509666 378467
rect 504738 378104 504766 378408
rect 505070 378104 505466 378408
rect 505770 378104 506138 378408
rect 508517 378284 508839 378288
rect 509217 378284 509539 378288
rect 509778 378284 509898 378684
rect 512150 378660 512726 378676
rect 512150 378596 512166 378660
rect 512230 378596 512246 378660
rect 512310 378596 512326 378660
rect 512390 378596 512406 378660
rect 512470 378596 512486 378660
rect 512550 378596 512566 378660
rect 512630 378596 512646 378660
rect 512710 378596 512726 378660
rect 512150 378580 512726 378596
rect 512850 378660 513426 378676
rect 512850 378596 512866 378660
rect 512930 378596 512946 378660
rect 513010 378596 513026 378660
rect 513090 378596 513106 378660
rect 513170 378596 513186 378660
rect 513250 378596 513266 378660
rect 513330 378596 513346 378660
rect 513410 378596 513426 378660
rect 512850 378580 513426 378596
rect 512277 378408 512599 378417
rect 512977 378408 513299 378417
rect 513538 378408 513658 378808
rect 515910 378660 516486 378676
rect 515910 378596 515926 378660
rect 515990 378596 516006 378660
rect 516070 378596 516086 378660
rect 516150 378596 516166 378660
rect 516230 378596 516246 378660
rect 516310 378596 516326 378660
rect 516390 378596 516406 378660
rect 516470 378596 516486 378660
rect 515910 378580 516486 378596
rect 516610 378660 517186 378676
rect 516610 378596 516626 378660
rect 516690 378596 516706 378660
rect 516770 378596 516786 378660
rect 516850 378596 516866 378660
rect 516930 378596 516946 378660
rect 517010 378596 517026 378660
rect 517090 378596 517106 378660
rect 517170 378596 517186 378660
rect 516610 378580 517186 378596
rect 516037 378408 516359 378417
rect 516737 378408 517059 378417
rect 517298 378408 517418 378808
rect 504738 378088 506138 378104
rect 504630 377941 505206 377957
rect 504630 377877 504646 377941
rect 504710 377877 504726 377941
rect 504790 377877 504806 377941
rect 504870 377877 504886 377941
rect 504950 377877 504966 377941
rect 505030 377877 505046 377941
rect 505110 377877 505126 377941
rect 505190 377877 505206 377941
rect 504630 377861 505206 377877
rect 505330 377941 505906 377957
rect 505330 377877 505346 377941
rect 505410 377877 505426 377941
rect 505490 377877 505506 377941
rect 505570 377877 505586 377941
rect 505650 377877 505666 377941
rect 505730 377877 505746 377941
rect 505810 377877 505826 377941
rect 505890 377877 505906 377941
rect 505330 377861 505906 377877
rect 506018 377858 506138 378088
rect 508498 378279 509898 378284
rect 508498 377975 508526 378279
rect 508830 377975 509226 378279
rect 509530 377975 509898 378279
rect 512258 378104 512286 378408
rect 512590 378104 512986 378408
rect 513290 378104 513658 378408
rect 512258 378088 513658 378104
rect 516018 378104 516046 378408
rect 516350 378104 516746 378408
rect 517050 378104 517418 378408
rect 516018 378088 517418 378104
rect 508498 377964 509898 377975
rect 508390 377812 508966 377828
rect 508390 377748 508406 377812
rect 508470 377748 508486 377812
rect 508550 377748 508566 377812
rect 508630 377748 508646 377812
rect 508710 377748 508726 377812
rect 508790 377748 508806 377812
rect 508870 377748 508886 377812
rect 508950 377748 508966 377812
rect 508390 377732 508966 377748
rect 509090 377812 509666 377828
rect 509090 377748 509106 377812
rect 509170 377748 509186 377812
rect 509250 377748 509266 377812
rect 509330 377748 509346 377812
rect 509410 377748 509426 377812
rect 509490 377748 509506 377812
rect 509570 377748 509586 377812
rect 509650 377748 509666 377812
rect 509090 377732 509666 377748
rect 508517 377564 508839 377569
rect 509217 377564 509539 377569
rect 509778 377564 509898 377964
rect 512150 377941 512726 377957
rect 512150 377877 512166 377941
rect 512230 377877 512246 377941
rect 512310 377877 512326 377941
rect 512390 377877 512406 377941
rect 512470 377877 512486 377941
rect 512550 377877 512566 377941
rect 512630 377877 512646 377941
rect 512710 377877 512726 377941
rect 512150 377861 512726 377877
rect 512850 377941 513426 377957
rect 512850 377877 512866 377941
rect 512930 377877 512946 377941
rect 513010 377877 513026 377941
rect 513090 377877 513106 377941
rect 513170 377877 513186 377941
rect 513250 377877 513266 377941
rect 513330 377877 513346 377941
rect 513410 377877 513426 377941
rect 512850 377861 513426 377877
rect 513538 377858 513658 378088
rect 515910 377941 516486 377957
rect 515910 377877 515926 377941
rect 515990 377877 516006 377941
rect 516070 377877 516086 377941
rect 516150 377877 516166 377941
rect 516230 377877 516246 377941
rect 516310 377877 516326 377941
rect 516390 377877 516406 377941
rect 516470 377877 516486 377941
rect 515910 377861 516486 377877
rect 516610 377941 517186 377957
rect 516610 377877 516626 377941
rect 516690 377877 516706 377941
rect 516770 377877 516786 377941
rect 516850 377877 516866 377941
rect 516930 377877 516946 377941
rect 517010 377877 517026 377941
rect 517090 377877 517106 377941
rect 517170 377877 517186 377941
rect 516610 377861 517186 377877
rect 517298 377858 517418 378088
rect 508498 377560 509898 377564
rect 506025 377404 506091 377405
rect 506025 377340 506026 377404
rect 506090 377402 506091 377404
rect 508498 377402 508526 377560
rect 506090 377342 508526 377402
rect 506090 377340 506091 377342
rect 506025 377339 506091 377340
rect 508498 377256 508526 377342
rect 508830 377256 509226 377560
rect 509530 377256 509898 377560
rect 508498 377244 509898 377256
rect 508390 377093 508966 377109
rect 508390 377029 508406 377093
rect 508470 377029 508486 377093
rect 508550 377029 508566 377093
rect 508630 377029 508646 377093
rect 508710 377029 508726 377093
rect 508790 377029 508806 377093
rect 508870 377029 508886 377093
rect 508950 377029 508966 377093
rect 508390 377013 508966 377029
rect 509090 377093 509666 377109
rect 509090 377029 509106 377093
rect 509170 377029 509186 377093
rect 509250 377029 509266 377093
rect 509330 377029 509346 377093
rect 509410 377029 509426 377093
rect 509490 377029 509506 377093
rect 509570 377029 509586 377093
rect 509650 377029 509666 377093
rect 509090 377013 509666 377029
rect 508517 376844 508839 376850
rect 509217 376844 509539 376850
rect 509778 376844 509898 377244
rect 508498 376841 509898 376844
rect 508498 376537 508526 376841
rect 508830 376537 509226 376841
rect 509530 376537 509898 376841
rect 508498 376524 509898 376537
rect 508390 376374 508966 376390
rect 508390 376310 508406 376374
rect 508470 376310 508486 376374
rect 508550 376310 508566 376374
rect 508630 376310 508646 376374
rect 508710 376310 508726 376374
rect 508790 376310 508806 376374
rect 508870 376310 508886 376374
rect 508950 376310 508966 376374
rect 508390 376294 508966 376310
rect 509090 376374 509666 376390
rect 509090 376310 509106 376374
rect 509170 376310 509186 376374
rect 509250 376310 509266 376374
rect 509330 376310 509346 376374
rect 509410 376310 509426 376374
rect 509490 376310 509506 376374
rect 509570 376310 509586 376374
rect 509650 376310 509666 376374
rect 509090 376294 509666 376310
rect 508517 376124 508839 376131
rect 509217 376124 509539 376131
rect 509778 376124 509898 376524
rect 508498 376122 509898 376124
rect 508498 375818 508526 376122
rect 508830 375818 509226 376122
rect 509530 375818 509898 376122
rect 508498 375804 509898 375818
rect 508390 375655 508966 375671
rect 508390 375591 508406 375655
rect 508470 375591 508486 375655
rect 508550 375591 508566 375655
rect 508630 375591 508646 375655
rect 508710 375591 508726 375655
rect 508790 375591 508806 375655
rect 508870 375591 508886 375655
rect 508950 375591 508966 375655
rect 508390 375575 508966 375591
rect 509090 375655 509666 375671
rect 509090 375591 509106 375655
rect 509170 375591 509186 375655
rect 509250 375591 509266 375655
rect 509330 375591 509346 375655
rect 509410 375591 509426 375655
rect 509490 375591 509506 375655
rect 509570 375591 509586 375655
rect 509650 375591 509666 375655
rect 509090 375575 509666 375591
rect 508517 375404 508839 375412
rect 509217 375404 509539 375412
rect 509778 375404 509898 375804
rect 508498 375403 509898 375404
rect 508498 375099 508526 375403
rect 508830 375099 509226 375403
rect 509530 375099 509898 375403
rect 508498 375084 509898 375099
rect 508390 374936 508966 374952
rect 508390 374872 508406 374936
rect 508470 374872 508486 374936
rect 508550 374872 508566 374936
rect 508630 374872 508646 374936
rect 508710 374872 508726 374936
rect 508790 374872 508806 374936
rect 508870 374872 508886 374936
rect 508950 374872 508966 374936
rect 508390 374856 508966 374872
rect 509090 374936 509666 374952
rect 509090 374872 509106 374936
rect 509170 374872 509186 374936
rect 509250 374872 509266 374936
rect 509330 374872 509346 374936
rect 509410 374872 509426 374936
rect 509490 374872 509506 374936
rect 509570 374872 509586 374936
rect 509650 374872 509666 374936
rect 509090 374856 509666 374872
rect 508517 374684 508839 374693
rect 509217 374684 509539 374693
rect 509778 374684 509898 375084
rect 508498 374380 508526 374684
rect 508830 374380 509226 374684
rect 509530 374380 509898 374684
rect 508498 374364 509898 374380
rect 508390 374217 508966 374233
rect 508390 374153 508406 374217
rect 508470 374153 508486 374217
rect 508550 374153 508566 374217
rect 508630 374153 508646 374217
rect 508710 374153 508726 374217
rect 508790 374153 508806 374217
rect 508870 374153 508886 374217
rect 508950 374153 508966 374217
rect 508390 374137 508966 374153
rect 509090 374217 509666 374233
rect 509090 374153 509106 374217
rect 509170 374153 509186 374217
rect 509250 374153 509266 374217
rect 509330 374153 509346 374217
rect 509410 374153 509426 374217
rect 509490 374153 509506 374217
rect 509570 374153 509586 374217
rect 509650 374153 509666 374217
rect 509090 374137 509666 374153
rect 509778 374134 509898 374364
rect 485484 361474 542060 361498
rect 485484 361440 493076 361474
rect 485484 359924 488838 361440
rect 490354 361410 493076 361440
rect 493140 361410 496836 361474
rect 496900 361410 500596 361474
rect 500660 361410 504356 361474
rect 504420 361410 508116 361474
rect 508180 361410 511876 361474
rect 511940 361410 515636 361474
rect 515700 361410 519396 361474
rect 519460 361410 523156 361474
rect 523220 361410 526916 361474
rect 526980 361410 530676 361474
rect 530740 361410 534436 361474
rect 534500 361440 542060 361474
rect 534500 361410 537222 361440
rect 490354 361394 537222 361410
rect 490354 361330 493076 361394
rect 493140 361330 496836 361394
rect 496900 361330 500596 361394
rect 500660 361330 504356 361394
rect 504420 361330 508116 361394
rect 508180 361330 511876 361394
rect 511940 361330 515636 361394
rect 515700 361330 519396 361394
rect 519460 361330 523156 361394
rect 523220 361330 526916 361394
rect 526980 361330 530676 361394
rect 530740 361330 534436 361394
rect 534500 361330 537222 361394
rect 490354 361314 537222 361330
rect 490354 361250 493076 361314
rect 493140 361250 496836 361314
rect 496900 361250 500596 361314
rect 500660 361250 504356 361314
rect 504420 361250 508116 361314
rect 508180 361250 511876 361314
rect 511940 361250 515636 361314
rect 515700 361250 519396 361314
rect 519460 361250 523156 361314
rect 523220 361250 526916 361314
rect 526980 361250 530676 361314
rect 530740 361250 534436 361314
rect 534500 361250 537222 361314
rect 490354 361234 537222 361250
rect 490354 361170 493076 361234
rect 493140 361170 496836 361234
rect 496900 361170 500596 361234
rect 500660 361170 504356 361234
rect 504420 361170 508116 361234
rect 508180 361170 511876 361234
rect 511940 361170 515636 361234
rect 515700 361170 519396 361234
rect 519460 361170 523156 361234
rect 523220 361170 526916 361234
rect 526980 361170 530676 361234
rect 530740 361170 534436 361234
rect 534500 361170 537222 361234
rect 490354 361154 537222 361170
rect 490354 361090 493076 361154
rect 493140 361090 496836 361154
rect 496900 361090 500596 361154
rect 500660 361090 504356 361154
rect 504420 361090 508116 361154
rect 508180 361090 511876 361154
rect 511940 361090 515636 361154
rect 515700 361090 519396 361154
rect 519460 361090 523156 361154
rect 523220 361090 526916 361154
rect 526980 361090 530676 361154
rect 530740 361090 534436 361154
rect 534500 361090 537222 361154
rect 490354 361074 537222 361090
rect 490354 361010 493076 361074
rect 493140 361010 496836 361074
rect 496900 361010 500596 361074
rect 500660 361010 504356 361074
rect 504420 361010 508116 361074
rect 508180 361010 511876 361074
rect 511940 361010 515636 361074
rect 515700 361010 519396 361074
rect 519460 361010 523156 361074
rect 523220 361010 526916 361074
rect 526980 361010 530676 361074
rect 530740 361010 534436 361074
rect 534500 361010 537222 361074
rect 490354 360994 537222 361010
rect 490354 360930 493076 360994
rect 493140 360930 496836 360994
rect 496900 360930 500596 360994
rect 500660 360930 504356 360994
rect 504420 360930 508116 360994
rect 508180 360930 511876 360994
rect 511940 360930 515636 360994
rect 515700 360930 519396 360994
rect 519460 360930 523156 360994
rect 523220 360930 526916 360994
rect 526980 360930 530676 360994
rect 530740 360930 534436 360994
rect 534500 360930 537222 360994
rect 490354 360914 537222 360930
rect 490354 360850 493076 360914
rect 493140 360850 496836 360914
rect 496900 360850 500596 360914
rect 500660 360850 504356 360914
rect 504420 360850 508116 360914
rect 508180 360850 511876 360914
rect 511940 360850 515636 360914
rect 515700 360850 519396 360914
rect 519460 360850 523156 360914
rect 523220 360850 526916 360914
rect 526980 360850 530676 360914
rect 530740 360850 534436 360914
rect 534500 360850 537222 360914
rect 490354 360834 537222 360850
rect 490354 360770 493076 360834
rect 493140 360770 496836 360834
rect 496900 360770 500596 360834
rect 500660 360770 504356 360834
rect 504420 360770 508116 360834
rect 508180 360770 511876 360834
rect 511940 360770 515636 360834
rect 515700 360770 519396 360834
rect 519460 360770 523156 360834
rect 523220 360770 526916 360834
rect 526980 360770 530676 360834
rect 530740 360770 534436 360834
rect 534500 360770 537222 360834
rect 490354 360754 537222 360770
rect 490354 360690 493076 360754
rect 493140 360690 496836 360754
rect 496900 360690 500596 360754
rect 500660 360690 504356 360754
rect 504420 360690 508116 360754
rect 508180 360690 511876 360754
rect 511940 360690 515636 360754
rect 515700 360690 519396 360754
rect 519460 360690 523156 360754
rect 523220 360690 526916 360754
rect 526980 360690 530676 360754
rect 530740 360690 534436 360754
rect 534500 360690 537222 360754
rect 490354 360674 537222 360690
rect 490354 360610 493076 360674
rect 493140 360610 496836 360674
rect 496900 360610 500596 360674
rect 500660 360610 504356 360674
rect 504420 360610 508116 360674
rect 508180 360610 511876 360674
rect 511940 360610 515636 360674
rect 515700 360610 519396 360674
rect 519460 360610 523156 360674
rect 523220 360610 526916 360674
rect 526980 360610 530676 360674
rect 530740 360610 534436 360674
rect 534500 360610 537222 360674
rect 490354 360594 537222 360610
rect 490354 360530 493076 360594
rect 493140 360530 496836 360594
rect 496900 360530 500596 360594
rect 500660 360530 504356 360594
rect 504420 360530 508116 360594
rect 508180 360530 511876 360594
rect 511940 360530 515636 360594
rect 515700 360530 519396 360594
rect 519460 360530 523156 360594
rect 523220 360530 526916 360594
rect 526980 360530 530676 360594
rect 530740 360530 534436 360594
rect 534500 360530 537222 360594
rect 490354 360514 537222 360530
rect 490354 360450 493076 360514
rect 493140 360450 496836 360514
rect 496900 360450 500596 360514
rect 500660 360450 504356 360514
rect 504420 360450 508116 360514
rect 508180 360450 511876 360514
rect 511940 360450 515636 360514
rect 515700 360450 519396 360514
rect 519460 360450 523156 360514
rect 523220 360450 526916 360514
rect 526980 360450 530676 360514
rect 530740 360450 534436 360514
rect 534500 360450 537222 360514
rect 490354 360434 537222 360450
rect 490354 360370 493076 360434
rect 493140 360370 496836 360434
rect 496900 360370 500596 360434
rect 500660 360370 504356 360434
rect 504420 360370 508116 360434
rect 508180 360370 511876 360434
rect 511940 360370 515636 360434
rect 515700 360370 519396 360434
rect 519460 360370 523156 360434
rect 523220 360370 526916 360434
rect 526980 360370 530676 360434
rect 530740 360370 534436 360434
rect 534500 360370 537222 360434
rect 490354 360354 537222 360370
rect 490354 360290 493076 360354
rect 493140 360290 496836 360354
rect 496900 360290 500596 360354
rect 500660 360290 504356 360354
rect 504420 360290 508116 360354
rect 508180 360290 511876 360354
rect 511940 360290 515636 360354
rect 515700 360290 519396 360354
rect 519460 360290 523156 360354
rect 523220 360290 526916 360354
rect 526980 360290 530676 360354
rect 530740 360290 534436 360354
rect 534500 360290 537222 360354
rect 490354 360274 537222 360290
rect 490354 360210 493076 360274
rect 493140 360210 496836 360274
rect 496900 360210 500596 360274
rect 500660 360210 504356 360274
rect 504420 360210 508116 360274
rect 508180 360210 511876 360274
rect 511940 360210 515636 360274
rect 515700 360210 519396 360274
rect 519460 360210 523156 360274
rect 523220 360210 526916 360274
rect 526980 360210 530676 360274
rect 530740 360210 534436 360274
rect 534500 360210 537222 360274
rect 490354 360194 537222 360210
rect 490354 360130 493076 360194
rect 493140 360130 496836 360194
rect 496900 360130 500596 360194
rect 500660 360130 504356 360194
rect 504420 360130 508116 360194
rect 508180 360130 511876 360194
rect 511940 360130 515636 360194
rect 515700 360130 519396 360194
rect 519460 360130 523156 360194
rect 523220 360130 526916 360194
rect 526980 360130 530676 360194
rect 530740 360130 534436 360194
rect 534500 360130 537222 360194
rect 490354 360114 537222 360130
rect 490354 360050 493076 360114
rect 493140 360050 496836 360114
rect 496900 360050 500596 360114
rect 500660 360050 504356 360114
rect 504420 360050 508116 360114
rect 508180 360050 511876 360114
rect 511940 360050 515636 360114
rect 515700 360050 519396 360114
rect 519460 360050 523156 360114
rect 523220 360050 526916 360114
rect 526980 360050 530676 360114
rect 530740 360050 534436 360114
rect 534500 360050 537222 360114
rect 490354 360034 537222 360050
rect 490354 359970 493076 360034
rect 493140 359970 496836 360034
rect 496900 359970 500596 360034
rect 500660 359970 504356 360034
rect 504420 359970 508116 360034
rect 508180 359970 511876 360034
rect 511940 359970 515636 360034
rect 515700 359970 519396 360034
rect 519460 359970 523156 360034
rect 523220 359970 526916 360034
rect 526980 359970 530676 360034
rect 530740 359970 534436 360034
rect 534500 359970 537222 360034
rect 490354 359954 537222 359970
rect 490354 359924 493076 359954
rect 485484 359890 493076 359924
rect 493140 359890 496836 359954
rect 496900 359890 500596 359954
rect 500660 359890 504356 359954
rect 504420 359890 508116 359954
rect 508180 359890 511876 359954
rect 511940 359890 515636 359954
rect 515700 359890 519396 359954
rect 519460 359890 523156 359954
rect 523220 359890 526916 359954
rect 526980 359890 530676 359954
rect 530740 359890 534436 359954
rect 534500 359924 537222 359954
rect 538738 359924 542060 361440
rect 534500 359890 542060 359924
rect 485484 359866 542060 359890
rect 551974 359050 560022 403192
rect 573537 403312 573889 403313
rect 573537 402980 573538 403312
rect 573888 402980 573889 403312
rect 573537 402979 573889 402980
rect 485484 359026 560022 359050
rect 485484 358992 491196 359026
rect 485484 357476 486390 358992
rect 487906 358962 491196 358992
rect 491260 358962 494956 359026
rect 495020 358962 498716 359026
rect 498780 358962 502476 359026
rect 502540 358962 506236 359026
rect 506300 358962 509996 359026
rect 510060 358962 513756 359026
rect 513820 358962 517516 359026
rect 517580 358962 521276 359026
rect 521340 358962 525036 359026
rect 525100 358962 528796 359026
rect 528860 358962 532556 359026
rect 532620 358962 536316 359026
rect 536380 358992 560022 359026
rect 536380 358962 539670 358992
rect 487906 358946 539670 358962
rect 487906 358882 491196 358946
rect 491260 358882 494956 358946
rect 495020 358882 498716 358946
rect 498780 358882 502476 358946
rect 502540 358882 506236 358946
rect 506300 358882 509996 358946
rect 510060 358882 513756 358946
rect 513820 358882 517516 358946
rect 517580 358882 521276 358946
rect 521340 358882 525036 358946
rect 525100 358882 528796 358946
rect 528860 358882 532556 358946
rect 532620 358882 536316 358946
rect 536380 358882 539670 358946
rect 487906 358866 539670 358882
rect 487906 358802 491196 358866
rect 491260 358802 494956 358866
rect 495020 358802 498716 358866
rect 498780 358802 502476 358866
rect 502540 358802 506236 358866
rect 506300 358802 509996 358866
rect 510060 358802 513756 358866
rect 513820 358802 517516 358866
rect 517580 358802 521276 358866
rect 521340 358802 525036 358866
rect 525100 358802 528796 358866
rect 528860 358802 532556 358866
rect 532620 358802 536316 358866
rect 536380 358802 539670 358866
rect 487906 358786 539670 358802
rect 487906 358722 491196 358786
rect 491260 358722 494956 358786
rect 495020 358722 498716 358786
rect 498780 358722 502476 358786
rect 502540 358722 506236 358786
rect 506300 358722 509996 358786
rect 510060 358722 513756 358786
rect 513820 358722 517516 358786
rect 517580 358722 521276 358786
rect 521340 358722 525036 358786
rect 525100 358722 528796 358786
rect 528860 358722 532556 358786
rect 532620 358722 536316 358786
rect 536380 358722 539670 358786
rect 487906 358706 539670 358722
rect 487906 358642 491196 358706
rect 491260 358642 494956 358706
rect 495020 358642 498716 358706
rect 498780 358642 502476 358706
rect 502540 358642 506236 358706
rect 506300 358642 509996 358706
rect 510060 358642 513756 358706
rect 513820 358642 517516 358706
rect 517580 358642 521276 358706
rect 521340 358642 525036 358706
rect 525100 358642 528796 358706
rect 528860 358642 532556 358706
rect 532620 358642 536316 358706
rect 536380 358642 539670 358706
rect 487906 358626 539670 358642
rect 487906 358562 491196 358626
rect 491260 358562 494956 358626
rect 495020 358562 498716 358626
rect 498780 358562 502476 358626
rect 502540 358562 506236 358626
rect 506300 358562 509996 358626
rect 510060 358562 513756 358626
rect 513820 358562 517516 358626
rect 517580 358562 521276 358626
rect 521340 358562 525036 358626
rect 525100 358562 528796 358626
rect 528860 358562 532556 358626
rect 532620 358562 536316 358626
rect 536380 358562 539670 358626
rect 487906 358546 539670 358562
rect 487906 358482 491196 358546
rect 491260 358482 494956 358546
rect 495020 358482 498716 358546
rect 498780 358482 502476 358546
rect 502540 358482 506236 358546
rect 506300 358482 509996 358546
rect 510060 358482 513756 358546
rect 513820 358482 517516 358546
rect 517580 358482 521276 358546
rect 521340 358482 525036 358546
rect 525100 358482 528796 358546
rect 528860 358482 532556 358546
rect 532620 358482 536316 358546
rect 536380 358482 539670 358546
rect 487906 358466 539670 358482
rect 487906 358402 491196 358466
rect 491260 358402 494956 358466
rect 495020 358402 498716 358466
rect 498780 358402 502476 358466
rect 502540 358402 506236 358466
rect 506300 358402 509996 358466
rect 510060 358402 513756 358466
rect 513820 358402 517516 358466
rect 517580 358402 521276 358466
rect 521340 358402 525036 358466
rect 525100 358402 528796 358466
rect 528860 358402 532556 358466
rect 532620 358402 536316 358466
rect 536380 358402 539670 358466
rect 487906 358386 539670 358402
rect 487906 358322 491196 358386
rect 491260 358322 494956 358386
rect 495020 358322 498716 358386
rect 498780 358322 502476 358386
rect 502540 358322 506236 358386
rect 506300 358322 509996 358386
rect 510060 358322 513756 358386
rect 513820 358322 517516 358386
rect 517580 358322 521276 358386
rect 521340 358322 525036 358386
rect 525100 358322 528796 358386
rect 528860 358322 532556 358386
rect 532620 358322 536316 358386
rect 536380 358322 539670 358386
rect 487906 358306 539670 358322
rect 487906 358242 491196 358306
rect 491260 358242 494956 358306
rect 495020 358242 498716 358306
rect 498780 358242 502476 358306
rect 502540 358242 506236 358306
rect 506300 358242 509996 358306
rect 510060 358242 513756 358306
rect 513820 358242 517516 358306
rect 517580 358242 521276 358306
rect 521340 358242 525036 358306
rect 525100 358242 528796 358306
rect 528860 358242 532556 358306
rect 532620 358242 536316 358306
rect 536380 358242 539670 358306
rect 487906 358226 539670 358242
rect 487906 358162 491196 358226
rect 491260 358162 494956 358226
rect 495020 358162 498716 358226
rect 498780 358162 502476 358226
rect 502540 358162 506236 358226
rect 506300 358162 509996 358226
rect 510060 358162 513756 358226
rect 513820 358162 517516 358226
rect 517580 358162 521276 358226
rect 521340 358162 525036 358226
rect 525100 358162 528796 358226
rect 528860 358162 532556 358226
rect 532620 358162 536316 358226
rect 536380 358162 539670 358226
rect 487906 358146 539670 358162
rect 487906 358082 491196 358146
rect 491260 358082 494956 358146
rect 495020 358082 498716 358146
rect 498780 358082 502476 358146
rect 502540 358082 506236 358146
rect 506300 358082 509996 358146
rect 510060 358082 513756 358146
rect 513820 358082 517516 358146
rect 517580 358082 521276 358146
rect 521340 358082 525036 358146
rect 525100 358082 528796 358146
rect 528860 358082 532556 358146
rect 532620 358082 536316 358146
rect 536380 358082 539670 358146
rect 487906 358066 539670 358082
rect 487906 358002 491196 358066
rect 491260 358002 494956 358066
rect 495020 358002 498716 358066
rect 498780 358002 502476 358066
rect 502540 358002 506236 358066
rect 506300 358002 509996 358066
rect 510060 358002 513756 358066
rect 513820 358002 517516 358066
rect 517580 358002 521276 358066
rect 521340 358002 525036 358066
rect 525100 358002 528796 358066
rect 528860 358002 532556 358066
rect 532620 358002 536316 358066
rect 536380 358002 539670 358066
rect 487906 357986 539670 358002
rect 487906 357922 491196 357986
rect 491260 357922 494956 357986
rect 495020 357922 498716 357986
rect 498780 357922 502476 357986
rect 502540 357922 506236 357986
rect 506300 357922 509996 357986
rect 510060 357922 513756 357986
rect 513820 357922 517516 357986
rect 517580 357922 521276 357986
rect 521340 357922 525036 357986
rect 525100 357922 528796 357986
rect 528860 357922 532556 357986
rect 532620 357922 536316 357986
rect 536380 357922 539670 357986
rect 487906 357906 539670 357922
rect 487906 357842 491196 357906
rect 491260 357842 494956 357906
rect 495020 357842 498716 357906
rect 498780 357842 502476 357906
rect 502540 357842 506236 357906
rect 506300 357842 509996 357906
rect 510060 357842 513756 357906
rect 513820 357842 517516 357906
rect 517580 357842 521276 357906
rect 521340 357842 525036 357906
rect 525100 357842 528796 357906
rect 528860 357842 532556 357906
rect 532620 357842 536316 357906
rect 536380 357842 539670 357906
rect 487906 357826 539670 357842
rect 487906 357762 491196 357826
rect 491260 357762 494956 357826
rect 495020 357762 498716 357826
rect 498780 357762 502476 357826
rect 502540 357762 506236 357826
rect 506300 357762 509996 357826
rect 510060 357762 513756 357826
rect 513820 357762 517516 357826
rect 517580 357762 521276 357826
rect 521340 357762 525036 357826
rect 525100 357762 528796 357826
rect 528860 357762 532556 357826
rect 532620 357762 536316 357826
rect 536380 357762 539670 357826
rect 487906 357746 539670 357762
rect 487906 357682 491196 357746
rect 491260 357682 494956 357746
rect 495020 357682 498716 357746
rect 498780 357682 502476 357746
rect 502540 357682 506236 357746
rect 506300 357682 509996 357746
rect 510060 357682 513756 357746
rect 513820 357682 517516 357746
rect 517580 357682 521276 357746
rect 521340 357682 525036 357746
rect 525100 357682 528796 357746
rect 528860 357682 532556 357746
rect 532620 357682 536316 357746
rect 536380 357682 539670 357746
rect 487906 357666 539670 357682
rect 487906 357602 491196 357666
rect 491260 357602 494956 357666
rect 495020 357602 498716 357666
rect 498780 357602 502476 357666
rect 502540 357602 506236 357666
rect 506300 357602 509996 357666
rect 510060 357602 513756 357666
rect 513820 357602 517516 357666
rect 517580 357602 521276 357666
rect 521340 357602 525036 357666
rect 525100 357602 528796 357666
rect 528860 357602 532556 357666
rect 532620 357602 536316 357666
rect 536380 357602 539670 357666
rect 487906 357586 539670 357602
rect 487906 357522 491196 357586
rect 491260 357522 494956 357586
rect 495020 357522 498716 357586
rect 498780 357522 502476 357586
rect 502540 357522 506236 357586
rect 506300 357522 509996 357586
rect 510060 357522 513756 357586
rect 513820 357522 517516 357586
rect 517580 357522 521276 357586
rect 521340 357522 525036 357586
rect 525100 357522 528796 357586
rect 528860 357522 532556 357586
rect 532620 357522 536316 357586
rect 536380 357522 539670 357586
rect 487906 357506 539670 357522
rect 487906 357476 491196 357506
rect 485484 357442 491196 357476
rect 491260 357442 494956 357506
rect 495020 357442 498716 357506
rect 498780 357442 502476 357506
rect 502540 357442 506236 357506
rect 506300 357442 509996 357506
rect 510060 357442 513756 357506
rect 513820 357442 517516 357506
rect 517580 357442 521276 357506
rect 521340 357442 525036 357506
rect 525100 357442 528796 357506
rect 528860 357442 532556 357506
rect 532620 357442 536316 357506
rect 536380 357476 539670 357506
rect 541186 358052 560022 358992
rect 541186 357844 559712 358052
rect 559920 357844 560022 358052
rect 541186 357476 560022 357844
rect 573539 357920 573879 357921
rect 573539 357594 573540 357920
rect 573878 357594 573879 357920
rect 573539 357593 573879 357594
rect 536380 357442 560022 357476
rect 485484 357418 560022 357442
rect 551974 311744 560022 357418
rect 551974 311536 559652 311744
rect 559860 311536 560022 311744
rect 551974 154934 560022 311536
rect 573491 311700 573835 311701
rect 573491 311420 573492 311700
rect 573834 311420 573835 311700
rect 573491 311419 573835 311420
<< via4 >>
rect 567306 640080 573722 644324
rect 567306 630012 573722 634256
rect 573564 491888 573874 492160
rect 486390 412480 487906 413996
rect 539670 412480 541186 413996
rect 488838 410032 490354 411548
rect 537222 410032 538738 411548
rect 488838 359924 490354 361440
rect 537222 359924 538738 361440
rect 573538 402980 573888 403312
rect 486390 357476 487906 358992
rect 539670 357476 541186 358992
rect 573540 357594 573878 357920
rect 573492 311420 573834 311700
<< metal5 >>
rect 567158 644324 573920 649062
rect 567158 640080 567306 644324
rect 573722 640080 573920 644324
rect 567158 634256 573920 640080
rect 567158 630012 567306 634256
rect 573722 630012 573920 634256
rect 567158 627314 573920 630012
rect 567156 621952 573942 627314
rect 567158 492160 573920 621952
rect 567158 491888 573564 492160
rect 573874 491888 573920 492160
rect 488780 422974 490412 423442
rect 567158 422974 573920 491888
rect 488780 421342 573920 422974
rect 486332 413996 487964 414954
rect 486332 412480 486390 413996
rect 487906 412480 487964 413996
rect 486332 358992 487964 412480
rect 486332 357476 486390 358992
rect 487906 357476 487964 358992
rect 486332 356442 487964 357476
rect 488780 411548 490412 421342
rect 536984 420968 573920 421342
rect 488780 410032 488838 411548
rect 490354 410032 490412 411548
rect 488780 361440 490412 410032
rect 488780 359924 488838 361440
rect 490354 359924 490412 361440
rect 488780 348924 490412 359924
rect 537164 411548 538796 420968
rect 537164 410032 537222 411548
rect 538738 410032 538796 411548
rect 537164 361440 538796 410032
rect 537164 359924 537222 361440
rect 538738 359924 538796 361440
rect 537164 348924 538796 359924
rect 539612 413996 541244 414954
rect 539612 412480 539670 413996
rect 541186 412480 541244 413996
rect 539612 358992 541244 412480
rect 539612 357476 539670 358992
rect 541186 357476 541244 358992
rect 539612 356442 541244 357476
rect 567158 403312 573920 420968
rect 567158 402980 573538 403312
rect 573888 402980 573920 403312
rect 567158 357920 573920 402980
rect 567158 357594 573540 357920
rect 573878 357594 573920 357920
rect 567158 348924 573920 357594
rect 488668 347292 573920 348924
rect 567158 311700 573920 347292
rect 567158 311420 573492 311700
rect 573834 311420 573920 311700
rect 567158 147385 573920 311420
<< labels >>
flabel metal3 510596 697782 515352 701406 1 FreeSans 8000 0 0 0 VSSA1
flabel metal3 574704 639800 581232 644606 1 FreeSans 8000 0 0 0 VCCD1
flabel metal1 565560 313022 565620 313082 1 FreeSans 800 0 0 0 nmos_flat_3/VPWR
flabel metal1 565560 311142 565620 311202 1 FreeSans 800 0 0 0 nmos_flat_3/VGND
flabel locali 560404 312862 560464 312922 1 FreeSans 800 0 0 0 nmos_flat_3/SOURCE
flabel locali 560404 311542 560464 311602 1 FreeSans 800 0 0 0 nmos_flat_3/DRAIN
flabel locali 560404 311376 560464 311436 1 FreeSans 800 0 0 0 nmos_flat_3/GATE
flabel nwell 580418 313092 580478 313152 1 FreeSans 800 0 0 0 pmos_flat_2/VPWR
flabel metal1 580320 311212 580478 311272 1 FreeSans 800 0 0 0 pmos_flat_2/VGND
flabel locali 575092 312932 575152 312972 1 FreeSans 800 0 0 0 pmos_flat_2/SOURCE
flabel locali 575092 311552 575152 311612 1 FreeSans 800 0 0 0 pmos_flat_2/DRAIN
flabel locali 575092 311390 575152 311450 1 FreeSans 800 0 0 0 pmos_flat_2/GATE
rlabel metal5 539612 413322 541244 414954 4 bgr_top_flat_0/VSS
rlabel metal5 537164 413322 538796 414954 4 bgr_top_flat_0/VDD
flabel metal1 534928 364678 535048 364798 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_2/Rin
flabel metal1 535888 364678 536008 364798 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_2/Rout
flabel metal1 534438 364858 534498 364918 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_2/VPWR
flabel metal1 536318 364858 536378 364918 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_2/VGND
flabel metal1 534928 370166 535048 370286 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_1/Rin
flabel metal1 535888 370166 536008 370286 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_1/Rout
flabel metal1 534438 370346 534498 370406 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_1/VPWR
flabel metal1 536318 370346 536378 370406 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_1/VGND
flabel metal1 534928 367422 535048 367542 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_0/Rin
flabel metal1 535888 367422 536008 367542 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_0/Rout
flabel metal1 534438 367602 534498 367662 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_0/VPWR
flabel metal1 536318 367602 536378 367662 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_0/VGND
flabel metal1 531168 370950 531288 371070 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_3/Rin
flabel metal1 532128 370950 532248 371070 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_3/Rout
flabel metal1 530678 371130 530738 371190 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_3/VPWR
flabel metal1 532558 371130 532618 371190 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_3/VGND
flabel metal1 531168 368206 531288 368326 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_4/Rin
flabel metal1 532128 368206 532248 368326 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_4/Rout
flabel metal1 530678 368386 530738 368446 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_4/VPWR
flabel metal1 532558 368386 532618 368446 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_4/VGND
flabel metal1 531168 365462 531288 365582 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_5/Rin
flabel metal1 532128 365462 532248 365582 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_5/Rout
flabel metal1 530678 365642 530738 365702 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_5/VPWR
flabel metal1 532558 365642 532618 365702 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_5/VGND
flabel metal1 527408 370852 527528 370972 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_6/Rin
flabel metal1 528368 370852 528488 370972 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_6/Rout
flabel metal1 526918 371032 526978 371092 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_6/VPWR
flabel metal1 528798 371032 528858 371092 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_6/VGND
flabel metal1 527408 368108 527528 368228 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_7/Rin
flabel metal1 528368 368108 528488 368228 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_7/Rout
flabel metal1 526918 368288 526978 368348 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_7/VPWR
flabel metal1 528798 368288 528858 368348 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_7/VGND
flabel metal1 527408 365364 527528 365484 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_8/Rin
flabel metal1 528368 365364 528488 365484 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_8/Rout
flabel metal1 526918 365544 526978 365604 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_8/VPWR
flabel metal1 528798 365544 528858 365604 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_8/VGND
flabel locali 524904 362516 524964 362576 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_60_0/GATE
flabel locali 523338 362516 523378 362576 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_60_0/SOURCE
flabel locali 524798 362516 524858 362576 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_60_0/DRAIN
flabel nwell 523158 390162 523218 390222 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_60_0/VPWR
flabel metal1 525038 390064 525098 390222 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_60_0/VGND
flabel metal1 519888 390844 520008 390964 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_10/Rin
flabel metal1 520848 390844 520968 390964 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_10/Rout
flabel metal1 519398 391024 519458 391084 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_10/VPWR
flabel metal1 521278 391024 521338 391084 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_10/VGND
flabel metal1 519888 387512 520008 387632 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_9/Rin
flabel metal1 520848 387512 520968 387632 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_9/Rout
flabel metal1 519398 387692 519458 387752 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_9/VPWR
flabel metal1 521278 387692 521338 387752 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_9/VGND
flabel metal1 519888 366344 520008 366464 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_15/Rin
flabel metal1 520848 366344 520968 366464 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_15/Rout
flabel metal1 519398 366524 519458 366584 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_15/VPWR
flabel metal1 521278 366524 521338 366584 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_15/VGND
flabel metal1 519888 374576 520008 374696 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_14/Rin
flabel metal1 520848 374576 520968 374696 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_14/Rout
flabel metal1 519398 374756 519458 374816 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_14/VPWR
flabel metal1 521278 374756 521338 374816 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_14/VGND
flabel metal1 519888 377320 520008 377440 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_13/Rin
flabel metal1 520848 377320 520968 377440 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_13/Rout
flabel metal1 519398 377500 519458 377560 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_13/VPWR
flabel metal1 521278 377500 521338 377560 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_13/VGND
flabel metal1 519888 381534 520008 381654 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_12/Rin
flabel metal1 520848 381534 520968 381654 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_12/Rout
flabel metal1 519398 381714 519458 381774 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_12/VPWR
flabel metal1 521278 381714 521338 381774 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_12/VGND
flabel metal1 519888 384768 520008 384888 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_11/Rin
flabel metal1 520848 384768 520968 384888 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_11/Rout
flabel metal1 519398 384948 519458 385008 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_11/VPWR
flabel metal1 521278 384948 521338 385008 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_11/VGND
flabel locali 517184 385356 517244 385416 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_9_0/GATE
flabel locali 515798 385356 515858 385416 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_9_0/SOURCE
flabel locali 517018 385356 517078 385416 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_9_0/DRAIN
flabel metal1 515638 389476 515698 389536 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_9_0/VPWR
flabel metal1 517518 389476 517578 389536 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_9_0/VGND
flabel metal1 516128 392314 516248 392434 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_16/Rin
flabel metal1 517088 392314 517208 392434 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_16/Rout
flabel metal1 515638 392494 515698 392554 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_16/VPWR
flabel metal1 517518 392494 517578 392554 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_16/VGND
flabel metal2 515898 384828 515978 385028 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_0/Cin
flabel metal4 517308 384846 517408 385006 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_0/Cout
flabel metal1 515638 384966 515698 385026 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_0/VPWR
flabel metal1 517518 384966 517578 385026 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_0/VGND
flabel metal1 516128 371832 516248 371952 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_19/Rin
flabel metal1 517088 371832 517208 371952 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_19/Rout
flabel metal1 515638 372012 515698 372072 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_19/VPWR
flabel metal1 517518 372012 517578 372072 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_19/VGND
flabel metal1 516128 374576 516248 374696 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_18/Rin
flabel metal1 517088 374576 517208 374696 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_18/Rout
flabel metal1 515638 374756 515698 374816 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_18/VPWR
flabel metal1 517518 374756 517578 374816 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_18/VGND
flabel metal1 516128 377320 516248 377440 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_17/Rin
flabel metal1 517088 377320 517208 377440 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_17/Rout
flabel metal1 515638 377500 515698 377560 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_17/VPWR
flabel metal1 517518 377500 517578 377560 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_17/VGND
flabel metal1 516128 366344 516248 366464 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rin
flabel metal1 517088 366344 517208 366464 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout
flabel metal1 515638 366524 515698 366584 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/VPWR
flabel metal1 517518 366524 517578 366584 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/VGND
flabel metal1 516128 369088 516248 369208 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_20/Rin
flabel metal1 517088 369088 517208 369208 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_20/Rout
flabel metal1 515638 369268 515698 369328 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_20/VPWR
flabel metal1 517518 369268 517578 369328 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_20/VGND
flabel metal1 512368 392706 512488 392826 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_25/Rin
flabel metal1 513328 392706 513448 392826 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_25/Rout
flabel metal1 511878 392886 511938 392946 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_25/VPWR
flabel metal1 513758 392886 513818 392946 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_25/VGND
flabel metal1 512368 398194 512488 398314 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_24/Rin
flabel metal1 513328 398194 513448 398314 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_24/Rout
flabel metal1 511878 398374 511938 398434 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_24/VPWR
flabel metal1 513758 398374 513818 398434 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_24/VGND
flabel metal1 512368 395450 512488 395570 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_23/Rin
flabel metal1 513328 395450 513448 395570 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_23/Rout
flabel metal1 511878 395630 511938 395690 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_23/VPWR
flabel metal1 513758 395630 513818 395690 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_23/VGND
flabel metal1 512368 387512 512488 387632 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_22/Rin
flabel metal1 513328 387512 513448 387632 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_22/Rout
flabel metal1 511878 387692 511938 387752 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_22/VPWR
flabel metal1 513758 387692 513818 387752 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_22/VGND
flabel metal2 512138 384828 512218 385028 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_1/Cin
flabel metal4 513548 384846 513648 385006 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_1/Cout
flabel metal1 511878 384966 511938 385026 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_1/VPWR
flabel metal1 513758 384966 513818 385026 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_1/VGND
flabel locali 513624 374606 513684 374666 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_0/GATE
flabel locali 512058 374606 512098 374666 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_0/SOURCE
flabel locali 513518 374606 513578 374666 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_0/DRAIN
flabel nwell 511878 377520 511938 377580 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_0/VPWR
flabel metal1 513758 377422 513818 377580 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_0/VGND
flabel locali 512788 362988 512892 363236 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Emitter
flabel locali 512217 363076 512266 363177 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector
flabel locali 512376 363082 512416 363200 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base
flabel locali 512788 364328 512892 364576 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 512217 364416 512266 364517 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 512376 364422 512416 364540 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 512788 365668 512892 365916 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 512217 365756 512266 365857 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 512376 365762 512416 365880 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 512788 367008 512892 367256 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 512217 367096 512266 367197 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 512376 367102 512416 367220 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 512788 368348 512892 368596 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 512217 368436 512266 368537 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 512376 368442 512416 368560 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 512788 369688 512892 369936 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 512217 369776 512266 369877 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 512376 369782 512416 369900 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 512788 371028 512892 371276 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 512217 371116 512266 371217 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 512376 371122 512416 371240 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 512788 372368 512892 372616 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/xm1/Emitter
flabel locali 512217 372456 512266 372557 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/xm1/Collector
flabel locali 512376 372462 512416 372580 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/xm1/Base
flabel metal1 512648 372390 512778 372630 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/Emitter
flabel metal1 512376 372740 512416 372980 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/Base
flabel metal1 512224 372904 512264 373144 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/Collector
flabel metal1 511878 373110 511938 373170 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/VPWR
flabel metal1 513758 373110 513818 373170 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_0/VGND
flabel metal2 508378 388552 508458 388752 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_2/Cin
flabel metal4 509788 388570 509888 388730 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_2/Cout
flabel metal1 508118 388690 508178 388750 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_2/VPWR
flabel metal1 509998 388690 510058 388750 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_2/VGND
flabel metal1 508608 392705 508728 392825 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_0/Rin
flabel metal1 509568 392705 509688 392825 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_0/Rout
flabel metal1 508118 392884 508178 392944 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_0/VPWR
flabel metal1 509998 392884 510058 392944 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_0/VGND
flabel metal1 508608 395450 508728 395570 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_26/Rin
flabel metal1 509568 395450 509688 395570 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_26/Rout
flabel metal1 508118 395630 508178 395690 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_26/VPWR
flabel metal1 509998 395630 510058 395690 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_26/VGND
flabel locali 509028 362988 509132 363236 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Emitter
flabel locali 508457 363076 508506 363177 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector
flabel locali 508616 363082 508656 363200 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base
flabel locali 509028 364328 509132 364576 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 508457 364416 508506 364517 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 508616 364422 508656 364540 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 509028 365668 509132 365916 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 508457 365756 508506 365857 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 508616 365762 508656 365880 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 509028 367008 509132 367256 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 508457 367096 508506 367197 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 508616 367102 508656 367220 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 509028 368348 509132 368596 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 508457 368436 508506 368537 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 508616 368442 508656 368560 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 509028 369688 509132 369936 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 508457 369776 508506 369877 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 508616 369782 508656 369900 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 509028 371028 509132 371276 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 508457 371116 508506 371217 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 508616 371122 508656 371240 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 509028 372368 509132 372616 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/xm1/Emitter
flabel locali 508457 372456 508506 372557 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/xm1/Collector
flabel locali 508616 372462 508656 372580 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/xm1/Base
flabel metal1 508888 372390 509018 372630 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/Emitter
flabel metal1 508616 372740 508656 372980 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/Base
flabel metal1 508464 372904 508504 373144 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/Collector
flabel metal1 508118 373110 508178 373170 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/VPWR
flabel metal1 509998 373110 510058 373170 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_1/VGND
flabel metal2 508378 381104 508458 381304 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_3/Cin
flabel metal4 509788 381122 509888 381282 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_3/Cout
flabel metal1 508118 381242 508178 381302 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_3/VPWR
flabel metal1 509998 381242 510058 381302 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_3/VGND
flabel metal1 504848 401036 504968 401156 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_27/Rin
flabel metal1 505808 401036 505928 401156 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_27/Rout
flabel metal1 504358 401216 504418 401276 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_27/VPWR
flabel metal1 506238 401216 506298 401276 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_27/VGND
flabel locali 505268 402160 505372 402408 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_1_0/xm1/Emitter
flabel locali 504697 402248 504746 402349 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_1_0/xm1/Collector
flabel locali 504856 402254 504896 402372 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_1_0/xm1/Base
flabel locali 505128 402172 505258 402400 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_1_0/Emitter
flabel locali 504856 402068 504896 402188 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_1_0/Base
flabel locali 504704 402032 504744 402152 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_1_0/Collector
flabel metal1 504358 402902 504418 402962 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_1_0/VPWR
flabel metal1 506238 402902 506298 402962 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_1_0/VGND
flabel metal1 504848 398292 504968 398412 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_28/Rin
flabel metal1 505808 398292 505928 398412 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_28/Rout
flabel metal1 504358 398472 504418 398532 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_28/VPWR
flabel metal1 506238 398472 506298 398532 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_28/VGND
flabel metal1 504848 395547 504968 395667 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_1/Rin
flabel metal1 505808 395547 505928 395667 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_1/Rout
flabel metal1 504358 395726 504418 395786 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_1/VPWR
flabel metal1 506238 395726 506298 395786 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_1/VGND
flabel locali 505904 385356 505964 385416 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_9_1/GATE
flabel locali 504518 385356 504578 385416 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_9_1/SOURCE
flabel locali 505738 385356 505798 385416 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_9_1/DRAIN
flabel metal1 504358 389476 504418 389536 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_9_1/VPWR
flabel metal1 506238 389476 506298 389536 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_9_1/VGND
flabel metal1 504848 392216 504968 392336 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_29/Rin
flabel metal1 505808 392216 505928 392336 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_29/Rout
flabel metal1 504358 392396 504418 392456 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_29/VPWR
flabel metal1 506238 392396 506298 392456 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_29/VGND
flabel metal2 504618 384828 504698 385028 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cin
flabel metal4 506028 384846 506128 385006 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout
flabel metal1 504358 384966 504418 385026 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/VPWR
flabel metal1 506238 384966 506298 385026 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/VGND
flabel locali 506104 374606 506164 374666 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE
flabel locali 504538 374606 504578 374666 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/SOURCE
flabel locali 505998 374606 506058 374666 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/DRAIN
flabel nwell 504358 377520 504418 377580 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/VPWR
flabel metal1 506238 377422 506298 377580 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/VGND
flabel locali 505268 362988 505372 363236 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Emitter
flabel locali 504697 363076 504746 363177 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector
flabel locali 504856 363082 504896 363200 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base
flabel locali 505268 364328 505372 364576 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 504697 364416 504746 364517 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 504856 364422 504896 364540 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 505268 365668 505372 365916 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 504697 365756 504746 365857 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 504856 365762 504896 365880 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 505268 367008 505372 367256 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 504697 367096 504746 367197 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 504856 367102 504896 367220 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 505268 368348 505372 368596 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 504697 368436 504746 368537 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 504856 368442 504896 368560 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 505268 369688 505372 369936 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 504697 369776 504746 369877 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 504856 369782 504896 369900 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 505268 371028 505372 371276 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 504697 371116 504746 371217 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 504856 371122 504896 371240 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 505268 372368 505372 372616 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/xm1/Emitter
flabel locali 504697 372456 504746 372557 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/xm1/Collector
flabel locali 504856 372462 504896 372580 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/xm1/Base
flabel metal1 505128 372390 505258 372630 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/Emitter
flabel metal1 504856 372740 504896 372980 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/Base
flabel metal1 504704 372904 504744 373144 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/Collector
flabel metal1 504358 373110 504418 373170 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/VPWR
flabel metal1 506238 373110 506298 373170 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_2/VGND
flabel metal2 500858 408446 500938 408646 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_5/Cin
flabel metal4 502268 408464 502368 408624 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_5/Cout
flabel metal1 500598 408584 500658 408644 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_5/VPWR
flabel metal1 502478 408584 502538 408644 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_5/VGND
flabel metal2 500858 399626 500938 399826 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_6/Cin
flabel metal4 502268 399644 502368 399804 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_6/Cout
flabel metal1 500598 399764 500658 399824 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_6/VPWR
flabel metal1 502478 399764 502538 399824 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_6/VGND
flabel locali 502344 386656 502404 386716 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_12_0/GATE
flabel locali 500778 386656 500818 386716 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_12_0/SOURCE
flabel locali 502238 386656 502298 386716 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_12_0/DRAIN
flabel nwell 500598 392318 500658 392378 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_12_0/VPWR
flabel metal1 502478 392220 502538 392378 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_12_0/VGND
flabel locali 502344 379992 502404 380052 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_12_1/GATE
flabel locali 500778 379992 500818 380052 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_12_1/SOURCE
flabel locali 502238 379992 502298 380052 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_12_1/DRAIN
flabel nwell 500598 385654 500658 385714 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_12_1/VPWR
flabel metal1 502478 385556 502538 385714 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_12_1/VGND
flabel locali 502144 373498 502204 373558 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_9_2/GATE
flabel locali 500758 373498 500818 373558 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_9_2/SOURCE
flabel locali 501978 373498 502038 373558 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_9_2/DRAIN
flabel metal1 500598 377618 500658 377678 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_9_2/VPWR
flabel metal1 502478 377618 502538 377678 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_9_2/VGND
flabel locali 501508 362988 501612 363236 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Emitter
flabel locali 500937 363076 500986 363177 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector
flabel locali 501096 363082 501136 363200 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base
flabel locali 501508 364328 501612 364576 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 500937 364416 500986 364517 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 501096 364422 501136 364540 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 501508 365668 501612 365916 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 500937 365756 500986 365857 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 501096 365762 501136 365880 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 501508 367008 501612 367256 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 500937 367096 500986 367197 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 501096 367102 501136 367220 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 501508 368348 501612 368596 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 500937 368436 500986 368537 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 501096 368442 501136 368560 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 501508 369688 501612 369936 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 500937 369776 500986 369877 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 501096 369782 501136 369900 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 501508 371028 501612 371276 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 500937 371116 500986 371217 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 501096 371122 501136 371240 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 501508 372368 501612 372616 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/xm1/Emitter
flabel locali 500937 372456 500986 372557 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/xm1/Collector
flabel locali 501096 372462 501136 372580 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/xm1/Base
flabel metal1 501368 372390 501498 372630 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/Emitter
flabel metal1 501096 372740 501136 372980 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/Base
flabel metal1 500944 372904 500984 373144 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/Collector
flabel metal1 500598 373110 500658 373170 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/VPWR
flabel metal1 502478 373110 502538 373170 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_8_3/VGND
flabel locali 498544 400320 498604 400380 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/GATE
flabel locali 496998 400320 497058 400380 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/SOURCE
flabel locali 498318 400320 498378 400380 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN
flabel metal1 496838 400776 496898 400836 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/VPWR
flabel metal1 498718 400776 498778 400836 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/VGND
flabel metal2 497098 408838 497178 409038 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_7/Cin
flabel metal4 498508 408856 498608 409016 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_7/Cout
flabel metal1 496838 408976 496898 409036 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_7/VPWR
flabel metal1 498718 408976 498778 409036 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_7/VGND
flabel locali 498584 372316 498644 372376 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_60_1/GATE
flabel locali 497018 372316 497058 372376 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_60_1/SOURCE
flabel locali 498478 372316 498538 372376 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_60_1/DRAIN
flabel nwell 496838 399962 496898 400022 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_60_1/VPWR
flabel metal1 498718 399864 498778 400022 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_60_1/VGND
flabel locali 497748 363152 497852 363400 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 497177 363240 497226 363341 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 497336 363246 497376 363364 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 497748 364492 497852 364740 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 497177 364580 497226 364681 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 497336 364586 497376 364704 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 497748 365832 497852 366080 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 497177 365920 497226 366021 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 497336 365926 497376 366044 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 497748 367172 497852 367420 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 497177 367260 497226 367361 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 497336 367266 497376 367384 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 497748 368512 497852 368760 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 497177 368600 497226 368701 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 497336 368606 497376 368724 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 497748 369852 497852 370100 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 497177 369940 497226 370041 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 497336 369946 497376 370064 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 497748 371192 497852 371440 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/xm1/Emitter
flabel locali 497177 371280 497226 371381 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/xm1/Collector
flabel locali 497336 371286 497376 371404 0 FreeSans 500 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/xm1/Base
flabel metal1 497608 371214 497738 371454 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/Emitter
flabel metal1 497336 371564 497376 371804 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/Base
flabel metal1 497184 371728 497224 371968 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/Collector
flabel metal1 496838 371934 496898 371994 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/VPWR
flabel metal1 498718 371934 498778 371994 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pnp_05v5_W3p40L3p40_7_0/VGND
flabel metal2 493338 401390 493418 401590 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_9/Cin
flabel metal4 494748 401408 494848 401568 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_9/Cout
flabel metal1 493078 401528 493138 401588 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_9/VPWR
flabel metal1 494958 401528 495018 401588 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_9/VGND
flabel metal2 493338 408838 493418 409038 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_8/Cin
flabel metal4 494748 408856 494848 409016 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_8/Cout
flabel metal1 493078 408976 493138 409036 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_8/VPWR
flabel metal1 494958 408976 495018 409036 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_8/VGND
flabel metal1 493568 393882 493688 394002 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_30/Rin
flabel metal1 494528 393882 494648 394002 7 FreeSans 600 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_30/Rout
flabel metal1 493078 394062 493138 394122 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_30/VPWR
flabel metal1 494958 394062 495018 394122 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_30/VGND
flabel locali 494784 390520 494844 390580 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE
flabel locali 493238 390520 493298 390580 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/SOURCE
flabel locali 494558 390520 494618 390580 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/DRAIN
flabel metal1 493078 390976 493138 391036 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/VPWR
flabel metal1 494958 390976 495018 391036 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/VGND
flabel locali 494824 362516 494884 362576 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_60_2/GATE
flabel locali 493258 362516 493298 362576 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_60_2/SOURCE
flabel locali 494718 362516 494778 362576 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_60_2/DRAIN
flabel nwell 493078 390162 493138 390222 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_60_2/VPWR
flabel metal1 494958 390064 495018 390222 7 FreeSans 1000 0 0 0 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_60_2/VGND
flabel metal2 541962 389410 542060 389438 7 FreeSans 8000 0 0 0 bgr_top_flat_0/porst
flabel metal2 541962 380578 542060 380606 7 FreeSans 8000 0 0 0 bgr_top_flat_0/vbg
flabel metal1 508622 356438 508658 356562 7 FreeSans 8000 0 0 0 bgr_top_flat_0/vb
flabel metal3 501026 414786 501086 414954 7 FreeSans 8000 0 0 0 bgr_top_flat_0/va
flabel metal1 565806 493790 565866 493850 1 FreeSans 800 0 0 0 nmos_flat_0/VPWR
flabel metal1 565806 491910 565866 491970 1 FreeSans 800 0 0 0 nmos_flat_0/VGND
flabel locali 560650 493630 560710 493690 1 FreeSans 800 0 0 0 nmos_flat_0/SOURCE
flabel locali 560650 492310 560710 492370 1 FreeSans 800 0 0 0 nmos_flat_0/DRAIN
flabel locali 560650 492144 560710 492204 1 FreeSans 800 0 0 0 nmos_flat_0/GATE
flabel metal1 560690 404648 560750 404708 1 FreeSans 800 0 0 0 nmos_flat_1/VPWR
flabel metal1 560690 402768 560750 402828 1 FreeSans 800 0 0 0 nmos_flat_1/VGND
flabel locali 565846 404488 565906 404548 1 FreeSans 800 0 0 0 nmos_flat_1/SOURCE
flabel locali 565846 403168 565906 403228 1 FreeSans 800 0 0 0 nmos_flat_1/DRAIN
flabel locali 565846 403002 565906 403062 1 FreeSans 800 0 0 0 nmos_flat_1/GATE
flabel metal1 565698 359330 565758 359390 1 FreeSans 800 0 0 0 nmos_flat_2/VPWR
flabel metal1 565698 357450 565758 357510 1 FreeSans 800 0 0 0 nmos_flat_2/VGND
flabel locali 560542 359170 560602 359230 1 FreeSans 800 0 0 0 nmos_flat_2/SOURCE
flabel locali 560542 357850 560602 357910 1 FreeSans 800 0 0 0 nmos_flat_2/DRAIN
flabel locali 560542 357684 560602 357744 1 FreeSans 800 0 0 0 nmos_flat_2/GATE
flabel nwell 579774 404688 579834 404748 1 FreeSans 800 0 0 0 pmos_flat_0/VPWR
flabel metal1 579676 402808 579834 402868 1 FreeSans 800 0 0 0 pmos_flat_0/VGND
flabel locali 574448 404528 574508 404568 1 FreeSans 800 0 0 0 pmos_flat_0/SOURCE
flabel locali 574448 403148 574508 403208 1 FreeSans 800 0 0 0 pmos_flat_0/DRAIN
flabel locali 574448 402986 574508 403046 1 FreeSans 800 0 0 0 pmos_flat_0/GATE
flabel nwell 579970 359260 580030 359320 1 FreeSans 800 0 0 0 pmos_flat_1/VPWR
flabel metal1 579872 357380 580030 357440 1 FreeSans 800 0 0 0 pmos_flat_1/VGND
flabel locali 574644 359100 574704 359140 1 FreeSans 800 0 0 0 pmos_flat_1/SOURCE
flabel locali 574644 357720 574704 357780 1 FreeSans 800 0 0 0 pmos_flat_1/DRAIN
flabel locali 574644 357558 574704 357618 1 FreeSans 800 0 0 0 pmos_flat_1/GATE
flabel nwell 580496 493564 580556 493624 1 FreeSans 800 0 0 0 pmos_flat_3/VPWR
flabel metal1 580398 491684 580556 491744 1 FreeSans 800 0 0 0 pmos_flat_3/VGND
flabel locali 575170 493404 575230 493444 1 FreeSans 800 0 0 0 pmos_flat_3/SOURCE
flabel locali 575170 492024 575230 492084 1 FreeSans 800 0 0 0 pmos_flat_3/DRAIN
flabel locali 575170 491862 575230 491922 1 FreeSans 800 0 0 0 pmos_flat_3/GATE
<< end >>
