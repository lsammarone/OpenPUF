* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_1 Y A VGND VPWR VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_1 Y B A VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 X A VGND VPWR VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_8 Y A VGND VPWR VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 Q RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_8 A X VGND VPWR VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_1 B Y A VGND VPWR VNB VPB a_109_297#
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 X A VGND VPWR VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VNB VPB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_6 Y A VPWR VGND VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_16 Y A VGND VPWR VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_4 Y A VPWR VGND VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_1#0 a_150_47# w_n38_261# a_68_47# a_68_297# w_42_21#
+ a_64_199# VSUBS
X0 a_150_47# a_64_199# a_68_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_150_47# a_64_199# a_68_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_hvt_UUWA33 a_n73_n100# a_15_n100# w_n109_n200# a_n33_n197#
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n109_n200# sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_PX9ZJG a_63_n65# a_n125_n65# a_15_87# a_n81_n153#
+ a_n33_n65# w_n151_n91# VSUBS
X0 a_n33_n65# a_n81_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_63_n65# a_15_87# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_hvt_SH6FHF w_n161_n200# a_n125_n100# a_63_n100# a_15_131#
+ a_n33_n100# a_n81_n197#
X0 a_63_n100# a_15_131# a_n33_n100# w_n161_n200# sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n33_n100# a_n81_n197# a_n125_n100# w_n161_n200# sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt mux 2/VSUBS w_n54_614# w_18_n122# m1_46_n2# m1_76_558# m1_188_418# m1_n50_88#
+ a_28_318# sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# VSUBS
X1 m1_188_418# m1_n50_88# a_28_318# m1_46_n2# m1_76_558# 1/w_n151_n91# 2/VSUBS sky130_fd_pr__nfet_01v8_PX9ZJG
X2 w_n54_614# m1_n50_88# m1_188_418# m1_46_n2# m1_76_558# a_28_318# sky130_fd_pr__pfet_01v8_hvt_SH6FHF
Xsky130_fd_pr__nfet_01v8_PX9ZJG_0 m1_188_418# m1_n50_88# a_28_318# m1_46_n2# m1_76_558#
+ sky130_fd_pr__nfet_01v8_PX9ZJG_0/w_n151_n91# 2/VSUBS sky130_fd_pr__nfet_01v8_PX9ZJG
Xsky130_fd_pr__nfet_01v8_PX9ZJG_1 m1_188_418# m1_n50_88# a_28_318# m1_46_n2# m1_76_558#
+ sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# 2/VSUBS sky130_fd_pr__nfet_01v8_PX9ZJG
Xsky130_fd_pr__pfet_01v8_hvt_SH6FHF_0 w_n54_614# m1_n50_88# m1_188_418# m1_46_n2#
+ m1_76_558# a_28_318# sky130_fd_pr__pfet_01v8_hvt_SH6FHF
Xsky130_fd_pr__pfet_01v8_hvt_SH6FHF_1 w_n54_614# m1_n50_88# m1_188_418# m1_46_n2#
+ m1_76_558# a_28_318# sky130_fd_pr__pfet_01v8_hvt_SH6FHF
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VNB VPB a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt demux m1_188_418# 2/VSUBS w_n54_614# w_18_n122# m1_46_n2# m1_76_558# a_28_318#
+ 1/w_n151_n91# m1_n50_88# VSUBS
X1 m1_188_418# m1_n50_88# a_28_318# m1_46_n2# m1_76_558# 1/w_n151_n91# 2/VSUBS sky130_fd_pr__nfet_01v8_PX9ZJG
X2 w_n54_614# m1_n50_88# m1_188_418# m1_46_n2# m1_76_558# a_28_318# sky130_fd_pr__pfet_01v8_hvt_SH6FHF
Xsky130_fd_pr__nfet_01v8_PX9ZJG_0 m1_188_418# m1_n50_88# a_28_318# m1_46_n2# m1_76_558#
+ 1/w_n151_n91# 2/VSUBS sky130_fd_pr__nfet_01v8_PX9ZJG
Xsky130_fd_pr__nfet_01v8_PX9ZJG_1 m1_188_418# m1_n50_88# a_28_318# m1_46_n2# m1_76_558#
+ 1/w_n151_n91# 2/VSUBS sky130_fd_pr__nfet_01v8_PX9ZJG
Xsky130_fd_pr__pfet_01v8_hvt_SH6FHF_0 w_n54_614# m1_n50_88# m1_188_418# m1_46_n2#
+ m1_76_558# a_28_318# sky130_fd_pr__pfet_01v8_hvt_SH6FHF
Xsky130_fd_pr__pfet_01v8_hvt_SH6FHF_1 w_n54_614# m1_n50_88# m1_188_418# m1_46_n2#
+ m1_76_558# a_28_318# sky130_fd_pr__pfet_01v8_hvt_SH6FHF
.ends

.subckt unitcell2buf sky130_fd_sc_hd__nor2_1_3/a_109_297# sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ sky130_fd_sc_hd__nor2_1_2/a_109_297# demux_0/w_18_n122# demux_0/1/w_n151_n91# sky130_fd_sc_hd__buf_1_1/X
+ li_n460_n386# sky130_fd_sc_hd__buf_1_1/a_27_47# mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__nor2_1_2/B li_80_172# sky130_fd_sc_hd__nor2_1_3/Y
+ m2_136_462# sky130_fd_sc_hd__buf_1_1/VPB mux_0/w_18_n122# sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__nor2_1_3/A a_24_n198# sky130_fd_sc_hd__nor2_1_2/Y sky130_fd_sc_hd__nor2_1_3/B
+ VSUBS
Xsky130_fd_sc_hd__inv_1#0_0 li_80_172# sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__inv_1#0_0/w_42_21# a_24_n198# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1#0_1 a_24_n198# sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__inv_1#0_1/w_42_21# li_n460_n386# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__nor2_1_3/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__nor2_1_3/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__nor2_1_2/Y
+ sky130_fd_sc_hd__nor2_1_3/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__nor2_1_2/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_2 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__nor2_1_2/Y
+ sky130_fd_sc_hd__nor2_1_3/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__nor2_1_2/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_3 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__nor2_1_3/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__nor2_1_3/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_pr__pfet_01v8_hvt_UUWA33_0 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__buf_1_1/VPB li_80_172# sky130_fd_pr__pfet_01v8_hvt_UUWA33
X1 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/VPB
+ li_80_172# sky130_fd_pr__pfet_01v8_hvt_UUWA33
Xsky130_fd_pr__pfet_01v8_hvt_UUWA33_1 sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__buf_1_1/VPB a_24_n198# sky130_fd_pr__pfet_01v8_hvt_UUWA33
X2 sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__buf_1_1/VPB
+ a_24_n198# sky130_fd_pr__pfet_01v8_hvt_UUWA33
Xmux_0 VSUBS sky130_fd_sc_hd__buf_1_1/VPB mux_0/w_18_n122# li_80_172# sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__nor2_1_2/Y a_24_n198# mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ mux_0/VSUBS mux
Xmux_1 VSUBS sky130_fd_sc_hd__buf_1_1/VPB mux_1/w_18_n122# li_80_172# sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__nor2_1_2/Y a_24_n198# mux_1/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ mux_1/VSUBS mux
Xsky130_fd_sc_hd__buf_1_0 VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/X
+ sky130_fd_sc_hd__buf_1_1/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__buf_1_1 VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/X
+ sky130_fd_sc_hd__buf_1_1/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__inv_1_0 li_80_172# sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__inv_1_0/w_42_21# a_24_n198# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1_1 a_24_n198# sky130_fd_sc_hd__buf_1_1/VPB VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__inv_1_1/w_42_21# li_n460_n386# VSUBS sky130_fd_sc_hd__inv_1#0
Xdemux_0 sky130_fd_sc_hd__nor2_1_3/B VSUBS sky130_fd_sc_hd__buf_1_1/VPB demux_0/w_18_n122#
+ li_80_172# m2_136_462# a_24_n198# demux_0/1/w_n151_n91# sky130_fd_sc_hd__nor2_1_2/B
+ demux_0/VSUBS demux
Xdemux_1 sky130_fd_sc_hd__nor2_1_3/B VSUBS sky130_fd_sc_hd__buf_1_1/VPB demux_1/w_18_n122#
+ li_80_172# m2_136_462# a_24_n198# demux_1/1/w_n151_n91# sky130_fd_sc_hd__nor2_1_2/B
+ demux_1/VSUBS demux
.ends

.subckt unitcell2bufcut sky130_fd_sc_hd__nor2_1_3/a_109_297# sky130_fd_sc_hd__inv_1_1/w_42_21#
+ sky130_fd_sc_hd__nor2_1_2/a_109_297# sky130_fd_sc_hd__nor2_1_2/B demux_1/1/w_n151_n91#
+ a_24_n198# li_n460_n386# sky130_fd_sc_hd__buf_1_1/a_27_47# mux_1/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ li_80_172# sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__nor2_1_2/Y m2_136_462# sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/X sky130_fd_sc_hd__inv_1_0/w_42_21#
+ sky130_fd_sc_hd__nor2_1_3/A sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__buf_1_1/VGND
+ VSUBS
Xsky130_fd_sc_hd__inv_1#0_0 li_80_172# sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/VGND
+ sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__inv_1_0/w_42_21# a_24_n198# VSUBS
+ sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1#0_1 a_24_n198# sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/VGND
+ sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__inv_1_1/w_42_21# li_n460_n386# VSUBS
+ sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__nor2_1_3/A sky130_fd_sc_hd__buf_1_1/VGND sky130_fd_sc_hd__buf_1_1/VPB
+ VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_3/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__nor2_1_2/Y
+ sky130_fd_sc_hd__nor2_1_3/A sky130_fd_sc_hd__buf_1_1/VGND sky130_fd_sc_hd__buf_1_1/VPB
+ VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_2/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_2 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__nor2_1_2/Y
+ sky130_fd_sc_hd__nor2_1_3/A sky130_fd_sc_hd__buf_1_1/VGND sky130_fd_sc_hd__buf_1_1/VPB
+ VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_2/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_3 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__nor2_1_3/A sky130_fd_sc_hd__buf_1_1/VGND sky130_fd_sc_hd__buf_1_1/VPB
+ VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_3/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_pr__pfet_01v8_hvt_UUWA33_0 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__buf_1_1/VPB li_80_172# sky130_fd_pr__pfet_01v8_hvt_UUWA33
X1 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/VPB
+ li_80_172# sky130_fd_pr__pfet_01v8_hvt_UUWA33
Xsky130_fd_pr__pfet_01v8_hvt_UUWA33_1 sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__buf_1_1/VPB a_24_n198# sky130_fd_pr__pfet_01v8_hvt_UUWA33
X2 sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__buf_1_1/VPB
+ a_24_n198# sky130_fd_pr__pfet_01v8_hvt_UUWA33
Xmux_0 mux_0/2/VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/VGND li_80_172#
+ sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__nor2_1_2/Y
+ a_24_n198# mux_1/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# VSUBS mux
Xmux_1 mux_1/2/VSUBS sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/VGND li_80_172#
+ sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__nor2_1_2/Y
+ a_24_n198# mux_1/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# VSUBS mux
Xsky130_fd_sc_hd__buf_1_0 sky130_fd_sc_hd__buf_1_1/VGND sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__buf_1_1/X sky130_fd_sc_hd__buf_1_1/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__buf_1_1/a_27_47# sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__buf_1_1 sky130_fd_sc_hd__buf_1_1/VGND sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__buf_1_1/X sky130_fd_sc_hd__buf_1_1/A VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__buf_1_1/a_27_47# sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__inv_1_0 li_80_172# sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/VGND
+ sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__inv_1_0/w_42_21# a_24_n198# VSUBS
+ sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1_1 a_24_n198# sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__buf_1_1/VGND
+ sky130_fd_sc_hd__buf_1_1/VPB sky130_fd_sc_hd__inv_1_1/w_42_21# li_n460_n386# VSUBS
+ sky130_fd_sc_hd__inv_1#0
Xdemux_0 sky130_fd_sc_hd__nor2_1_3/B demux_0/2/VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__buf_1_1/VGND li_80_172# m2_136_462# a_24_n198# demux_1/1/w_n151_n91#
+ sky130_fd_sc_hd__nor2_1_2/B VSUBS demux
Xdemux_1 sky130_fd_sc_hd__nor2_1_3/B demux_1/2/VSUBS sky130_fd_sc_hd__buf_1_1/VPB
+ sky130_fd_sc_hd__buf_1_1/VGND li_80_172# m2_136_462# a_24_n198# demux_1/1/w_n151_n91#
+ sky130_fd_sc_hd__nor2_1_2/B VSUBS demux
.ends

.subckt brbufhalf unitcell2buf_7/li_n460_n386# unitcell2bufcut_3/li_n460_n386# sky130_fd_sc_hd__inv_16_7/A
+ unitcell2buf_2/li_n460_n386# unitcell2buf_24/li_n460_n386# sky130_fd_sc_hd__inv_16_6/VGND
+ unitcell2buf_5/li_n460_n386# unitcell2buf_27/li_n460_n386# unitcell2buf_8/li_n460_n386#
+ unitcell2buf_0/li_n460_n386# unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_7/VGND unitcell2buf_25/li_n460_n386# unitcell2bufcut_2/li_n460_n386#
+ unitcell2buf_6/li_n460_n386# sky130_fd_sc_hd__inv_16_4/VGND unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_9/li_n460_n386# unitcell2buf_1/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_5/A
+ unitcell2buf_26/m2_136_462# sky130_fd_sc_hd__inv_16_5/VGND VSUBS unitcell2buf_26/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_7/VPB
Xunitcell2buf_1 unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_1/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_1/demux_0/w_18_n122#
+ unitcell2buf_1/demux_0/1/w_n151_n91# unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_1/li_n460_n386#
+ unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_1/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_1/li_80_172# unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_1/mux_0/w_18_n122# unitcell2buf_1/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_1/a_24_n198# unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/A
+ sky130_fd_sc_hd__inv_16_7/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_2 unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_2/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_2/demux_0/w_18_n122#
+ unitcell2buf_2/demux_0/1/w_n151_n91# unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_2/li_n460_n386#
+ unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_2/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_2/li_80_172# unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_2/mux_0/w_18_n122# unitcell2buf_2/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_2/a_24_n198# unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_4 sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_5/A
+ sky130_fd_sc_hd__inv_16_4/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_5 sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_5/A
+ sky130_fd_sc_hd__inv_16_5/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_3 unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_3/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_3/demux_0/w_18_n122#
+ unitcell2buf_3/demux_0/1/w_n151_n91# unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_3/li_n460_n386#
+ unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_3/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_3/li_80_172# unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_3/mux_0/w_18_n122# unitcell2buf_3/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_3/a_24_n198# unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_6 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/A
+ sky130_fd_sc_hd__inv_16_6/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_4 unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_4/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_4/demux_0/w_18_n122#
+ unitcell2buf_4/demux_0/1/w_n151_n91# unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_4/li_n460_n386#
+ unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_4/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_4/li_80_172# unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB VSUBS unitcell2buf_4/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_4/a_24_n198# unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_7 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/A
+ sky130_fd_sc_hd__inv_16_7/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_5 unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_5/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_5/demux_0/w_18_n122#
+ unitcell2buf_5/demux_0/1/w_n151_n91# unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_5/li_n460_n386#
+ unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_5/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_5/li_80_172# unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_5/mux_0/w_18_n122# unitcell2buf_5/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_5/a_24_n198# unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_6 unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_6/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_6/demux_0/w_18_n122#
+ unitcell2buf_6/demux_0/1/w_n151_n91# unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_6/li_n460_n386#
+ unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_6/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_6/li_80_172# unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/Y unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_6/mux_0/w_18_n122# unitcell2buf_6/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_6/a_24_n198# unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_7 unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_7/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_7/demux_0/w_18_n122#
+ unitcell2buf_7/demux_0/1/w_n151_n91# unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_7/li_n460_n386#
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_7/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_7/li_80_172# unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_7/mux_0/w_18_n122# unitcell2buf_7/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_7/a_24_n198# unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_8 unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_8/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_8/demux_0/w_18_n122#
+ unitcell2buf_8/demux_0/1/w_n151_n91# unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_8/li_n460_n386#
+ unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_8/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_8/li_80_172# unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_8/mux_0/w_18_n122# unitcell2buf_8/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_8/a_24_n198# unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_9 unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_9/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_9/demux_0/w_18_n122#
+ unitcell2buf_9/demux_0/1/w_n151_n91# unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_9/li_n460_n386#
+ unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_9/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_9/li_80_172# unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_9/mux_0/w_18_n122# unitcell2buf_9/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_9/a_24_n198# unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_20 unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_6/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_6/demux_0/w_18_n122#
+ unitcell2buf_6/demux_0/1/w_n151_n91# unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_6/li_n460_n386#
+ unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_6/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_6/li_80_172# unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/Y unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_20/mux_0/w_18_n122# unitcell2buf_6/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_6/a_24_n198# unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_21 unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_7/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_7/demux_0/w_18_n122#
+ unitcell2buf_7/demux_0/1/w_n151_n91# unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_7/li_n460_n386#
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_7/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_7/li_80_172# unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB VSUBS unitcell2buf_7/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_7/a_24_n198# unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_22 unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_8/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_8/demux_0/w_18_n122#
+ unitcell2buf_8/demux_0/1/w_n151_n91# unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_8/li_n460_n386#
+ unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_8/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_8/li_80_172# unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_22/mux_0/w_18_n122# unitcell2buf_8/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_8/a_24_n198# unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_10 unitcell2buf_24/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_24/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_24/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_24/demux_0/w_18_n122#
+ unitcell2buf_24/demux_0/1/w_n151_n91# unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/X
+ unitcell2buf_24/li_n460_n386# unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_24/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_24/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_24/li_80_172# unitcell2buf_24/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_10/mux_0/w_18_n122#
+ unitcell2buf_24/sky130_fd_sc_hd__inv_1#0_0/w_42_21# sky130_fd_sc_hd__inv_16_7/Y
+ unitcell2buf_24/a_24_n198# unitcell2buf_24/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_24/sky130_fd_sc_hd__nor2_1_3/B
+ VSUBS unitcell2buf
Xunitcell2buf_11 unitcell2buf_25/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_25/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_25/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_25/demux_0/w_18_n122#
+ unitcell2buf_25/demux_0/1/w_n151_n91# unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/X
+ unitcell2buf_25/li_n460_n386# unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_25/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_25/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_25/li_80_172# unitcell2buf_25/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_11/mux_0/w_18_n122#
+ unitcell2buf_25/sky130_fd_sc_hd__inv_1#0_0/w_42_21# sky130_fd_sc_hd__inv_16_7/Y
+ unitcell2buf_25/a_24_n198# unitcell2buf_25/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_25/sky130_fd_sc_hd__nor2_1_3/B
+ VSUBS unitcell2buf
Xunitcell2buf_23 unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_9/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_9/demux_0/w_18_n122#
+ unitcell2buf_9/demux_0/1/w_n151_n91# unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_9/li_n460_n386#
+ unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_9/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_9/li_80_172# unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB VSUBS unitcell2buf_9/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_9/a_24_n198# unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_12 unitcell2buf_26/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_26/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_26/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_26/demux_0/w_18_n122#
+ unitcell2buf_26/demux_0/1/w_n151_n91# unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/X
+ unitcell2buf_26/li_n460_n386# unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_26/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_26/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_26/li_80_172# unitcell2buf_26/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2buf_26/m2_136_462# sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_26/mux_0/w_18_n122#
+ unitcell2buf_26/sky130_fd_sc_hd__inv_1#0_0/w_42_21# sky130_fd_sc_hd__inv_16_7/Y
+ unitcell2buf_26/a_24_n198# unitcell2buf_26/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_26/sky130_fd_sc_hd__nor2_1_3/B
+ VSUBS unitcell2buf
Xunitcell2buf_24 unitcell2buf_24/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_24/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_24/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_24/demux_0/w_18_n122#
+ unitcell2buf_24/demux_0/1/w_n151_n91# unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/X
+ unitcell2buf_24/li_n460_n386# unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_24/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_24/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_24/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_24/li_80_172# unitcell2buf_24/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB VSUBS unitcell2buf_24/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_24/a_24_n198# unitcell2buf_24/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_24/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_13 unitcell2buf_27/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_27/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_27/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_27/demux_0/w_18_n122#
+ unitcell2buf_27/demux_0/1/w_n151_n91# unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/X
+ unitcell2buf_27/li_n460_n386# unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_27/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_27/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_27/li_80_172# unitcell2buf_27/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_13/mux_0/w_18_n122#
+ unitcell2buf_27/sky130_fd_sc_hd__inv_1#0_0/w_42_21# sky130_fd_sc_hd__inv_16_7/Y
+ unitcell2buf_27/a_24_n198# unitcell2buf_27/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_27/sky130_fd_sc_hd__nor2_1_3/B
+ VSUBS unitcell2buf
Xunitcell2buf_14 unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_0/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_0/demux_0/w_18_n122#
+ unitcell2buf_0/demux_0/1/w_n151_n91# unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_0/li_n460_n386#
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_0/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_0/li_80_172# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_0/mux_0/w_18_n122# unitcell2buf_0/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_0/a_24_n198# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_25 unitcell2buf_25/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_25/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_25/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_25/demux_0/w_18_n122#
+ unitcell2buf_25/demux_0/1/w_n151_n91# unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/X
+ unitcell2buf_25/li_n460_n386# unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_25/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_25/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_25/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_25/li_80_172# unitcell2buf_25/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_25/mux_0/w_18_n122#
+ unitcell2buf_25/sky130_fd_sc_hd__inv_1#0_0/w_42_21# sky130_fd_sc_hd__inv_16_7/Y
+ unitcell2buf_25/a_24_n198# unitcell2buf_25/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_25/sky130_fd_sc_hd__nor2_1_3/B
+ VSUBS unitcell2buf
Xunitcell2buf_15 unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_1/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_1/demux_0/w_18_n122#
+ unitcell2buf_1/demux_0/1/w_n151_n91# unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_1/li_n460_n386#
+ unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_1/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_1/li_80_172# unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_1/mux_0/w_18_n122# unitcell2buf_1/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_1/a_24_n198# unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_26 unitcell2buf_26/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_26/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_26/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_26/demux_0/w_18_n122#
+ unitcell2buf_26/demux_0/1/w_n151_n91# unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/X
+ unitcell2buf_26/li_n460_n386# unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_26/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_26/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_26/li_80_172# unitcell2buf_26/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2buf_26/m2_136_462# sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_26/mux_0/w_18_n122#
+ unitcell2buf_26/sky130_fd_sc_hd__inv_1#0_0/w_42_21# sky130_fd_sc_hd__inv_16_7/Y
+ unitcell2buf_26/a_24_n198# unitcell2buf_26/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_26/sky130_fd_sc_hd__nor2_1_3/B
+ VSUBS unitcell2buf
Xunitcell2buf_16 unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_2/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_2/demux_0/w_18_n122#
+ unitcell2buf_2/demux_0/1/w_n151_n91# unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_2/li_n460_n386#
+ unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_2/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_2/li_80_172# unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB VSUBS unitcell2buf_2/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_2/a_24_n198# unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_27 unitcell2buf_27/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_27/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_27/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_27/demux_0/w_18_n122#
+ unitcell2buf_27/demux_0/1/w_n151_n91# unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/X
+ unitcell2buf_27/li_n460_n386# unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_27/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_27/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_27/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_27/li_80_172# unitcell2buf_27/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2buf_26/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_7/VPB VSUBS unitcell2buf_27/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_27/a_24_n198# unitcell2buf_27/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_27/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_17 unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_3/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_3/demux_0/w_18_n122#
+ unitcell2buf_3/demux_0/1/w_n151_n91# unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_3/li_n460_n386#
+ unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_3/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_3/li_80_172# unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_17/mux_0/w_18_n122# unitcell2buf_3/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_3/a_24_n198# unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_18 unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_4/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_4/demux_0/w_18_n122#
+ unitcell2buf_4/demux_0/1/w_n151_n91# unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_4/li_n460_n386#
+ unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_4/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_4/li_80_172# unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB VSUBS unitcell2buf_4/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_4/a_24_n198# unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_19 unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_5/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_5/demux_0/w_18_n122#
+ unitcell2buf_5/demux_0/1/w_n151_n91# unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_5/li_n460_n386#
+ unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_5/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_5/li_80_172# unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB VSUBS unitcell2buf_5/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_5/a_24_n198# unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2bufcut_0 unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2bufcut_2/sky130_fd_sc_hd__inv_1_1/w_42_21#
+ unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2bufcut_2/demux_1/1/w_n151_n91# unitcell2bufcut_2/a_24_n198# unitcell2bufcut_2/li_n460_n386#
+ unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2bufcut_2/mux_1/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2bufcut_2/li_80_172# unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X unitcell2bufcut_2/sky130_fd_sc_hd__inv_1_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_3/B VSUBS
+ VSUBS unitcell2bufcut
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_5/A
+ sky130_fd_sc_hd__inv_16_4/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2bufcut_1 unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2bufcut_3/sky130_fd_sc_hd__inv_1_1/w_42_21#
+ unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2bufcut_3/demux_1/1/w_n151_n91# unitcell2bufcut_3/a_24_n198# unitcell2bufcut_3/li_n460_n386#
+ unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2bufcut_3/mux_1/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2bufcut_3/li_80_172# unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/X unitcell2bufcut_3/sky130_fd_sc_hd__inv_1_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_7/Y unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_3/B VSUBS
+ VSUBS unitcell2bufcut
Xunitcell2bufcut_2 unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2bufcut_2/sky130_fd_sc_hd__inv_1_1/w_42_21#
+ unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2bufcut_2/demux_1/1/w_n151_n91# unitcell2bufcut_2/a_24_n198# unitcell2bufcut_2/li_n460_n386#
+ unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2bufcut_2/mux_1/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2bufcut_2/li_80_172# unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X unitcell2bufcut_2/sky130_fd_sc_hd__inv_1_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2bufcut_2/sky130_fd_sc_hd__nor2_1_3/B VSUBS
+ VSUBS unitcell2bufcut
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_5/Y sky130_fd_sc_hd__inv_16_5/A
+ sky130_fd_sc_hd__inv_16_5/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_0 unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_0/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_0/demux_0/w_18_n122#
+ unitcell2buf_0/demux_0/1/w_n151_n91# unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_0/li_n460_n386#
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_0/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_0/li_80_172# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2buf_0/mux_0/w_18_n122# unitcell2buf_0/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_5/Y unitcell2buf_0/a_24_n198# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2bufcut_3 unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2bufcut_3/sky130_fd_sc_hd__inv_1_1/w_42_21#
+ unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2bufcut_3/demux_1/1/w_n151_n91# unitcell2bufcut_3/a_24_n198# unitcell2bufcut_3/li_n460_n386#
+ unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2bufcut_3/mux_1/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2bufcut_3/li_80_172# unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__inv_16_7/VPB unitcell2bufcut_3/sky130_fd_sc_hd__buf_1_1/X unitcell2bufcut_3/sky130_fd_sc_hd__inv_1_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_7/Y unitcell2bufcut_3/sky130_fd_sc_hd__nor2_1_3/B VSUBS
+ VSUBS unitcell2bufcut
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/A
+ sky130_fd_sc_hd__inv_16_6/VGND sky130_fd_sc_hd__inv_16_7/VPB VSUBS sky130_fd_sc_hd__inv_16_7/VPB
+ sky130_fd_sc_hd__inv_16
.ends

.subckt brbufhalf_64 unitcell2buf_7/li_n460_n386# unitcell2buf_2/li_n460_n386# unitcell2buf_10/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_2/VGND unitcell2buf_5/li_n460_n386# unitcell2buf_13/li_n460_n386#
+ unitcell2buf_8/li_n460_n386# sky130_fd_sc_hd__inv_16_1/A unitcell2buf_0/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/A unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/VGND unitcell2buf_11/li_n460_n386# sky130_fd_sc_hd__inv_16_0/VGND
+ unitcell2bufcut_0/li_n460_n386# unitcell2buf_6/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ unitcell2buf_9/li_n460_n386# unitcell2buf_1/li_n460_n386# unitcell2buf_4/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_1/VGND unitcell2buf_12/m2_136_462# VSUBS unitcell2buf_12/li_n460_n386#
Xunitcell2buf_1 unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_1/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_1/demux_0/w_18_n122#
+ unitcell2buf_1/demux_0/1/w_n151_n91# unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_1/li_n460_n386#
+ unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_1/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_1/li_80_172# unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_1/mux_0/w_18_n122# unitcell2buf_1/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_1/a_24_n198# unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16_3/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_2 unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_2/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_2/demux_0/w_18_n122#
+ unitcell2buf_2/demux_0/1/w_n151_n91# unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_2/li_n460_n386#
+ unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_2/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_2/li_80_172# unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_2/mux_0/w_18_n122# unitcell2buf_2/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_2/a_24_n198# unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_3 unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_3/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_3/demux_0/w_18_n122#
+ unitcell2buf_3/demux_0/1/w_n151_n91# unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_3/li_n460_n386#
+ unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_3/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_3/li_80_172# unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_3/mux_0/w_18_n122# unitcell2buf_3/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_3/a_24_n198# unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_4 unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_4/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_4/demux_0/w_18_n122#
+ unitcell2buf_4/demux_0/1/w_n151_n91# unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_4/li_n460_n386#
+ unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_4/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_4/li_80_172# unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_4/mux_0/w_18_n122# unitcell2buf_4/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_4/a_24_n198# unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_5 unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_5/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_5/demux_0/w_18_n122#
+ unitcell2buf_5/demux_0/1/w_n151_n91# unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_5/li_n460_n386#
+ unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_5/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_5/li_80_172# unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_5/mux_0/w_18_n122# unitcell2buf_5/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_5/a_24_n198# unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_6 unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_6/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_6/demux_0/w_18_n122#
+ unitcell2buf_6/demux_0/1/w_n151_n91# unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_6/li_n460_n386#
+ unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_6/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_6/li_80_172# unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/Y unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_6/mux_0/w_18_n122# unitcell2buf_6/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_6/a_24_n198# unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_7 unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_7/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_7/demux_0/w_18_n122#
+ unitcell2buf_7/demux_0/1/w_n151_n91# unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_7/li_n460_n386#
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_7/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_7/li_80_172# unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_7/mux_0/w_18_n122# unitcell2buf_7/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_7/a_24_n198# unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_8 unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_8/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_8/demux_0/w_18_n122#
+ unitcell2buf_8/demux_0/1/w_n151_n91# unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_8/li_n460_n386#
+ unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_8/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_8/li_80_172# unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_8/mux_0/w_18_n122# unitcell2buf_8/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_8/a_24_n198# unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_9 unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_9/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_9/demux_0/w_18_n122#
+ unitcell2buf_9/demux_0/1/w_n151_n91# unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_9/li_n460_n386#
+ unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_9/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_9/li_80_172# unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_9/mux_0/w_18_n122# unitcell2buf_9/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_9/a_24_n198# unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_10 unitcell2buf_10/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_10/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_10/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_10/demux_0/w_18_n122#
+ unitcell2buf_10/demux_0/1/w_n151_n91# unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/X
+ unitcell2buf_10/li_n460_n386# unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_10/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_10/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_10/li_80_172# unitcell2buf_10/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_10/mux_0/w_18_n122#
+ unitcell2buf_10/sky130_fd_sc_hd__inv_1#0_0/w_42_21# sky130_fd_sc_hd__inv_16_3/Y
+ unitcell2buf_10/a_24_n198# unitcell2buf_10/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_10/sky130_fd_sc_hd__nor2_1_3/B
+ VSUBS unitcell2buf
Xunitcell2buf_11 unitcell2buf_11/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_11/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_11/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_11/demux_0/w_18_n122#
+ unitcell2buf_11/demux_0/1/w_n151_n91# unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/X
+ unitcell2buf_11/li_n460_n386# unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_11/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_11/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_11/li_80_172# unitcell2buf_11/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2buf_13/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_11/mux_0/w_18_n122#
+ unitcell2buf_11/sky130_fd_sc_hd__inv_1#0_0/w_42_21# sky130_fd_sc_hd__inv_16_3/Y
+ unitcell2buf_11/a_24_n198# unitcell2buf_11/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_11/sky130_fd_sc_hd__nor2_1_3/B
+ VSUBS unitcell2buf
Xunitcell2buf_12 unitcell2buf_12/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_12/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_12/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_12/demux_0/w_18_n122#
+ unitcell2buf_12/demux_0/1/w_n151_n91# unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/X
+ unitcell2buf_12/li_n460_n386# unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_12/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_12/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_12/li_80_172# unitcell2buf_12/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2buf_12/m2_136_462# sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_12/mux_0/w_18_n122#
+ unitcell2buf_12/sky130_fd_sc_hd__inv_1#0_0/w_42_21# sky130_fd_sc_hd__inv_16_3/Y
+ unitcell2buf_12/a_24_n198# unitcell2buf_12/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_12/sky130_fd_sc_hd__nor2_1_3/B
+ VSUBS unitcell2buf
Xunitcell2buf_13 unitcell2buf_13/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_13/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_13/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_13/demux_0/w_18_n122#
+ unitcell2buf_13/demux_0/1/w_n151_n91# unitcell2buf_13/sky130_fd_sc_hd__buf_1_1/X
+ unitcell2buf_13/li_n460_n386# unitcell2buf_13/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_13/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_13/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_13/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_13/li_80_172# unitcell2buf_13/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_13/mux_0/w_18_n122#
+ unitcell2buf_13/sky130_fd_sc_hd__inv_1#0_0/w_42_21# sky130_fd_sc_hd__inv_16_3/Y
+ unitcell2buf_13/a_24_n198# unitcell2buf_13/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_13/sky130_fd_sc_hd__nor2_1_3/B
+ VSUBS unitcell2buf
Xunitcell2bufcut_0 unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2bufcut_0/sky130_fd_sc_hd__inv_1_1/w_42_21#
+ unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2bufcut_0/demux_1/1/w_n151_n91# unitcell2bufcut_0/a_24_n198# unitcell2bufcut_0/li_n460_n386#
+ unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2bufcut_0/mux_1/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2bufcut_0/li_80_172# unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/X unitcell2bufcut_0/sky130_fd_sc_hd__inv_1_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_3/Y unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_3/B VSUBS
+ VSUBS unitcell2bufcut
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_0/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_1/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_0 unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_0/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_0/demux_0/w_18_n122#
+ unitcell2buf_0/demux_0/1/w_n151_n91# unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_0/li_n460_n386#
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_0/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_0/li_80_172# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_0/mux_0/w_18_n122# unitcell2buf_0/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_0/a_24_n198# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16_2/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
.ends

.subckt BR64 OUT VDD RESET C[0] C[1] C[2] C[3] C[4] C[5] C[6] C[7] C[8] C[9] C[10]
+ C[11] C[12] C[13] C[14] C[15] C[16] C[17] C[18] C[19] C[20] C[21] C[22] C[23] C[24]
+ C[25] C[26] C[27] C[28] C[29] C[30] C[31] C[32] C[33] C[34] C[35] C[36] C[37] C[38]
+ C[39] C[40] C[41] C[42] C[43] C[44] C[45] C[46] C[47] C[48] C[49] C[50] C[51] C[52]
+ C[53] C[54] C[55] C[56] C[57] C[58] C[59] C[60] C[61] C[62] C[63] VSS
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__inv_16_4/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_4 sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__inv_16_4/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_4_0 sky130_fd_sc_hd__inv_4_0/Y RESET VDD VSS VSS VDD sky130_fd_sc_hd__inv_4
Xbrbufhalf_0 C[6] C[7] sky130_fd_sc_hd__inv_16_1/Y C[12] C[3] VSS C[9] C[1] C[5] C[14]
+ brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X C[11] VSS C[2] C[15] C[8]
+ VSS brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A brbufhalf_0/sky130_fd_sc_hd__inv_16_7/Y
+ C[4] C[13] brbufhalf_0/sky130_fd_sc_hd__inv_16_5/Y C[10] sky130_fd_sc_hd__inv_16_1/Y
+ brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A VSS VSS C[0] VDD brbufhalf
Xbrbufhalf_1 C[54] C[55] sky130_fd_sc_hd__inv_16_1/Y C[60] C[51] VSS C[57] C[49] C[53]
+ C[62] OUT C[59] VSS C[50] C[63] C[56] VSS brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_1/sky130_fd_sc_hd__inv_16_7/Y C[52] C[61] brbufhalf_1/sky130_fd_sc_hd__inv_16_5/Y
+ C[58] sky130_fd_sc_hd__inv_16_1/Y brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ VSS VSS C[48] VDD brbufhalf
Xbrbufhalf_2 C[38] C[39] sky130_fd_sc_hd__inv_16_4/Y C[44] C[35] VSS C[41] C[33] C[37]
+ C[46] brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X C[43] VSS C[34] C[47]
+ C[40] VSS brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A brbufhalf_2/sky130_fd_sc_hd__inv_16_7/Y
+ C[36] C[45] brbufhalf_2/sky130_fd_sc_hd__inv_16_5/Y C[42] sky130_fd_sc_hd__inv_16_4/Y
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A VSS VSS C[32] VDD brbufhalf
Xbrbufhalf_64_0 C[22] C[28] C[19] VSS C[25] C[17] C[21] sky130_fd_sc_hd__inv_16_4/Y
+ C[30] sky130_fd_sc_hd__inv_16_4/Y brbufhalf_64_0/unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ C[27] VSS C[18] VSS C[23] C[24] VDD C[20] C[29] C[26] VSS brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ VSS C[16] brbufhalf_64
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_4/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_4/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_4_0/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xunitcell2buf_0 unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_0/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_0/demux_0/w_18_n122#
+ unitcell2buf_0/demux_0/1/w_n151_n91# unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/X C[31]
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_0/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_0/li_80_172# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/Y brbufhalf_64_0/unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ VDD unitcell2buf_0/mux_0/w_18_n122# unitcell2buf_0/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ brbufhalf_2/sky130_fd_sc_hd__inv_16_7/Y unitcell2buf_0/a_24_n198# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/B VSS unitcell2buf
.ends

.subckt sky130_fd_sc_hd__nand2_2 Y A B VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt unitcell2bufcut_32 IN C VDD OUT buf_out sky130_fd_sc_hd__nor2_1_1/A VSS VSUBS
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_1_0/B sky130_fd_sc_hd__nor2_1_0/Y
+ sky130_fd_sc_hd__nor2_1_1/A VSS VDD VSUBS VDD sky130_fd_sc_hd__nor2_1_0/a_109_297#
+ sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_1/B sky130_fd_sc_hd__nor2_1_1/Y
+ sky130_fd_sc_hd__nor2_1_1/A VSS VDD VSUBS VDD sky130_fd_sc_hd__nor2_1_1/a_109_297#
+ sky130_fd_sc_hd__nor2_1
X1 sky130_fd_sc_hd__nor2_1_0/B VDD VDD li_80_172# sky130_fd_pr__pfet_01v8_hvt_UUWA33
X2 VDD sky130_fd_sc_hd__nor2_1_1/B VDD a_24_n198# sky130_fd_pr__pfet_01v8_hvt_UUWA33
Xmux_0 mux_0/2/VSUBS VDD VSS li_80_172# OUT sky130_fd_sc_hd__nor2_1_1/Y sky130_fd_sc_hd__nor2_1_0/Y
+ a_24_n198# mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# VSUBS mux
Xsky130_fd_sc_hd__buf_1_0 VSS VDD buf_out OUT VSUBS VDD sky130_fd_sc_hd__buf_1_0/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__inv_1_0 li_80_172# VDD VSS VDD sky130_fd_sc_hd__inv_1_0/w_42_21#
+ a_24_n198# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1_1 a_24_n198# VDD VSS VDD sky130_fd_sc_hd__inv_1_1/w_42_21#
+ C VSUBS sky130_fd_sc_hd__inv_1#0
Xdemux_0 sky130_fd_sc_hd__nor2_1_1/B demux_0/2/VSUBS VDD VSS li_80_172# IN a_24_n198#
+ demux_0/1/w_n151_n91# sky130_fd_sc_hd__nor2_1_0/B VSUBS demux
.ends

.subckt unitcell2buf_32 IN C OUT buf_out VDD RESET VSS VSUBS
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_1_0/B sky130_fd_sc_hd__nor2_1_0/Y
+ RESET VSS VDD VSUBS VDD sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_1/B sky130_fd_sc_hd__nor2_1_1/Y
+ RESET VSS VDD VSUBS VDD sky130_fd_sc_hd__nor2_1_1/a_109_297# sky130_fd_sc_hd__nor2_1
X1 sky130_fd_sc_hd__nor2_1_0/B VDD VDD li_80_172# sky130_fd_pr__pfet_01v8_hvt_UUWA33
X2 VDD sky130_fd_sc_hd__nor2_1_1/B VDD a_24_n198# sky130_fd_pr__pfet_01v8_hvt_UUWA33
Xmux_0 mux_0/2/VSUBS VDD VSS li_80_172# OUT sky130_fd_sc_hd__nor2_1_1/Y sky130_fd_sc_hd__nor2_1_0/Y
+ a_24_n198# mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# VSUBS mux
Xsky130_fd_sc_hd__buf_1_0 VSS VDD buf_out OUT VSUBS VDD sky130_fd_sc_hd__buf_1_0/a_27_47#
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__inv_1_0 li_80_172# VDD VSS VDD sky130_fd_sc_hd__inv_1_0/w_42_21#
+ a_24_n198# VSUBS sky130_fd_sc_hd__inv_1#0
Xsky130_fd_sc_hd__inv_1_1 a_24_n198# VDD VSS VDD sky130_fd_sc_hd__inv_1_1/w_42_21#
+ C VSUBS sky130_fd_sc_hd__inv_1#0
Xdemux_0 sky130_fd_sc_hd__nor2_1_1/B demux_0/2/VSUBS VDD VSS li_80_172# IN a_24_n198#
+ demux_0/1/w_n151_n91# sky130_fd_sc_hd__nor2_1_0/B VSUBS demux
.ends

.subckt brbufhalf_32 unitcell2buf_32_9/C unitcell2buf_32_0/C unitcell2bufcut_32_0/buf_out
+ unitcell2buf_32_10/C unitcell2buf_32_2/C unitcell2buf_32_12/C unitcell2buf_32_4/C
+ unitcell2bufcut_32_1/C unitcell2buf_32_6/C unitcell2buf_32_8/C sky130_fd_sc_hd__inv_16_3/A
+ unitcell2buf_32_1/C unitcell2buf_32_11/C sky130_fd_sc_hd__inv_16_3/VGND unitcell2buf_32_3/C
+ unitcell2bufcut_32_0/C unitcell2buf_32_5/C unitcell2buf_32_11/IN unitcell2bufcut_32_0/OUT
+ unitcell2buf_32_7/C sky130_fd_sc_hd__inv_16_1/A unitcell2buf_32_9/RESET unitcell2buf_32_9/VSS
+ sky130_fd_sc_hd__inv_16_1/VGND unitcell2buf_32_9/VDD VSUBS
Xsky130_fd_sc_hd__inv_16_3 unitcell2buf_32_9/RESET sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__inv_16_3/VGND
+ unitcell2buf_32_9/VDD VSUBS unitcell2buf_32_9/VDD sky130_fd_sc_hd__inv_16
Xunitcell2bufcut_32_0 unitcell2buf_32_0/OUT unitcell2bufcut_32_0/C unitcell2buf_32_9/VDD
+ unitcell2bufcut_32_0/OUT unitcell2bufcut_32_0/buf_out unitcell2buf_32_6/RESET unitcell2buf_32_9/VSS
+ VSUBS unitcell2bufcut_32
Xunitcell2buf_32_0 unitcell2buf_32_0/IN unitcell2buf_32_0/C unitcell2buf_32_0/OUT
+ unitcell2buf_32_0/buf_out unitcell2buf_32_9/VDD unitcell2buf_32_6/RESET unitcell2buf_32_9/VSS
+ VSUBS unitcell2buf_32
Xunitcell2buf_32_1 unitcell2buf_32_1/IN unitcell2buf_32_1/C unitcell2buf_32_0/IN unitcell2buf_32_1/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_6/RESET unitcell2buf_32_9/VSS VSUBS unitcell2buf_32
Xunitcell2bufcut_32_1 unitcell2buf_32_7/OUT unitcell2bufcut_32_1/C unitcell2buf_32_9/VDD
+ unitcell2buf_32_6/IN unitcell2bufcut_32_1/buf_out unitcell2buf_32_9/RESET unitcell2buf_32_9/VSS
+ VSUBS unitcell2bufcut_32
Xunitcell2buf_32_10 unitcell2buf_32_10/IN unitcell2buf_32_10/C unitcell2buf_32_9/IN
+ unitcell2buf_32_10/buf_out unitcell2buf_32_9/VDD unitcell2buf_32_9/RESET unitcell2buf_32_9/VSS
+ VSUBS unitcell2buf_32
Xunitcell2buf_32_2 unitcell2buf_32_2/IN unitcell2buf_32_2/C unitcell2buf_32_1/IN unitcell2buf_32_2/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_6/RESET unitcell2buf_32_9/VSS VSUBS unitcell2buf_32
Xunitcell2buf_32_12 unitcell2buf_32_12/IN unitcell2buf_32_12/C unitcell2buf_32_10/IN
+ unitcell2buf_32_12/buf_out unitcell2buf_32_9/VDD unitcell2buf_32_9/RESET unitcell2buf_32_9/VSS
+ VSUBS unitcell2buf_32
Xunitcell2buf_32_11 unitcell2buf_32_11/IN unitcell2buf_32_11/C unitcell2buf_32_12/IN
+ unitcell2buf_32_11/buf_out unitcell2buf_32_9/VDD unitcell2buf_32_9/RESET unitcell2buf_32_9/VSS
+ VSUBS unitcell2buf_32
Xunitcell2buf_32_3 unitcell2buf_32_3/IN unitcell2buf_32_3/C unitcell2buf_32_2/IN unitcell2buf_32_3/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_6/RESET unitcell2buf_32_9/VSS VSUBS unitcell2buf_32
Xunitcell2buf_32_4 unitcell2buf_32_4/IN unitcell2buf_32_4/C unitcell2buf_32_3/IN unitcell2buf_32_4/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_6/RESET unitcell2buf_32_9/VSS VSUBS unitcell2buf_32
Xunitcell2buf_32_5 unitcell2buf_32_5/IN unitcell2buf_32_5/C unitcell2buf_32_4/IN unitcell2buf_32_5/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_6/RESET unitcell2buf_32_9/VSS VSUBS unitcell2buf_32
Xunitcell2buf_32_6 unitcell2buf_32_6/IN unitcell2buf_32_6/C unitcell2buf_32_5/IN unitcell2buf_32_6/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_6/RESET unitcell2buf_32_9/VSS VSUBS unitcell2buf_32
Xunitcell2buf_32_7 unitcell2buf_32_7/IN unitcell2buf_32_7/C unitcell2buf_32_7/OUT
+ unitcell2buf_32_7/buf_out unitcell2buf_32_9/VDD unitcell2buf_32_9/RESET unitcell2buf_32_9/VSS
+ VSUBS unitcell2buf_32
Xunitcell2buf_32_8 unitcell2buf_32_8/IN unitcell2buf_32_8/C unitcell2buf_32_7/IN unitcell2buf_32_8/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_9/RESET unitcell2buf_32_9/VSS VSUBS unitcell2buf_32
Xunitcell2buf_32_9 unitcell2buf_32_9/IN unitcell2buf_32_9/C unitcell2buf_32_8/IN unitcell2buf_32_9/buf_out
+ unitcell2buf_32_9/VDD unitcell2buf_32_9/RESET unitcell2buf_32_9/VSS VSUBS unitcell2buf_32
Xsky130_fd_sc_hd__inv_16_0 unitcell2buf_32_6/RESET sky130_fd_sc_hd__inv_16_1/A sky130_fd_sc_hd__inv_16_1/VGND
+ unitcell2buf_32_9/VDD VSUBS unitcell2buf_32_9/VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 unitcell2buf_32_6/RESET sky130_fd_sc_hd__inv_16_1/A sky130_fd_sc_hd__inv_16_1/VGND
+ unitcell2buf_32_9/VDD VSUBS unitcell2buf_32_9/VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 unitcell2buf_32_9/RESET sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__inv_16_3/VGND
+ unitcell2buf_32_9/VDD VSUBS unitcell2buf_32_9/VDD sky130_fd_sc_hd__inv_16
.ends

.subckt sky130_fd_sc_hd__inv_8 A Y VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_2 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt invcell sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_8_0/VGND
+ sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__inv_8_0/VPWR sky130_fd_sc_hd__inv_8_0/VPB
+ VSUBS
Xsky130_fd_sc_hd__inv_8_0 sky130_fd_sc_hd__inv_8_0/A sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_8_0/VGND
+ sky130_fd_sc_hd__inv_8_0/VPWR VSUBS sky130_fd_sc_hd__inv_8_0/VPB sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__inv_2_0 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_8_0/A sky130_fd_sc_hd__inv_8_0/VPWR
+ sky130_fd_sc_hd__inv_8_0/VGND VSUBS sky130_fd_sc_hd__inv_8_0/VPB sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__inv_8_0/Y
+ sky130_fd_sc_hd__inv_8_0/VGND sky130_fd_sc_hd__inv_8_0/VPWR VSUBS sky130_fd_sc_hd__inv_8_0/VPB
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_8_0/Y
+ sky130_fd_sc_hd__inv_8_0/VGND sky130_fd_sc_hd__inv_8_0/VPWR VSUBS sky130_fd_sc_hd__inv_8_0/VPB
+ sky130_fd_sc_hd__inv_16
.ends

.subckt BR32 C[31] C[30] C[29] C[28] C[27] C[26] C[25] C[24] C[23] C[22] C[21] C[20]
+ C[19] C[18] C[17] C[16] C[15] C[14] C[13] C[12] C[11] C[10] C[9] C[8] C[7] C[6]
+ C[5] C[4] C[3] C[2] C[1] C[0] VSS VDD RESET OUT
Xbrbufhalf_32_0 C[20] C[30] OUT C[19] C[28] C[18] C[26] C[23] C[24] C[21] invcell_0/sky130_fd_sc_hd__inv_16_1/Y
+ C[29] C[17] VSS C[27] C[31] C[25] unitcell2buf_32_1/OUT brbufhalf_32_1/unitcell2buf_32_11/IN
+ C[22] invcell_0/sky130_fd_sc_hd__inv_16_0/Y unitcell2buf_32_1/RESET VSS VSS VDD
+ VSS brbufhalf_32
Xbrbufhalf_32_1 C[3] C[13] brbufhalf_32_1/unitcell2bufcut_32_0/buf_out C[2] C[11]
+ C[1] C[9] C[6] C[7] C[4] invcell_0/sky130_fd_sc_hd__inv_16_0/Y C[12] C[0] VSS C[10]
+ C[14] C[8] brbufhalf_32_1/unitcell2buf_32_11/IN unitcell2buf_32_0/IN C[5] invcell_0/sky130_fd_sc_hd__inv_16_1/Y
+ brbufhalf_32_1/unitcell2buf_32_9/RESET VSS VSS VDD VSS brbufhalf_32
Xinvcell_0 RESET invcell_0/sky130_fd_sc_hd__inv_16_1/Y VSS invcell_0/sky130_fd_sc_hd__inv_16_0/Y
+ VDD VDD VSS invcell
Xunitcell2buf_32_0 unitcell2buf_32_0/IN C[15] unitcell2buf_32_1/IN unitcell2buf_32_0/buf_out
+ VDD unitcell2buf_32_1/RESET VSS VSS unitcell2buf_32
Xunitcell2buf_32_1 unitcell2buf_32_1/IN C[16] unitcell2buf_32_1/OUT unitcell2buf_32_1/buf_out
+ VDD unitcell2buf_32_1/RESET VSS VSS unitcell2buf_32
.ends

.subckt sky130_fd_sc_hd__o22ai_1 A2 B1 Y A1 B2 VGND VPWR VNB VPB
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A1 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_307_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 A1 B1 Y VNB VPB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt brbufhalf_128 unitcell2bufcut_1/li_n460_n386# unitcell2buf_7/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/A unitcell2buf_2/li_n460_n386# unitcell2buf_11/m2_136_462#
+ sky130_fd_sc_hd__inv_16_2/VGND unitcell2buf_10/li_n460_n386# unitcell2buf_5/li_n460_n386#
+ unitcell2buf_8/li_n460_n386# unitcell2buf_0/li_n460_n386# sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_3/VGND unitcell2buf_3/li_n460_n386# unitcell2buf_11/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16_0/VGND unitcell2buf_6/li_n460_n386#
+ unitcell2bufcut_0/li_n460_n386# unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_9/li_n460_n386#
+ unitcell2buf_1/li_n460_n386# unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_1/VGND
+ VSUBS unitcell2buf_12/li_n460_n386#
Xunitcell2buf_1 unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_1/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_1/demux_0/w_18_n122#
+ unitcell2buf_1/demux_0/1/w_n151_n91# unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_1/li_n460_n386#
+ unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_1/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_1/li_80_172# unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_1/mux_0/w_18_n122# unitcell2buf_1/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_1/a_24_n198# unitcell2buf_1/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_1/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16_3/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_2 unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_2/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_2/demux_0/w_18_n122#
+ unitcell2buf_2/demux_0/1/w_n151_n91# unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_2/li_n460_n386#
+ unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_2/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_2/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_2/li_80_172# unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_2/mux_0/w_18_n122# unitcell2buf_2/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_2/a_24_n198# unitcell2buf_2/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_2/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_3 unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_3/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_3/demux_0/w_18_n122#
+ unitcell2buf_3/demux_0/1/w_n151_n91# unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_3/li_n460_n386#
+ unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_3/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_3/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_3/li_80_172# unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_3/mux_0/w_18_n122# unitcell2buf_3/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_3/a_24_n198# unitcell2buf_3/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_3/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_4 unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_4/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_4/demux_0/w_18_n122#
+ unitcell2buf_4/demux_0/1/w_n151_n91# unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_4/li_n460_n386#
+ unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_4/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_4/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_4/li_80_172# unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_4/mux_0/w_18_n122# unitcell2buf_4/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_4/a_24_n198# unitcell2buf_4/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_4/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_5 unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_5/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_5/demux_0/w_18_n122#
+ unitcell2buf_5/demux_0/1/w_n151_n91# unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_5/li_n460_n386#
+ unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_5/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_5/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_5/li_80_172# unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_5/mux_0/w_18_n122# unitcell2buf_5/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_5/a_24_n198# unitcell2buf_5/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_5/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_6 unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_6/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_6/demux_0/w_18_n122#
+ unitcell2buf_6/demux_0/1/w_n151_n91# unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_6/li_n460_n386#
+ unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_6/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_6/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_6/li_80_172# unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/Y unitcell2bufcut_1/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_6/mux_0/w_18_n122# unitcell2buf_6/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_6/a_24_n198# unitcell2buf_6/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_6/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_7 unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_7/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_7/demux_0/w_18_n122#
+ unitcell2buf_7/demux_0/1/w_n151_n91# unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_7/li_n460_n386#
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_7/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_7/li_80_172# unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_7/mux_0/w_18_n122# unitcell2buf_7/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_7/a_24_n198# unitcell2buf_7/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_7/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_8 unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_8/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_8/demux_0/w_18_n122#
+ unitcell2buf_8/demux_0/1/w_n151_n91# unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_8/li_n460_n386#
+ unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_8/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_8/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_8/li_80_172# unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_8/mux_0/w_18_n122# unitcell2buf_8/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_8/a_24_n198# unitcell2buf_8/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_8/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_9 unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_9/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_9/demux_0/w_18_n122#
+ unitcell2buf_9/demux_0/1/w_n151_n91# unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_9/li_n460_n386#
+ unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_9/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_9/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_9/li_80_172# unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_9/mux_0/w_18_n122# unitcell2buf_9/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_3/Y unitcell2buf_9/a_24_n198# unitcell2buf_9/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_9/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xunitcell2buf_10 unitcell2buf_10/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_10/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_10/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_10/demux_0/w_18_n122#
+ unitcell2buf_10/demux_0/1/w_n151_n91# unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/X
+ unitcell2buf_10/li_n460_n386# unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_10/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_10/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_10/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_10/li_80_172# unitcell2buf_10/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_10/mux_0/w_18_n122#
+ unitcell2buf_10/sky130_fd_sc_hd__inv_1#0_0/w_42_21# sky130_fd_sc_hd__inv_16_3/Y
+ unitcell2buf_10/a_24_n198# unitcell2buf_10/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_10/sky130_fd_sc_hd__nor2_1_3/B
+ VSUBS unitcell2buf
Xunitcell2buf_11 unitcell2buf_11/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_11/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_11/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_11/demux_0/w_18_n122#
+ unitcell2buf_11/demux_0/1/w_n151_n91# unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/X
+ unitcell2buf_11/li_n460_n386# unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_11/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_11/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_11/li_80_172# unitcell2buf_11/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2buf_11/m2_136_462# sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_11/mux_0/w_18_n122#
+ unitcell2buf_11/sky130_fd_sc_hd__inv_1#0_0/w_42_21# sky130_fd_sc_hd__inv_16_3/Y
+ unitcell2buf_11/a_24_n198# unitcell2buf_11/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_11/sky130_fd_sc_hd__nor2_1_3/B
+ VSUBS unitcell2buf
Xunitcell2buf_12 unitcell2buf_12/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_12/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_12/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_12/demux_0/w_18_n122#
+ unitcell2buf_12/demux_0/1/w_n151_n91# unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/X
+ unitcell2buf_12/li_n460_n386# unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_12/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_12/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_12/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_12/li_80_172# unitcell2buf_12/sky130_fd_sc_hd__nor2_1_3/Y
+ unitcell2buf_11/sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_12/mux_0/w_18_n122#
+ unitcell2buf_12/sky130_fd_sc_hd__inv_1#0_0/w_42_21# sky130_fd_sc_hd__inv_16_3/Y
+ unitcell2buf_12/a_24_n198# unitcell2buf_12/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_12/sky130_fd_sc_hd__nor2_1_3/B
+ VSUBS unitcell2buf
Xunitcell2bufcut_0 unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2bufcut_0/sky130_fd_sc_hd__inv_1_1/w_42_21#
+ unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2bufcut_0/demux_1/1/w_n151_n91# unitcell2bufcut_0/a_24_n198# unitcell2bufcut_0/li_n460_n386#
+ unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2bufcut_0/mux_1/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2bufcut_0/li_80_172# unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/X unitcell2bufcut_0/sky130_fd_sc_hd__inv_1_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2bufcut_0/sky130_fd_sc_hd__nor2_1_3/B VSUBS
+ VSUBS unitcell2bufcut
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_0/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2bufcut_1 unitcell2bufcut_1/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2bufcut_1/sky130_fd_sc_hd__inv_1_1/w_42_21#
+ unitcell2bufcut_1/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2bufcut_1/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2bufcut_1/demux_1/1/w_n151_n91# unitcell2bufcut_1/a_24_n198# unitcell2bufcut_1/li_n460_n386#
+ unitcell2bufcut_1/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2bufcut_1/mux_1/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2bufcut_1/li_80_172# unitcell2bufcut_1/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut_1/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_7/sky130_fd_sc_hd__buf_1_1/A unitcell2bufcut_1/sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2bufcut_1/sky130_fd_sc_hd__buf_1_1/X unitcell2bufcut_1/sky130_fd_sc_hd__inv_1_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_3/Y unitcell2bufcut_1/sky130_fd_sc_hd__nor2_1_3/B VSUBS
+ VSUBS unitcell2bufcut
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_1/A
+ sky130_fd_sc_hd__inv_16_1/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
Xunitcell2buf_0 unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_0/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_0/demux_0/w_18_n122#
+ unitcell2buf_0/demux_0/1/w_n151_n91# unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/X unitcell2buf_0/li_n460_n386#
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/a_27_47# unitcell2buf_0/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91#
+ unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/B
+ unitcell2buf_0/li_80_172# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/Y unitcell2buf_1/sky130_fd_sc_hd__buf_1_1/A
+ sky130_fd_sc_hd__inv_16_3/VPB unitcell2buf_0/mux_0/w_18_n122# unitcell2buf_0/sky130_fd_sc_hd__inv_1#0_0/w_42_21#
+ sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_0/a_24_n198# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/Y
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/B VSUBS unitcell2buf
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16_2/VGND sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB
+ sky130_fd_sc_hd__inv_16
.ends

.subckt BR128half_bottom brbufhalf_128_0/unitcell2bufcut_0/li_n460_n386# brbufhalf_2/unitcell2buf_4/li_n460_n386#
+ brbufhalf_0/unitcell2bufcut_3/li_n460_n386# brbufhalf_128_0/unitcell2buf_4/li_n460_n386#
+ brbufhalf_2/unitcell2buf_26/m2_136_462# brbufhalf_0/unitcell2buf_3/li_n460_n386#
+ brbufhalf_1/unitcell2buf_9/li_n460_n386# brbufhalf_2/unitcell2buf_26/li_n460_n386#
+ brbufhalf_2/unitcell2bufcut_2/li_n460_n386# brbufhalf_1/unitcell2buf_1/li_n460_n386#
+ brbufhalf_0/unitcell2buf_24/li_n460_n386# brbufhalf_2/unitcell2buf_7/li_n460_n386#
+ brbufhalf_128_0/unitcell2buf_7/li_n460_n386# brbufhalf_128_0/unitcell2buf_11/li_n460_n386#
+ brbufhalf_0/unitcell2buf_6/li_n460_n386# brbufhalf_0/unitcell2buf_27/li_n460_n386#
+ brbufhalf_1/unitcell2buf_4/li_n460_n386# brbufhalf_1/unitcell2buf_24/li_n460_n386#
+ brbufhalf_1/unitcell2bufcut_3/li_n460_n386# sky130_fd_sc_hd__inv_16_3/A brbufhalf_2/unitcell2buf_2/li_n460_n386#
+ brbufhalf_0/unitcell2buf_9/li_n460_n386# brbufhalf_128_0/unitcell2buf_11/m2_136_462#
+ brbufhalf_128_0/unitcell2buf_2/li_n460_n386# brbufhalf_0/unitcell2buf_1/li_n460_n386#
+ brbufhalf_1/unitcell2buf_7/li_n460_n386# brbufhalf_1/unitcell2buf_27/li_n460_n386#
+ brbufhalf_128_0/unitcell2bufcut_1/li_n460_n386# brbufhalf_2/unitcell2buf_24/li_n460_n386#
+ brbufhalf_2/unitcell2buf_5/li_n460_n386# brbufhalf_128_0/unitcell2buf_5/li_n460_n386#
+ brbufhalf_0/unitcell2buf_4/li_n460_n386# brbufhalf_0/unitcell2buf_25/li_n460_n386#
+ brbufhalf_2/unitcell2buf_27/li_n460_n386# brbufhalf_1/unitcell2buf_2/li_n460_n386#
+ brbufhalf_2/unitcell2bufcut_3/li_n460_n386# brbufhalf_2/unitcell2buf_8/li_n460_n386#
+ brbufhalf_128_0/unitcell2buf_8/li_n460_n386# brbufhalf_2/unitcell2buf_0/li_n460_n386#
+ brbufhalf_128_0/unitcell2buf_12/li_n460_n386# brbufhalf_0/unitcell2buf_7/li_n460_n386#
+ brbufhalf_128_0/unitcell2buf_0/li_n460_n386# brbufhalf_1/unitcell2buf_5/li_n460_n386#
+ brbufhalf_1/unitcell2buf_25/li_n460_n386# brbufhalf_2/unitcell2buf_3/li_n460_n386#
+ brbufhalf_0/unitcell2bufcut_2/li_n460_n386# brbufhalf_128_0/unitcell2buf_3/li_n460_n386#
+ brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A brbufhalf_0/unitcell2buf_2/li_n460_n386#
+ brbufhalf_1/unitcell2buf_8/li_n460_n386# brbufhalf_2/unitcell2buf_25/li_n460_n386#
+ brbufhalf_2/unitcell2buf_6/li_n460_n386# brbufhalf_1/unitcell2buf_0/li_n460_n386#
+ brbufhalf_128_0/unitcell2buf_6/li_n460_n386# brbufhalf_128_0/unitcell2buf_10/li_n460_n386#
+ brbufhalf_0/unitcell2buf_5/li_n460_n386# brbufhalf_0/unitcell2buf_26/li_n460_n386#
+ brbufhalf_1/unitcell2buf_3/li_n460_n386# brbufhalf_2/unitcell2buf_9/li_n460_n386#
+ brbufhalf_1/unitcell2bufcut_2/li_n460_n386# brbufhalf_128_0/unitcell2buf_9/li_n460_n386#
+ brbufhalf_2/unitcell2buf_1/li_n460_n386# brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_0/unitcell2buf_8/li_n460_n386# brbufhalf_128_0/unitcell2buf_1/li_n460_n386#
+ brbufhalf_0/unitcell2buf_0/li_n460_n386# brbufhalf_1/unitcell2buf_6/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/VPB VSUBS brbufhalf_1/unitcell2buf_26/li_n460_n386#
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xbrbufhalf_0 brbufhalf_0/unitcell2buf_7/li_n460_n386# brbufhalf_0/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_1/Y brbufhalf_0/unitcell2buf_2/li_n460_n386# brbufhalf_0/unitcell2buf_24/li_n460_n386#
+ VSUBS brbufhalf_0/unitcell2buf_5/li_n460_n386# brbufhalf_0/unitcell2buf_27/li_n460_n386#
+ brbufhalf_0/unitcell2buf_8/li_n460_n386# brbufhalf_0/unitcell2buf_0/li_n460_n386#
+ brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X brbufhalf_0/unitcell2buf_3/li_n460_n386#
+ VSUBS brbufhalf_0/unitcell2buf_25/li_n460_n386# brbufhalf_0/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_0/unitcell2buf_6/li_n460_n386# VSUBS brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_0/sky130_fd_sc_hd__inv_16_7/Y brbufhalf_0/unitcell2buf_9/li_n460_n386#
+ brbufhalf_0/unitcell2buf_1/li_n460_n386# brbufhalf_0/sky130_fd_sc_hd__inv_16_5/Y
+ brbufhalf_0/unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_1/Y brbufhalf_128_0/unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS VSUBS brbufhalf_0/unitcell2buf_26/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ brbufhalf
Xbrbufhalf_1 brbufhalf_1/unitcell2buf_7/li_n460_n386# brbufhalf_1/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/Y brbufhalf_1/unitcell2buf_2/li_n460_n386# brbufhalf_1/unitcell2buf_24/li_n460_n386#
+ VSUBS brbufhalf_1/unitcell2buf_5/li_n460_n386# brbufhalf_1/unitcell2buf_27/li_n460_n386#
+ brbufhalf_1/unitcell2buf_8/li_n460_n386# brbufhalf_1/unitcell2buf_0/li_n460_n386#
+ brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X brbufhalf_1/unitcell2buf_3/li_n460_n386#
+ VSUBS brbufhalf_1/unitcell2buf_25/li_n460_n386# brbufhalf_1/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_1/unitcell2buf_6/li_n460_n386# VSUBS brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_1/sky130_fd_sc_hd__inv_16_7/Y brbufhalf_1/unitcell2buf_9/li_n460_n386#
+ brbufhalf_1/unitcell2buf_1/li_n460_n386# brbufhalf_1/sky130_fd_sc_hd__inv_16_5/Y
+ brbufhalf_1/unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_3/Y brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS VSUBS brbufhalf_1/unitcell2buf_26/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ brbufhalf
Xbrbufhalf_2 brbufhalf_2/unitcell2buf_7/li_n460_n386# brbufhalf_2/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_1/Y brbufhalf_2/unitcell2buf_2/li_n460_n386# brbufhalf_2/unitcell2buf_24/li_n460_n386#
+ VSUBS brbufhalf_2/unitcell2buf_5/li_n460_n386# brbufhalf_2/unitcell2buf_27/li_n460_n386#
+ brbufhalf_2/unitcell2buf_8/li_n460_n386# brbufhalf_2/unitcell2buf_0/li_n460_n386#
+ brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X brbufhalf_2/unitcell2buf_3/li_n460_n386#
+ VSUBS brbufhalf_2/unitcell2buf_25/li_n460_n386# brbufhalf_2/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_2/unitcell2buf_6/li_n460_n386# VSUBS brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_2/sky130_fd_sc_hd__inv_16_7/Y brbufhalf_2/unitcell2buf_9/li_n460_n386#
+ brbufhalf_2/unitcell2buf_1/li_n460_n386# brbufhalf_2/sky130_fd_sc_hd__inv_16_5/Y
+ brbufhalf_2/unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_1/Y brbufhalf_2/unitcell2buf_26/m2_136_462#
+ VSUBS VSUBS brbufhalf_2/unitcell2buf_26/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ brbufhalf
Xbrbufhalf_128_0 brbufhalf_128_0/unitcell2bufcut_1/li_n460_n386# brbufhalf_128_0/unitcell2buf_7/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/Y brbufhalf_128_0/unitcell2buf_2/li_n460_n386# brbufhalf_128_0/unitcell2buf_11/m2_136_462#
+ VSUBS brbufhalf_128_0/unitcell2buf_10/li_n460_n386# brbufhalf_128_0/unitcell2buf_5/li_n460_n386#
+ brbufhalf_128_0/unitcell2buf_8/li_n460_n386# brbufhalf_128_0/unitcell2buf_0/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/Y VSUBS brbufhalf_128_0/unitcell2buf_3/li_n460_n386# brbufhalf_128_0/unitcell2buf_11/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/VPB VSUBS brbufhalf_128_0/unitcell2buf_6/li_n460_n386#
+ brbufhalf_128_0/unitcell2bufcut_0/li_n460_n386# brbufhalf_128_0/unitcell2bufcut_0/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_128_0/unitcell2buf_9/li_n460_n386# brbufhalf_128_0/unitcell2buf_1/li_n460_n386#
+ brbufhalf_128_0/unitcell2buf_4/li_n460_n386# VSUBS VSUBS brbufhalf_128_0/unitcell2buf_12/li_n460_n386#
+ brbufhalf_128
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
.ends

.subckt BR128half brbufhalf_2/unitcell2buf_4/li_n460_n386# brbufhalf_0/unitcell2bufcut_3/li_n460_n386#
+ brbufhalf_0/unitcell2buf_3/li_n460_n386# brbufhalf_3/unitcell2buf_2/li_n460_n386#
+ brbufhalf_1/unitcell2buf_9/li_n460_n386# brbufhalf_2/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_2/unitcell2buf_26/li_n460_n386# brbufhalf_1/unitcell2buf_1/li_n460_n386#
+ brbufhalf_0/unitcell2buf_24/li_n460_n386# brbufhalf_2/unitcell2buf_7/li_n460_n386#
+ brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A brbufhalf_0/unitcell2buf_6/li_n460_n386#
+ brbufhalf_3/unitcell2buf_5/li_n460_n386# brbufhalf_1/unitcell2buf_4/li_n460_n386#
+ brbufhalf_0/unitcell2buf_27/li_n460_n386# brbufhalf_1/unitcell2buf_24/li_n460_n386#
+ brbufhalf_3/unitcell2buf_26/li_n460_n386# brbufhalf_1/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/A brbufhalf_1/unitcell2buf_26/m2_136_462# brbufhalf_2/unitcell2buf_2/li_n460_n386#
+ brbufhalf_0/unitcell2buf_9/li_n460_n386# brbufhalf_3/unitcell2buf_8/li_n460_n386#
+ brbufhalf_3/unitcell2buf_0/li_n460_n386# brbufhalf_0/unitcell2buf_1/li_n460_n386#
+ brbufhalf_3/unitcell2bufcut_2/li_n460_n386# brbufhalf_1/unitcell2buf_7/li_n460_n386#
+ brbufhalf_1/unitcell2buf_27/li_n460_n386# brbufhalf_2/unitcell2buf_24/li_n460_n386#
+ brbufhalf_2/unitcell2buf_5/li_n460_n386# brbufhalf_0/unitcell2buf_4/li_n460_n386#
+ brbufhalf_3/unitcell2buf_3/li_n460_n386# brbufhalf_2/unitcell2bufcut_3/li_n460_n386#
+ brbufhalf_2/unitcell2buf_27/li_n460_n386# brbufhalf_0/unitcell2buf_25/li_n460_n386#
+ brbufhalf_1/unitcell2buf_2/li_n460_n386# brbufhalf_2/unitcell2buf_8/li_n460_n386#
+ brbufhalf_3/unitcell2buf_24/li_n460_n386# brbufhalf_2/unitcell2buf_0/li_n460_n386#
+ brbufhalf_3/unitcell2buf_6/li_n460_n386# brbufhalf_0/unitcell2buf_7/li_n460_n386#
+ brbufhalf_1/unitcell2buf_5/li_n460_n386# brbufhalf_3/unitcell2buf_27/li_n460_n386#
+ brbufhalf_1/unitcell2buf_25/li_n460_n386# brbufhalf_3/unitcell2buf_9/li_n460_n386#
+ brbufhalf_2/unitcell2buf_3/li_n460_n386# brbufhalf_0/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A brbufhalf_0/unitcell2buf_2/li_n460_n386#
+ brbufhalf_3/unitcell2buf_1/li_n460_n386# brbufhalf_1/unitcell2buf_8/li_n460_n386#
+ brbufhalf_3/unitcell2bufcut_3/li_n460_n386# brbufhalf_2/unitcell2buf_25/li_n460_n386#
+ brbufhalf_2/unitcell2buf_6/li_n460_n386# brbufhalf_1/unitcell2buf_0/li_n460_n386#
+ brbufhalf_0/unitcell2buf_5/li_n460_n386# brbufhalf_3/unitcell2buf_4/li_n460_n386#
+ brbufhalf_2/sky130_fd_sc_hd__inv_16_5/Y brbufhalf_3/unitcell2buf_26/m2_136_462#
+ brbufhalf_0/unitcell2buf_26/li_n460_n386# brbufhalf_1/unitcell2buf_3/li_n460_n386#
+ brbufhalf_2/unitcell2buf_9/li_n460_n386# brbufhalf_3/unitcell2buf_25/li_n460_n386#
+ brbufhalf_1/unitcell2bufcut_2/li_n460_n386# brbufhalf_2/unitcell2buf_1/li_n460_n386#
+ brbufhalf_3/unitcell2buf_7/li_n460_n386# brbufhalf_0/unitcell2buf_8/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/VPB brbufhalf_0/unitcell2buf_0/li_n460_n386# brbufhalf_1/unitcell2buf_6/li_n460_n386#
+ VSUBS brbufhalf_1/unitcell2buf_26/li_n460_n386#
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xbrbufhalf_0 brbufhalf_0/unitcell2buf_7/li_n460_n386# brbufhalf_0/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_1/Y brbufhalf_0/unitcell2buf_2/li_n460_n386# brbufhalf_0/unitcell2buf_24/li_n460_n386#
+ VSUBS brbufhalf_0/unitcell2buf_5/li_n460_n386# brbufhalf_0/unitcell2buf_27/li_n460_n386#
+ brbufhalf_0/unitcell2buf_8/li_n460_n386# brbufhalf_0/unitcell2buf_0/li_n460_n386#
+ brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X brbufhalf_0/unitcell2buf_3/li_n460_n386#
+ VSUBS brbufhalf_0/unitcell2buf_25/li_n460_n386# brbufhalf_0/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_0/unitcell2buf_6/li_n460_n386# VSUBS brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_0/sky130_fd_sc_hd__inv_16_7/Y brbufhalf_0/unitcell2buf_9/li_n460_n386#
+ brbufhalf_0/unitcell2buf_1/li_n460_n386# brbufhalf_0/sky130_fd_sc_hd__inv_16_5/Y
+ brbufhalf_0/unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_1/Y brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS VSUBS brbufhalf_0/unitcell2buf_26/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ brbufhalf
Xbrbufhalf_1 brbufhalf_1/unitcell2buf_7/li_n460_n386# brbufhalf_1/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/Y brbufhalf_1/unitcell2buf_2/li_n460_n386# brbufhalf_1/unitcell2buf_24/li_n460_n386#
+ VSUBS brbufhalf_1/unitcell2buf_5/li_n460_n386# brbufhalf_1/unitcell2buf_27/li_n460_n386#
+ brbufhalf_1/unitcell2buf_8/li_n460_n386# brbufhalf_1/unitcell2buf_0/li_n460_n386#
+ brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X brbufhalf_1/unitcell2buf_3/li_n460_n386#
+ VSUBS brbufhalf_1/unitcell2buf_25/li_n460_n386# brbufhalf_1/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_1/unitcell2buf_6/li_n460_n386# VSUBS brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_1/sky130_fd_sc_hd__inv_16_7/Y brbufhalf_1/unitcell2buf_9/li_n460_n386#
+ brbufhalf_1/unitcell2buf_1/li_n460_n386# brbufhalf_1/sky130_fd_sc_hd__inv_16_5/Y
+ brbufhalf_1/unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_3/Y brbufhalf_1/unitcell2buf_26/m2_136_462#
+ VSUBS VSUBS brbufhalf_1/unitcell2buf_26/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ brbufhalf
Xbrbufhalf_2 brbufhalf_2/unitcell2buf_7/li_n460_n386# brbufhalf_2/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_3/Y brbufhalf_2/unitcell2buf_2/li_n460_n386# brbufhalf_2/unitcell2buf_24/li_n460_n386#
+ VSUBS brbufhalf_2/unitcell2buf_5/li_n460_n386# brbufhalf_2/unitcell2buf_27/li_n460_n386#
+ brbufhalf_2/unitcell2buf_8/li_n460_n386# brbufhalf_2/unitcell2buf_0/li_n460_n386#
+ brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X brbufhalf_2/unitcell2buf_3/li_n460_n386#
+ VSUBS brbufhalf_2/unitcell2buf_25/li_n460_n386# brbufhalf_2/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_2/unitcell2buf_6/li_n460_n386# VSUBS brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_2/sky130_fd_sc_hd__inv_16_7/Y brbufhalf_2/unitcell2buf_9/li_n460_n386#
+ brbufhalf_2/unitcell2buf_1/li_n460_n386# brbufhalf_2/sky130_fd_sc_hd__inv_16_5/Y
+ brbufhalf_2/unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_3/Y brbufhalf_3/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ VSUBS VSUBS brbufhalf_2/unitcell2buf_26/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ brbufhalf
Xbrbufhalf_3 brbufhalf_3/unitcell2buf_7/li_n460_n386# brbufhalf_3/unitcell2bufcut_3/li_n460_n386#
+ sky130_fd_sc_hd__inv_16_1/Y brbufhalf_3/unitcell2buf_2/li_n460_n386# brbufhalf_3/unitcell2buf_24/li_n460_n386#
+ VSUBS brbufhalf_3/unitcell2buf_5/li_n460_n386# brbufhalf_3/unitcell2buf_27/li_n460_n386#
+ brbufhalf_3/unitcell2buf_8/li_n460_n386# brbufhalf_3/unitcell2buf_0/li_n460_n386#
+ brbufhalf_3/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/X brbufhalf_3/unitcell2buf_3/li_n460_n386#
+ VSUBS brbufhalf_3/unitcell2buf_25/li_n460_n386# brbufhalf_3/unitcell2bufcut_2/li_n460_n386#
+ brbufhalf_3/unitcell2buf_6/li_n460_n386# VSUBS brbufhalf_3/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ brbufhalf_3/sky130_fd_sc_hd__inv_16_7/Y brbufhalf_3/unitcell2buf_9/li_n460_n386#
+ brbufhalf_3/unitcell2buf_1/li_n460_n386# brbufhalf_3/sky130_fd_sc_hd__inv_16_5/Y
+ brbufhalf_3/unitcell2buf_4/li_n460_n386# sky130_fd_sc_hd__inv_16_1/Y brbufhalf_3/unitcell2buf_26/m2_136_462#
+ VSUBS VSUBS brbufhalf_3/unitcell2buf_26/li_n460_n386# sky130_fd_sc_hd__inv_16_3/VPB
+ brbufhalf
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_16_3/Y sky130_fd_sc_hd__inv_16_3/A
+ VSUBS sky130_fd_sc_hd__inv_16_3/VPB VSUBS sky130_fd_sc_hd__inv_16_3/VPB sky130_fd_sc_hd__inv_16
.ends

.subckt BR128 RESET VDD C[0] C[1] C[2] C[3] C[4] C[5] C[7] C[8] C[9] C[10] C[11] C[12]
+ C[13] C[14] C[15] C[16] C[17] C[18] C[19] C[20] C[21] C[22] C[23] C[24] C[25] C[26]
+ C[27] C[28] C[29] C[30] C[6] C[31] C[32] C[33] C[34] C[35] C[36] C[37] C[38] C[39]
+ C[40] C[41] C[42] C[43] C[44] C[45] C[46] C[47] C[48] C[49] C[50] C[51] C[52] C[53]
+ C[54] C[55] C[56] C[57] C[58] C[59] C[60] C[61] C[62] C[95] C[96] C[97] C[98] C[99]
+ C[100] C[101] C[102] C[103] C[104] C[105] C[106] C[107] C[108] C[109] C[110] C[111]
+ C[112] C[113] C[114] C[115] C[116] C[117] C[118] C[119] C[120] C[121] C[122] C[123]
+ C[124] C[125] C[126] C[127] C[63] C[64] C[65] C[66] C[67] C[68] C[69] C[70] C[71]
+ C[72] C[73] C[74] C[75] C[76] C[77] C[78] C[79] C[80] C[81] C[82] C[83] C[84] C[85]
+ C[86] C[87] C[88] C[89] C[90] C[91] C[92] C[93] C[94] OUT VSS
XBR128half_bottom_0 C[46] C[73] C[54] C[41] BR128half_bottom_0/brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ C[58] C[83] C[63] C[78] C[92] C[50] C[69] C[37] C[32] C[55] C[48] C[89] C[82] C[86]
+ sky130_fd_sc_hd__inv_16_1/Y C[75] C[51] BR128half_0/brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ C[43] C[60] C[85] C[80] C[38] C[66] C[72] C[40] C[57] C[49] C[64] C[91] C[70] C[68]
+ C[36] C[77] C[33] C[53] C[45] C[88] C[81] C[74] C[62] C[42] BR128half_bottom_0/brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ C[59] C[84] C[65] C[71] C[93] C[39] C[34] C[56] C[47] C[90] C[67] C[94] C[35] C[76]
+ BR128half_bottom_0/brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A C[52]
+ C[44] C[61] C[87] VDD VSS C[79] BR128half_bottom
Xsky130_fd_sc_hd__inv_8_0 sky130_fd_sc_hd__inv_8_0/A sky130_fd_sc_hd__inv_8_0/Y VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__buf_2_0 VDD VSS sky130_fd_sc_hd__inv_8_0/A RESET VSS VDD sky130_fd_sc_hd__buf_2
XBR128half_0 C[121] C[23] C[27] C[107] C[4] C[126] C[111] C[13] C[19] C[117] BR128half_0/brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A
+ C[24] C[104] C[10] C[17] C[3] C[95] C[7] sky130_fd_sc_hd__inv_16_1/Y unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ C[123] C[20] C[100] C[109] C[29] C[110] C[6] C[1] C[114] C[120] C[26] C[106] C[118]
+ C[112] C[18] C[12] C[116] C[98] C[125] C[103] C[22] C[9] C[96] C[2] C[99] C[122]
+ C[31] BR128half_0/brbufhalf_0/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A C[28]
+ C[108] C[5] C[102] C[113] C[119] C[14] C[25] C[105] unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/A
+ BR128half_bottom_0/brbufhalf_1/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A C[16]
+ C[11] C[115] C[97] C[15] C[124] C[101] C[21] VDD C[30] C[8] VSS C[0] BR128half
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_8_0/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_8_0/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_16
Xunitcell2buf_0 unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/a_109_297# unitcell2buf_0/sky130_fd_sc_hd__inv_1#0_1/w_42_21#
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/a_109_297# unitcell2buf_0/demux_0/w_18_n122#
+ unitcell2buf_0/demux_0/1/w_n151_n91# OUT C[127] unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/a_27_47#
+ unitcell2buf_0/mux_0/sky130_fd_pr__nfet_01v8_PX9ZJG_1/w_n151_n91# unitcell2buf_0/sky130_fd_sc_hd__buf_1_1/A
+ unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/B unitcell2buf_0/li_80_172# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/Y
+ BR128half_0/brbufhalf_2/unitcell2bufcut_2/sky130_fd_sc_hd__buf_1_1/A VDD unitcell2buf_0/mux_0/w_18_n122#
+ unitcell2buf_0/sky130_fd_sc_hd__inv_1#0_0/w_42_21# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/A
+ unitcell2buf_0/a_24_n198# unitcell2buf_0/sky130_fd_sc_hd__nor2_1_2/Y unitcell2buf_0/sky130_fd_sc_hd__nor2_1_3/B
+ VSS unitcell2buf
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=5.36e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__buf_12 A X VGND VPWR VNB VPB
X0 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__nand2b_1 Y A_N B VGND VPWR VNB VPB
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_2 B1 Y A2 A1 VGND VPWR VNB VPB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_0 VGND VPWR Y B1 A2 A1 VNB VPB
X0 a_120_369# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 Y A2 a_120_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt puf_super reset clk si puf_sel1 puf_sel0 length1 length0 out so vccd1 rstn
+ vssd1
Xsky130_fd_sc_hd__decap_12_1780 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1791 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_7 vssd1 vccd1 BR128_3/C[126] BR128_2/C[126] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_7 sky130_fd_sc_hd__inv_6_0/A BR32_1/C[1] vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1010 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1021 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1032 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1043 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1054 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1065 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1076 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1087 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1098 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1609 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_9 sky130_fd_sc_hd__nand2_1_9/Y BR128_2/OUT sky130_fd_sc_hd__nor2_1_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_10 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_21 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_32 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_43 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_54 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_65 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_76 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_87 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_98 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_407 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_418 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_429 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1406 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1417 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1428 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1439 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_930 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_941 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_952 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_963 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_974 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_985 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_996 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_8_1 BR64_3/C[8] sky130_fd_sc_hd__clkbuf_8_1/A vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__decap_12_204 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_215 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_226 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_237 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_248 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_259 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1203 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1214 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1225 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1236 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1247 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1258 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1269 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_1 sky130_fd_sc_hd__clkinv_8_4/A sky130_fd_sc_hd__clkinv_8_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_760 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_771 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_782 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_793 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1770 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1781 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1792 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_8 vssd1 vccd1 BR128_3/C[117] BR128_2/C[117] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_8 sky130_fd_sc_hd__inv_6_1/A BR32_1/C[9] vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1000 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1011 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1022 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1033 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1044 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1055 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1066 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1077 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1088 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1099 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_590 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_11 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_22 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_33 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_44 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_55 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_66 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_77 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_88 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_99 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_408 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_419 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1407 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1418 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1429 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_920 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_931 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_942 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_953 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_964 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_975 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_986 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_997 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_8_2 BR64_3/C[6] sky130_fd_sc_hd__clkbuf_8_2/A vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__decap_12_205 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_216 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_227 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_238 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_249 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1204 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1215 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1226 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1237 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1248 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1259 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_2 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__clkinv_8_4/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_750 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_761 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_772 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_783 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_794 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1760 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1771 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1782 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1793 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_9 vssd1 vccd1 BR128_3/C[121] BR128_2/C[121] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_9 sky130_fd_sc_hd__clkinv_4_2/A BR32_2/C[5] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1001 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1012 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1023 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1034 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1045 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1056 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1067 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1078 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1089 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_580 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_591 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1590 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_10 sky130_fd_sc_hd__clkinv_4_3/A BR32_2/C[4] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_12 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_23 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_34 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_45 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_56 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_67 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_78 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_89 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_409 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1408 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1419 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_910 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_921 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_932 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_943 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_954 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_965 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_976 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_987 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_998 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_206 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_217 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_228 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_239 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_90 BR64_1/C[37] sky130_fd_sc_hd__clkbuf_4_1/A BR64_3/C[36]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1205 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1216 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1227 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1238 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1249 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_3 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__clkinv_8_4/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_740 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_751 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_762 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_773 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_784 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_795 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1750 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1761 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1772 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1783 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1794 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1002 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1013 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1024 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1035 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1046 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1057 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1068 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1079 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_570 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_581 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_592 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1580 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1591 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_1_11 sky130_fd_sc_hd__clkinv_4_4/A BR32_2/C[3] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__buf_8_0 BR32_2/C[13] BR64_3/C[13] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__decap_12_13 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_24 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_35 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_46 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_57 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_68 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_79 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1409 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_900 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_911 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_922 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_933 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_944 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_955 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_966 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_977 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_988 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_999 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_207 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_218 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_229 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_80 BR64_1/C[47] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[46]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_91 BR64_1/C[36] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[35]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1206 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1217 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1228 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1239 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_4 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__clkinv_8_4/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_730 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_741 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_752 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_763 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_774 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_785 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_796 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1740 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1751 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1762 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1773 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1784 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1795 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1003 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1014 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1025 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1036 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1047 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1058 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1069 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_560 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_571 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_582 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_593 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1570 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1581 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1592 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_390 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_14 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_25 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_36 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_47 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_58 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_69 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_901 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_912 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_923 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_934 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_945 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_956 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_967 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_978 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_989 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_208 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_219 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_70 BR64_1/C[57] sky130_fd_sc_hd__clkbuf_4_1/X BR64_3/C[56]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_81 BR64_1/C[46] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[45]
+ sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_92 BR64_1/C[35] sky130_fd_sc_hd__clkbuf_4_1/A BR64_3/C[34]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1207 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1218 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1229 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_5 sky130_fd_sc_hd__clkinv_8_8/A sky130_fd_sc_hd__clkinv_8_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_720 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_731 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_742 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_753 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_764 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_775 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_786 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_797 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1730 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1741 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1752 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1763 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1774 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1785 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1796 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1004 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1015 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1026 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1037 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1048 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1059 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_550 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_561 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_572 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_583 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_594 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1560 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1571 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1582 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1593 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_380 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_391 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1390 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_15 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_26 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_37 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_48 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_59 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nor2_1_0 reset sky130_fd_sc_hd__nor2_1_0/Y puf_sel1 vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_902 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_913 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_924 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_935 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_946 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_957 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_968 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_979 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_60 BR128_2/C[67] sky130_fd_sc_hd__clkbuf_4_1/X BR128_2/C[66]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_71 BR64_1/C[56] sky130_fd_sc_hd__clkbuf_4_1/X BR64_3/C[55]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_82 BR64_1/C[45] sky130_fd_sc_hd__clkbuf_4_1/A BR64_3/C[44]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_93 BR64_1/C[34] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[33]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1208 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1219 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_6 sky130_fd_sc_hd__clkinv_8_6/Y sky130_fd_sc_hd__clkinv_8_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_710 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_721 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_732 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_743 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_754 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_765 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_776 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_787 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_798 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1720 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1731 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1742 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1753 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1764 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1775 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1786 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1797 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1005 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1016 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1027 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1038 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1049 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_540 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_551 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_562 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_573 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_584 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_595 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1550 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1561 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1572 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1583 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1594 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_0 sky130_fd_sc_hd__clkbuf_4_1/A rstn vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_4_0 sky130_fd_sc_hd__clkinv_4_0/A BR64_3/C[31] vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_370 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_381 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_392 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1380 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1391 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_16 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_27 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_38 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_49 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_0 vccd1 vssd1 BR64_3/C[47] BR64_1/C[47] vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__inv_6_0 BR64_3/C[1] sky130_fd_sc_hd__inv_6_0/A vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__inv_6
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_1/B sky130_fd_sc_hd__nor2_1_1/Y
+ reset vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_1/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_903 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_914 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_925 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_936 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_947 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_958 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_969 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_50 sky130_fd_sc_hd__buf_6_9/A sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_0/C[76] sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_61 BR128_2/C[66] sky130_fd_sc_hd__clkbuf_4_1/X BR128_1/C[65]
+ sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_72 BR64_1/C[55] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[54]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_83 sky130_fd_sc_hd__buf_6_1/A sky130_fd_sc_hd__clkbuf_4_1/A
+ BR64_1/C[43] sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_94 BR64_1/C[33] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[32]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_7 sky130_fd_sc_hd__clkinv_8_7/Y sky130_fd_sc_hd__clkinv_8_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_700 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_711 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_722 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_733 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_744 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_755 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_766 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_777 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_788 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_799 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1710 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1721 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1732 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1743 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1754 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1765 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1776 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1787 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1798 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1006 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1017 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1028 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1039 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_530 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_541 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_552 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_563 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_574 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_585 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_596 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1540 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1551 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1562 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1573 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1584 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1595 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_1 sky130_fd_sc_hd__clkbuf_4_1/X sky130_fd_sc_hd__clkbuf_4_1/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_4_1 clk sky130_fd_sc_hd__clkinv_8_0/A vccd1 vssd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_360 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_371 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_382 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_393 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1370 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1381 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1392 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_190 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR64_0 BR64_0/OUT vccd1 BR64_0/RESET BR64_3/C[0] BR64_3/C[1] BR64_3/C[2] BR64_3/C[3]
+ BR64_3/C[4] BR64_3/C[5] BR64_3/C[6] BR64_3/C[7] BR64_3/C[8] BR64_3/C[9] BR64_3/C[10]
+ BR64_3/C[11] BR64_3/C[12] BR64_3/C[13] BR64_1/C[14] BR64_1/C[15] BR64_1/C[16] BR64_1/C[17]
+ BR64_1/C[18] BR64_1/C[19] BR64_1/C[20] BR64_1/C[21] BR64_1/C[22] BR64_3/C[23] BR64_1/C[24]
+ BR64_1/C[25] BR64_3/C[26] BR64_1/C[27] BR64_1/C[28] BR64_1/C[29] BR64_1/C[30] BR64_3/C[31]
+ BR64_1/C[32] BR64_1/C[33] BR64_1/C[34] BR64_1/C[35] BR64_1/C[36] BR64_1/C[37] BR64_1/C[38]
+ BR64_1/C[39] BR64_1/C[40] BR64_1/C[41] BR64_1/C[42] BR64_1/C[43] BR64_3/C[44] BR64_1/C[45]
+ BR64_1/C[46] BR64_1/C[47] BR64_1/C[48] BR64_1/C[49] BR64_1/C[50] BR64_1/C[51] BR64_1/C[52]
+ BR64_1/C[53] BR64_1/C[54] BR64_1/C[55] BR64_1/C[56] BR64_1/C[57] BR64_1/C[58] BR64_1/C[59]
+ BR64_1/C[60] BR64_1/C[61] BR64_1/C[62] BR64_1/C[63] vssd1 BR64
Xsky130_fd_sc_hd__decap_12_17 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_28 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_39 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_1 vccd1 vssd1 BR64_3/C[44] sky130_fd_sc_hd__buf_6_1/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__inv_6_1 BR64_3/C[9] sky130_fd_sc_hd__inv_6_1/A vccd1 vssd1 vssd1
+ vccd1 sky130_fd_sc_hd__inv_6
Xsky130_fd_sc_hd__nor2_1_2 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__nor2_1_2/Y
+ length1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_2/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_12_904 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_915 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_926 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_937 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_948 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_959 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_40 BR128_0/C[87] sky130_fd_sc_hd__clkbuf_4_1/A BR128_0/C[86]
+ sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_51 BR128_0/C[76] sky130_fd_sc_hd__clkbuf_4_1/X BR128_3/C[75]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_62 BR128_1/C[65] sky130_fd_sc_hd__clkbuf_4_1/X BR128_1/C[64]
+ sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_73 BR64_1/C[54] sky130_fd_sc_hd__clkbuf_4_1/X BR64_3/C[53]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_84 BR64_1/C[43] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[42]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_95 BR64_1/C[32] sky130_fd_sc_hd__clkbuf_4_1/A BR64_3/C[31]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkinv_8_8 sky130_fd_sc_hd__clkinv_8_8/Y sky130_fd_sc_hd__clkinv_8_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_701 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_712 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_723 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_734 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_745 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_756 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_767 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_778 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_789 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1700 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1711 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1722 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1733 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1744 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1755 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1766 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1777 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1788 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_2_0 sky130_fd_sc_hd__nor2_1_2/B puf_sel0 sky130_fd_sc_hd__nor2_1_1/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__decap_12_1799 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1007 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1018 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1029 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_520 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_531 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_542 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_553 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_564 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_575 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_586 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_597 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1530 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1541 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1552 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1563 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1574 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1585 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1596 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_2 BR64_3/C[60] BR64_1/C[60] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_4_2 sky130_fd_sc_hd__clkinv_4_2/A BR64_3/C[5] vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_350 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_361 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_372 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_383 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_394 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1360 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1371 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1382 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1393 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_180 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_10 BR32_2/RESET sky130_fd_sc_hd__o22ai_1_5/B1 sky130_fd_sc_hd__nor2_1_4/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_191 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1190 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR64_1 BR64_1/OUT vccd1 BR64_1/RESET BR64_3/C[0] BR64_3/C[1] BR64_3/C[2] BR64_3/C[3]
+ BR64_3/C[4] BR64_3/C[5] BR64_3/C[6] BR64_3/C[7] BR64_3/C[8] BR64_3/C[9] BR64_3/C[10]
+ BR64_3/C[11] BR64_3/C[12] BR64_3/C[13] BR64_1/C[14] BR64_1/C[15] BR64_1/C[16] BR64_1/C[17]
+ BR64_1/C[18] BR64_1/C[19] BR64_1/C[20] BR64_1/C[21] BR64_1/C[22] BR64_3/C[23] BR64_1/C[24]
+ BR64_1/C[25] BR64_3/C[26] BR64_1/C[27] BR64_1/C[28] BR64_1/C[29] BR64_1/C[30] BR64_3/C[31]
+ BR64_1/C[32] BR64_1/C[33] BR64_1/C[34] BR64_1/C[35] BR64_1/C[36] BR64_1/C[37] BR64_1/C[38]
+ BR64_1/C[39] BR64_1/C[40] BR64_1/C[41] BR64_1/C[42] BR64_1/C[43] BR64_3/C[44] BR64_1/C[45]
+ BR64_1/C[46] BR64_1/C[47] BR64_1/C[48] BR64_1/C[49] BR64_1/C[50] BR64_1/C[51] BR64_1/C[52]
+ BR64_1/C[53] BR64_1/C[54] BR64_1/C[55] BR64_1/C[56] BR64_1/C[57] BR64_1/C[58] BR64_1/C[59]
+ BR64_1/C[60] BR64_1/C[61] BR64_1/C[62] BR64_1/C[63] vssd1 BR64
Xsky130_fd_sc_hd__decap_12_18 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_29 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_2 vccd1 vssd1 BR64_3/C[26] sky130_fd_sc_hd__buf_6_2/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__nor2_1_3 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__nor2_1_5/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_3/a_109_297#
+ sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_3_0 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_12_905 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_916 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_927 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_938 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_949 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_30 BR128_1/C[97] rstn BR128_1/C[96] sky130_fd_sc_hd__clkinv_8_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_41 BR128_0/C[86] sky130_fd_sc_hd__clkbuf_4_1/A BR128_3/C[85]
+ sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_52 sky130_fd_sc_hd__buf_6_5/A sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_3/C[74] sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_63 BR128_1/C[64] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[63]
+ sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_74 BR64_1/C[53] sky130_fd_sc_hd__clkbuf_4_1/X BR64_3/C[52]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_85 BR64_1/C[42] sky130_fd_sc_hd__clkbuf_4_1/A BR64_3/C[41]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_96 BR32_2/C[31] sky130_fd_sc_hd__clkbuf_4_1/A BR64_3/C[30]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_702 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_713 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_724 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_735 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_746 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_757 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_120 sky130_fd_sc_hd__buf_12_1/A sky130_fd_sc_hd__clkbuf_4_1/A
+ BR64_3/C[6] sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_768 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_779 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1701 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1712 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1723 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1734 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1745 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1756 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1767 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1778 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1789 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1008 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1019 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_510 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_521 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_532 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_543 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_554 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_565 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_576 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_587 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_598 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1520 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1531 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1542 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1553 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1564 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1575 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1586 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1597 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_3 BR64_3/C[56] BR64_1/C[56] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_4_3 sky130_fd_sc_hd__clkinv_4_3/A BR64_3/C[4] vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_340 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_351 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_362 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_373 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_384 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_395 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1350 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1361 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1372 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1383 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1394 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_170 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_181 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_11 BR64_2/RESET sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__nand2_1_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_192 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1180 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1191 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR64_2 BR64_2/OUT vccd1 BR64_2/RESET BR64_3/C[0] BR64_3/C[1] BR64_3/C[2] BR64_3/C[3]
+ BR64_3/C[4] BR64_3/C[5] BR64_3/C[6] BR64_3/C[7] BR64_3/C[8] BR64_3/C[9] BR64_3/C[10]
+ BR64_3/C[11] BR64_3/C[12] BR64_3/C[13] BR64_3/C[14] BR64_3/C[15] BR64_3/C[16] BR64_3/C[17]
+ BR64_3/C[18] BR64_3/C[19] BR64_3/C[20] BR64_3/C[21] BR64_3/C[22] BR64_3/C[23] BR64_3/C[24]
+ BR64_3/C[25] BR64_3/C[26] BR64_3/C[27] BR64_3/C[28] BR64_3/C[29] BR64_3/C[30] BR64_3/C[31]
+ BR64_3/C[32] BR64_3/C[33] BR64_3/C[34] BR64_3/C[35] BR64_3/C[36] BR64_3/C[37] BR64_3/C[38]
+ BR64_3/C[39] BR64_3/C[40] BR64_3/C[41] BR64_3/C[42] BR64_3/C[43] BR64_3/C[44] BR64_3/C[45]
+ BR64_3/C[46] BR64_3/C[47] BR64_3/C[48] BR64_3/C[49] BR64_3/C[50] BR64_3/C[51] BR64_3/C[52]
+ BR64_3/C[53] BR64_3/C[54] BR64_3/C[55] BR64_3/C[56] BR64_3/C[57] BR64_3/C[58] BR64_3/C[59]
+ BR64_3/C[60] BR64_3/C[61] BR64_3/C[62] BR64_3/C[63] vssd1 BR64
Xsky130_fd_sc_hd__decap_12_19 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_3 vccd1 vssd1 BR64_3/C[23] sky130_fd_sc_hd__buf_6_3/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__nor2_1_4 sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__nor2_1_4/Y
+ sky130_fd_sc_hd__nor2_1_5/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_4/a_109_297#
+ sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_3_1 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_12_906 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_917 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_928 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_939 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_20 BR128_1/C[107] rstn BR128_1/C[106] sky130_fd_sc_hd__clkinv_8_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_31 BR128_1/C[96] sky130_fd_sc_hd__clkbuf_4_1/A BR128_1/C[95]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_42 BR128_0/C[85] sky130_fd_sc_hd__clkbuf_4_1/A BR128_0/C[84]
+ sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_53 sky130_fd_sc_hd__buf_6_6/A sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_3/C[73] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_64 BR64_1/C[63] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[62]
+ sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_75 BR64_1/C[52] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[51]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_86 BR64_1/C[41] sky130_fd_sc_hd__clkbuf_4_1/A BR64_3/C[40]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_97 BR64_1/C[30] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[29]
+ sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_703 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_714 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_725 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_736 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_747 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_110 sky130_fd_sc_hd__dfrtp_2_110/Q sky130_fd_sc_hd__clkbuf_4_1/A
+ BR32_2/C[16] sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_758 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_121 sky130_fd_sc_hd__clkbuf_8_2/A sky130_fd_sc_hd__clkbuf_4_1/X
+ BR32_2/C[5] sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_769 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1702 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1713 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1724 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1735 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1746 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1757 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1768 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1779 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1009 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR32_0 BR64_3/C[31] BR64_1/C[30] BR64_1/C[29] BR64_1/C[28] BR64_1/C[27] BR64_3/C[26]
+ BR64_1/C[25] BR64_1/C[24] BR64_3/C[23] BR64_1/C[22] BR64_1/C[21] BR64_1/C[20] BR64_1/C[19]
+ BR64_1/C[18] BR64_1/C[17] BR64_1/C[16] BR64_1/C[15] BR64_1/C[14] BR64_3/C[13] BR64_3/C[12]
+ BR64_3/C[11] BR64_3/C[10] BR32_1/C[9] BR64_3/C[8] BR64_3/C[7] BR64_3/C[6] BR64_3/C[5]
+ BR64_3/C[4] BR64_3/C[3] BR64_3/C[2] BR64_3/C[1] BR32_1/C[0] vssd1 vccd1 BR32_0/RESET
+ BR32_0/OUT BR32
Xsky130_fd_sc_hd__decap_12_500 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_511 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_522 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_533 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_544 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_555 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_566 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_577 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_588 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_599 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1510 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1521 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1532 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1543 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1554 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1565 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1576 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1587 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1598 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_4 BR64_3/C[55] BR64_1/C[55] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkinv_4_4 sky130_fd_sc_hd__clkinv_4_4/A BR64_3/C[3] vccd1 vssd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_12_330 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_341 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_352 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_363 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_374 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_385 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_396 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1340 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1351 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1362 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1373 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1384 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1395 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_160 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_171 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_182 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_12 sky130_fd_sc_hd__o21ai_1_1/B1 BR128_3/OUT sky130_fd_sc_hd__nor2_1_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_193 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1170 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1181 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1192 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR64_3 BR64_3/OUT vccd1 BR64_3/RESET BR64_3/C[0] BR64_3/C[1] BR64_3/C[2] BR64_3/C[3]
+ BR64_3/C[4] BR64_3/C[5] BR64_3/C[6] BR64_3/C[7] BR64_3/C[8] BR64_3/C[9] BR64_3/C[10]
+ BR64_3/C[11] BR64_3/C[12] BR64_3/C[13] BR64_3/C[14] BR64_3/C[15] BR64_3/C[16] BR64_3/C[17]
+ BR64_3/C[18] BR64_3/C[19] BR64_3/C[20] BR64_3/C[21] BR64_3/C[22] BR64_3/C[23] BR64_3/C[24]
+ BR64_3/C[25] BR64_3/C[26] BR64_3/C[27] BR64_3/C[28] BR64_3/C[29] BR64_3/C[30] BR64_3/C[31]
+ BR64_3/C[32] BR64_3/C[33] BR64_3/C[34] BR64_3/C[35] BR64_3/C[36] BR64_3/C[37] BR64_3/C[38]
+ BR64_3/C[39] BR64_3/C[40] BR64_3/C[41] BR64_3/C[42] BR64_3/C[43] BR64_3/C[44] BR64_3/C[45]
+ BR64_3/C[46] BR64_3/C[47] BR64_3/C[48] BR64_3/C[49] BR64_3/C[50] BR64_3/C[51] BR64_3/C[52]
+ BR64_3/C[53] BR64_3/C[54] BR64_3/C[55] BR64_3/C[56] BR64_3/C[57] BR64_3/C[58] BR64_3/C[59]
+ BR64_3/C[60] BR64_3/C[61] BR64_3/C[62] BR64_3/C[63] vssd1 BR64
Xsky130_fd_sc_hd__buf_6_4 vccd1 vssd1 BR64_3/C[0] BR32_1/C[0] vssd1 vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__nor2_1_5 sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__nor2_1_5/Y
+ sky130_fd_sc_hd__nor2_1_5/A vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_5/a_109_297#
+ sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_3_2 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_12_907 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_918 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_929 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_10 BR128_2/C[117] sky130_fd_sc_hd__clkbuf_4_1/X BR128_2/C[116]
+ sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_21 BR128_1/C[106] rstn BR128_1/C[105] sky130_fd_sc_hd__clkinv_8_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_32 BR128_1/C[95] sky130_fd_sc_hd__clkbuf_4_1/A BR128_1/C[94]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_43 BR128_0/C[84] sky130_fd_sc_hd__clkbuf_4_1/A BR128_3/C[83]
+ sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_54 sky130_fd_sc_hd__dfrtp_2_54/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_3/C[72] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_65 BR64_1/C[62] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[61]
+ sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_76 BR64_1/C[51] sky130_fd_sc_hd__clkbuf_4_1/X BR64_3/C[50]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_87 BR64_1/C[40] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[39]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_98 BR64_1/C[29] sky130_fd_sc_hd__clkbuf_4_1/A BR64_3/C[28]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_704 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_715 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_726 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_737 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_100 BR64_1/C[27] sky130_fd_sc_hd__clkbuf_4_1/A BR64_3/C[26]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_748 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_111 BR32_2/C[16] sky130_fd_sc_hd__clkbuf_4_1/A BR32_2/C[15]
+ sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_759 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_122 BR32_2/C[5] sky130_fd_sc_hd__clkbuf_4_1/X BR32_2/C[4]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1703 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1714 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1725 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1736 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1747 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1758 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1769 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR32_1 BR32_2/C[31] BR64_1/C[30] BR64_1/C[29] BR64_1/C[28] BR64_1/C[27] BR64_3/C[26]
+ BR64_1/C[25] BR64_1/C[24] BR64_3/C[23] BR64_1/C[22] BR64_1/C[21] BR64_1/C[20] BR64_1/C[19]
+ BR64_1/C[18] BR64_1/C[17] BR64_1/C[16] BR64_1/C[15] BR32_2/C[14] BR32_2/C[13] BR32_1/C[12]
+ BR64_3/C[11] BR64_3/C[10] BR32_1/C[9] BR64_3/C[8] BR64_3/C[7] BR64_3/C[6] BR32_2/C[5]
+ BR32_2/C[4] BR32_2/C[3] BR64_3/C[2] BR32_1/C[1] BR32_1/C[0] vssd1 vccd1 BR32_1/RESET
+ BR32_1/OUT BR32
Xsky130_fd_sc_hd__decap_12_501 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_512 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_523 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_534 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_545 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_556 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_567 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_578 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_589 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1500 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1511 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1522 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1533 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1544 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1555 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1566 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1577 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1588 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1599 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o22ai_1_0 sky130_fd_sc_hd__o22ai_1_2/Y sky130_fd_sc_hd__nor2_1_1/B
+ sky130_fd_sc_hd__o22ai_1_0/Y puf_sel1 sky130_fd_sc_hd__o22ai_1_1/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkbuf_4_5 BR64_3/C[53] BR64_1/C[53] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_320 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_331 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_342 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_353 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_364 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_375 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_386 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_397 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1330 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1341 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1352 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1363 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1374 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1385 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1396 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_150 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_161 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_172 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_183 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_13 BR32_3/RESET sky130_fd_sc_hd__o22ai_1_6/B1 sky130_fd_sc_hd__nor2_1_5/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_194 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1160 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1171 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1182 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1193 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_5 vccd1 vssd1 BR128_3/C[75] sky130_fd_sc_hd__buf_6_5/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__decap_3_3 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_12_908 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_919 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_11 BR128_2/C[116] sky130_fd_sc_hd__clkbuf_4_1/X BR128_2/C[115]
+ sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_22 BR128_1/C[105] sky130_fd_sc_hd__clkbuf_4_1/A BR128_1/C[104]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_33 BR128_1/C[94] sky130_fd_sc_hd__clkbuf_4_1/A BR128_1/C[93]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_44 BR128_0/C[83] sky130_fd_sc_hd__clkbuf_4_1/X BR128_3/C[82]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_55 sky130_fd_sc_hd__dfrtp_2_55/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_3/C[71] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_66 BR64_1/C[61] sky130_fd_sc_hd__clkbuf_4_1/X BR64_3/C[60]
+ sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_77 BR64_1/C[50] sky130_fd_sc_hd__clkbuf_4_1/X BR64_3/C[49]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_88 BR64_1/C[39] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[38]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_99 BR64_1/C[28] sky130_fd_sc_hd__clkbuf_4_1/A BR64_3/C[27]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_705 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_716 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_727 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_738 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_101 sky130_fd_sc_hd__buf_6_2/A sky130_fd_sc_hd__clkbuf_4_1/A
+ BR64_3/C[25] sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_749 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_112 BR32_2/C[15] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[14]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_123 BR32_2/C[4] sky130_fd_sc_hd__clkbuf_4_1/X BR32_2/C[3]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1704 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1715 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1726 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1737 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1748 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1759 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR32_2 BR32_2/C[31] BR64_3/C[30] BR64_3/C[29] BR64_3/C[28] BR64_3/C[27] BR64_3/C[26]
+ BR64_3/C[25] BR64_3/C[24] BR64_3/C[23] BR64_3/C[22] BR64_3/C[21] BR64_3/C[20] BR64_3/C[19]
+ BR64_3/C[18] BR64_3/C[17] BR32_2/C[16] BR32_2/C[15] BR32_2/C[14] BR32_2/C[13] BR64_3/C[12]
+ BR64_3/C[11] BR64_3/C[10] BR64_3/C[9] BR64_3/C[8] BR64_3/C[7] BR64_3/C[6] BR32_2/C[5]
+ BR32_2/C[4] BR32_2/C[3] BR64_3/C[2] BR64_3/C[1] BR64_3/C[0] vssd1 vccd1 BR32_2/RESET
+ BR32_2/OUT BR32
Xsky130_fd_sc_hd__decap_12_502 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_513 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_524 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_535 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_546 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_568 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_579 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1501 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1512 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1523 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1534 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1545 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1556 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1567 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1578 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1589 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o22ai_1_1 sky130_fd_sc_hd__o22ai_1_1/A2 sky130_fd_sc_hd__nand2_1_2/B
+ sky130_fd_sc_hd__o22ai_1_1/Y puf_sel0 sky130_fd_sc_hd__o22ai_1_1/B2 vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkbuf_4_6 BR64_3/C[52] BR64_1/C[52] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_310 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_321 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_332 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_343 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_354 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_365 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_376 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_387 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_398 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1320 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1331 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1342 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1353 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1364 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1375 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1386 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1397 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_0 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_5/A sky130_fd_sc_hd__o22ai_1_5/Y
+ sky130_fd_sc_hd__nand2_1_9/Y sky130_fd_sc_hd__o21ai_1_0/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_140 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_151 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_162 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_173 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_184 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_14 BR64_3/RESET sky130_fd_sc_hd__nor2_1_5/Y sky130_fd_sc_hd__nand2_1_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_195 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1150 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1161 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1172 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1183 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1194 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_6 vccd1 vssd1 BR128_3/C[74] sky130_fd_sc_hd__buf_6_6/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__decap_12_909 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_12 BR128_2/C[115] sky130_fd_sc_hd__clkbuf_4_1/X BR128_3/C[114]
+ sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_23 BR128_1/C[104] sky130_fd_sc_hd__clkbuf_4_1/A BR128_1/C[103]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_34 BR128_1/C[93] sky130_fd_sc_hd__clkbuf_4_1/A BR128_1/C[92]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_45 BR128_0/C[82] sky130_fd_sc_hd__clkbuf_4_1/X BR128_0/C[81]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_56 sky130_fd_sc_hd__dfrtp_2_56/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_3/C[70] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_67 BR64_1/C[60] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[59]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_78 BR64_1/C[49] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[48]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_89 BR64_1/C[38] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[37]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkbuf_4_70 BR128_3/C[84] BR128_0/C[84] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_706 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_717 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_728 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_739 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_102 BR64_1/C[25] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[24]
+ sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_113 BR32_2/C[14] sky130_fd_sc_hd__clkbuf_4_1/A BR32_2/C[13]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_124 BR32_2/C[3] sky130_fd_sc_hd__clkbuf_4_1/X sky130_fd_sc_hd__buf_6_8/A
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1705 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1716 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1727 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1738 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1749 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_0 vccd1 vssd1 BR128_3/C[69] BR128_2/C[69] vssd1 vccd1 sky130_fd_sc_hd__buf_2
XBR32_3 BR64_3/C[31] BR64_3/C[30] BR64_3/C[29] BR64_3/C[28] BR64_3/C[27] BR64_3/C[26]
+ BR64_3/C[25] BR64_3/C[24] BR64_3/C[23] BR64_3/C[22] BR64_3/C[21] BR64_3/C[20] BR64_3/C[19]
+ BR64_3/C[18] BR64_3/C[17] BR64_3/C[16] BR64_3/C[15] BR32_3/C[14] BR64_3/C[13] BR64_3/C[12]
+ BR64_3/C[11] BR64_3/C[10] BR64_3/C[9] BR64_3/C[8] BR64_3/C[7] BR64_3/C[6] BR64_3/C[5]
+ BR64_3/C[4] BR64_3/C[3] BR64_3/C[2] BR64_3/C[1] BR64_3/C[0] vssd1 vccd1 BR32_3/RESET
+ BR32_3/OUT BR32
Xsky130_fd_sc_hd__decap_12_503 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_514 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_525 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_536 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_547 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_558 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_569 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1502 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1513 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1524 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1535 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1546 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1568 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1579 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o22ai_1_2 sky130_fd_sc_hd__o21ai_1_1/Y sky130_fd_sc_hd__nand2_1_2/B
+ sky130_fd_sc_hd__o22ai_1_2/Y puf_sel0 sky130_fd_sc_hd__o21ai_1_0/Y vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkbuf_4_7 BR64_3/C[50] BR64_1/C[50] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_300 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_311 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_322 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_333 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_344 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_355 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_366 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_377 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_388 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_399 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1310 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1321 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1332 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1343 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1354 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1365 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1376 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1387 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1398 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o21ai_1_1 vssd1 vccd1 sky130_fd_sc_hd__nor2_1_5/A sky130_fd_sc_hd__o22ai_1_6/Y
+ sky130_fd_sc_hd__o21ai_1_1/B1 sky130_fd_sc_hd__o21ai_1_1/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_12_130 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_141 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_152 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_163 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_174 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_185 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_196 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1140 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1151 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1162 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1173 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1184 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1195 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_7 vccd1 vssd1 BR128_3/C[89] sky130_fd_sc_hd__buf_6_7/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__dfrtp_2_13 sky130_fd_sc_hd__dfrtp_2_13/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_3/C[113] sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_24 BR128_1/C[103] rstn BR128_1/C[102] sky130_fd_sc_hd__clkinv_8_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_35 BR128_1/C[92] sky130_fd_sc_hd__clkbuf_4_1/A BR128_3/C[91]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_46 BR128_0/C[81] sky130_fd_sc_hd__clkbuf_4_1/X BR128_0/C[80]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_57 sky130_fd_sc_hd__dfrtp_2_57/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_1/C[69] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_68 BR64_1/C[59] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[58]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_79 BR64_1/C[48] sky130_fd_sc_hd__clkbuf_4_1/X BR64_3/C[47]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkbuf_4_60 BR64_1/C[16] BR32_2/C[16] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_71 BR128_3/C[86] BR128_0/C[86] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_707 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_718 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_729 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_103 BR64_1/C[24] sky130_fd_sc_hd__clkbuf_4_1/A BR64_3/C[23]
+ sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_114 BR32_2/C[13] sky130_fd_sc_hd__clkbuf_4_1/A BR32_1/C[12]
+ sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_125 sky130_fd_sc_hd__buf_6_8/A sky130_fd_sc_hd__clkbuf_4_1/X
+ BR64_3/C[1] sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1706 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1717 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1728 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1739 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_1 vccd1 vssd1 BR128_3/C[68] BR128_2/C[68] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_504 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_515 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_526 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_537 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_548 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_559 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1503 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1514 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1525 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1536 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1547 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1558 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1569 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o22ai_1_3 BR32_0/OUT sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__o22ai_1_3/Y
+ length0 BR64_0/OUT vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkbuf_4_8 BR64_3/C[49] BR64_1/C[49] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_301 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_312 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_323 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_334 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_345 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_356 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_367 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_378 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_389 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1300 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1311 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1322 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1333 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1344 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1355 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1366 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1377 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1388 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1399 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_890 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_120 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_131 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_142 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_153 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_164 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_175 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_186 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_197 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1130 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1141 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1152 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1163 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1174 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1185 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1196 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_8 vccd1 vssd1 BR64_3/C[2] sky130_fd_sc_hd__buf_6_8/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__dfrtp_2_14 BR128_0/C[113] sky130_fd_sc_hd__clkbuf_4_1/X BR128_3/C[112]
+ sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_25 BR128_1/C[102] rstn BR128_1/C[101] sky130_fd_sc_hd__clkinv_8_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_36 sky130_fd_sc_hd__dfrtp_2_36/Q sky130_fd_sc_hd__clkbuf_4_1/A
+ BR128_3/C[90] sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_47 BR128_0/C[80] sky130_fd_sc_hd__clkbuf_4_1/X BR128_0/C[79]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_58 BR128_1/C[69] sky130_fd_sc_hd__clkbuf_4_1/X BR128_2/C[68]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_69 BR64_1/C[58] sky130_fd_sc_hd__clkbuf_4_1/X BR64_1/C[57]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkbuf_4_50 BR64_3/C[38] BR64_1/C[38] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_61 BR64_3/C[16] BR32_2/C[16] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_72 BR128_3/C[76] BR128_0/C[76] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_708 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_719 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_104 sky130_fd_sc_hd__buf_6_3/A sky130_fd_sc_hd__clkbuf_4_1/A
+ BR64_3/C[22] sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_115 BR32_1/C[12] sky130_fd_sc_hd__clkbuf_4_1/A BR64_3/C[11]
+ sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_126 BR32_1/C[1] sky130_fd_sc_hd__clkbuf_4_1/X BR64_3/C[0]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1707 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1718 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1729 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_2 vccd1 vssd1 BR128_3/C[113] BR128_0/C[113] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_505 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_516 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_527 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_538 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_549 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1504 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1515 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1526 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1537 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1548 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1559 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o22ai_1_4 BR32_1/OUT sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__o22ai_1_4/Y
+ sky130_fd_sc_hd__nand2_1_8/A BR64_1/OUT vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__clkbuf_4_9 BR64_3/C[41] BR64_1/C[41] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_302 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_313 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_324 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_335 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_346 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_357 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_368 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_379 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1301 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1312 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1323 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1334 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1345 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1356 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1367 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1378 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1389 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_880 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_891 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_110 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_121 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_132 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_143 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_154 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_165 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_176 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_187 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_198 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1120 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1131 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1142 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1153 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1164 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1175 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1186 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1197 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_0 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_6_9 vccd1 vssd1 BR128_3/C[77] sky130_fd_sc_hd__buf_6_9/A vssd1
+ vccd1 sky130_fd_sc_hd__buf_6
Xsky130_fd_sc_hd__dfrtp_2_15 sky130_fd_sc_hd__dfrtp_2_15/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_0/C[111] sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_26 BR128_1/C[101] rstn BR128_1/C[100] sky130_fd_sc_hd__clkinv_8_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_37 sky130_fd_sc_hd__dfrtp_2_37/Q sky130_fd_sc_hd__clkbuf_4_1/A
+ BR128_3/C[89] sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_48 BR128_0/C[79] sky130_fd_sc_hd__clkbuf_4_1/X BR128_3/C[78]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_59 BR128_2/C[68] sky130_fd_sc_hd__clkbuf_4_1/X BR128_2/C[67]
+ sky130_fd_sc_hd__clkinv_8_6/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkbuf_4_40 sky130_fd_sc_hd__nand2_1_8/A length0 vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_51 BR64_3/C[37] BR64_1/C[37] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_62 BR64_1/C[15] BR32_2/C[15] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_73 BR128_3/C[87] BR128_0/C[87] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_709 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_105 BR64_1/C[22] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[21]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_116 sky130_fd_sc_hd__clkbuf_8_0/A sky130_fd_sc_hd__clkbuf_4_1/A
+ BR64_3/C[10] sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_127 BR32_1/C[0] sky130_fd_sc_hd__clkbuf_4_1/X si sky130_fd_sc_hd__clkinv_8_7/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1708 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1719 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_3 vccd1 vssd1 so BR128_1/C[127] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_506 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_517 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_528 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_539 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1505 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1516 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1527 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1538 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1549 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o22ai_1_5 BR32_2/OUT sky130_fd_sc_hd__o22ai_1_5/B1 sky130_fd_sc_hd__o22ai_1_5/Y
+ sky130_fd_sc_hd__nand2_1_8/A BR64_2/OUT vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__decap_12_303 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_314 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_325 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_336 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_347 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_358 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_369 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1302 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1313 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1324 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1335 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1346 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1357 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1368 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1379 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_870 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_881 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_892 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_100 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_111 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_122 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_133 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_144 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_155 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_166 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_177 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_188 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_199 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1110 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1121 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1132 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1143 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1154 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1165 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1176 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1187 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1198 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_16 BR128_0/C[111] sky130_fd_sc_hd__clkbuf_4_1/X BR128_1/C[110]
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_27 BR128_1/C[100] rstn BR128_1/C[99] sky130_fd_sc_hd__clkinv_8_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_38 sky130_fd_sc_hd__buf_6_7/A sky130_fd_sc_hd__clkbuf_4_1/A
+ BR128_0/C[88] sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_49 BR128_0/C[78] sky130_fd_sc_hd__clkbuf_4_1/X sky130_fd_sc_hd__buf_6_9/A
+ sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkbuf_4_30 BR64_1/C[17] sky130_fd_sc_hd__dfrtp_2_110/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_41 BR64_3/C[57] BR64_1/C[57] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_52 BR64_3/C[35] BR64_1/C[35] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_63 BR64_3/C[15] BR32_2/C[15] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_74 BR128_3/C[88] BR128_0/C[88] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__dfrtp_2_106 BR64_1/C[21] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[20]
+ sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_117 sky130_fd_sc_hd__buf_12_0/A sky130_fd_sc_hd__clkbuf_4_1/A
+ BR32_1/C[9] sky130_fd_sc_hd__clkinv_8_3/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1709 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_4 vccd1 vssd1 BR128_3/C[111] BR128_0/C[111] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_507 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_518 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_529 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1506 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1517 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1528 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1539 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__o22ai_1_6 BR32_3/OUT sky130_fd_sc_hd__o22ai_1_6/B1 sky130_fd_sc_hd__o22ai_1_6/Y
+ sky130_fd_sc_hd__nand2_1_8/A BR64_3/OUT vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1
Xsky130_fd_sc_hd__decap_12_304 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_315 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_326 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_337 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_348 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_359 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1303 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1314 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1325 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1336 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1347 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1358 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1369 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_860 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_871 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_882 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_893 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1870 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_101 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_112 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_123 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_134 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_145 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_156 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_167 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_178 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_189 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1100 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1111 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1122 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1133 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1144 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1155 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1166 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1177 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1188 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1199 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_690 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_17 BR128_1/C[110] sky130_fd_sc_hd__clkbuf_4_1/A BR128_1/C[109]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_28 BR128_1/C[99] rstn BR128_1/C[98] sky130_fd_sc_hd__clkinv_8_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_39 BR128_0/C[88] sky130_fd_sc_hd__clkbuf_4_1/A BR128_0/C[87]
+ sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkbuf_4_20 BR128_3/C[83] BR128_0/C[83] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_31 BR128_3/C[123] sky130_fd_sc_hd__dfrtp_2_4/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_42 BR64_3/C[54] BR64_1/C[54] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_53 BR64_3/C[32] BR64_1/C[32] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_64 BR64_3/C[14] BR64_1/C[14] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__dfrtp_2_107 BR64_1/C[20] sky130_fd_sc_hd__clkbuf_4_1/A BR64_1/C[19]
+ sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_118 BR32_1/C[9] sky130_fd_sc_hd__clkbuf_4_1/A BR64_3/C[8]
+ sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__buf_2_5 vccd1 vssd1 BR128_3/C[110] BR128_1/C[110] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_508 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_519 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1507 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1518 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1529 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_10 vssd1 vccd1 sky130_fd_sc_hd__o22ai_1_1/A2 sky130_fd_sc_hd__o21ai_2_0/Y
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_12_305 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_316 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_327 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_338 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_349 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1304 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1315 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1326 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1337 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1348 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1359 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_850 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_861 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_872 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_883 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_894 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1860 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1871 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_102 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_113 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_124 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_135 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_146 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_157 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_168 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_179 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1101 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1112 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1123 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1134 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1145 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1156 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1167 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1178 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1189 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_680 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_691 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR128_0 BR128_0/RESET vccd1 BR64_3/C[0] BR64_3/C[1] BR64_3/C[2] BR64_3/C[3] BR64_3/C[4]
+ BR64_3/C[5] BR64_3/C[7] BR64_3/C[8] BR64_3/C[9] BR64_3/C[10] BR64_3/C[11] BR64_3/C[12]
+ BR64_3/C[13] BR64_1/C[14] BR64_1/C[15] BR64_1/C[16] BR64_1/C[17] BR64_1/C[18] BR64_1/C[19]
+ BR64_1/C[20] BR64_1/C[21] BR64_1/C[22] BR64_3/C[23] BR64_1/C[24] BR64_1/C[25] BR64_3/C[26]
+ BR64_1/C[27] BR64_1/C[28] BR64_1/C[29] BR64_1/C[30] BR64_3/C[6] BR64_3/C[31] BR64_1/C[32]
+ BR64_1/C[33] BR64_1/C[34] BR64_1/C[35] BR64_1/C[36] BR64_1/C[37] BR64_1/C[38] BR64_1/C[39]
+ BR64_1/C[40] BR64_1/C[41] BR64_1/C[42] BR64_1/C[43] BR64_3/C[44] BR64_1/C[45] BR64_1/C[46]
+ BR64_1/C[47] BR64_1/C[48] BR64_1/C[49] BR64_1/C[50] BR64_1/C[51] BR64_1/C[52] BR64_1/C[53]
+ BR64_1/C[54] BR64_1/C[55] BR64_1/C[56] BR64_1/C[57] BR64_1/C[58] BR64_1/C[59] BR64_1/C[60]
+ BR64_1/C[61] BR64_1/C[62] BR128_1/C[95] BR128_1/C[96] BR128_1/C[97] BR128_1/C[98]
+ BR128_1/C[99] BR128_1/C[100] BR128_1/C[101] BR128_1/C[102] BR128_1/C[103] BR128_1/C[104]
+ BR128_1/C[105] BR128_1/C[106] BR128_1/C[107] BR128_1/C[108] BR128_1/C[109] BR128_1/C[110]
+ BR128_0/C[111] BR128_3/C[112] BR128_0/C[113] BR128_3/C[114] BR128_2/C[115] BR128_2/C[116]
+ BR128_2/C[117] BR128_2/C[118] BR128_3/C[119] BR128_3/C[120] BR128_2/C[121] BR128_3/C[122]
+ BR128_3/C[123] BR128_3/C[124] BR128_2/C[125] BR128_2/C[126] BR128_1/C[127] BR64_1/C[63]
+ BR128_1/C[64] BR128_1/C[65] BR128_2/C[66] BR128_2/C[67] BR128_2/C[68] BR128_1/C[69]
+ BR128_3/C[70] BR128_3/C[71] BR128_3/C[72] BR128_3/C[73] BR128_3/C[74] BR128_3/C[75]
+ BR128_0/C[76] BR128_3/C[77] BR128_0/C[78] BR128_0/C[79] BR128_0/C[80] BR128_0/C[81]
+ BR128_0/C[82] BR128_0/C[83] BR128_0/C[84] BR128_0/C[85] BR128_0/C[86] BR128_0/C[87]
+ BR128_0/C[88] BR128_3/C[89] BR128_3/C[90] BR128_3/C[91] BR128_1/C[92] BR128_1/C[93]
+ BR128_1/C[94] BR128_0/OUT vssd1 BR128
Xsky130_fd_sc_hd__decap_12_1690 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_0 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__diode_2_0 BR128_3/OUT vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__dfrtp_2_18 BR128_1/C[109] sky130_fd_sc_hd__clkbuf_4_1/A BR128_1/C[108]
+ sky130_fd_sc_hd__clkinv_8_2/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_29 BR128_1/C[98] rstn BR128_1/C[97] sky130_fd_sc_hd__clkinv_8_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkbuf_4_10 BR64_3/C[40] BR64_1/C[40] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_21 BR128_3/C[78] BR128_0/C[78] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_32 BR128_3/C[124] sky130_fd_sc_hd__dfrtp_2_3/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_43 BR64_3/C[51] BR64_1/C[51] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_54 BR64_3/C[29] BR64_1/C[29] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_65 sky130_fd_sc_hd__o22ai_1_1/B2 sky130_fd_sc_hd__o21ai_0_0/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__dfrtp_2_108 sky130_fd_sc_hd__dfrtp_2_108/Q sky130_fd_sc_hd__clkbuf_4_1/A
+ BR64_1/C[18] sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__dfrtp_2_119 sky130_fd_sc_hd__clkbuf_8_1/A sky130_fd_sc_hd__clkbuf_4_1/A
+ BR64_3/C[7] sky130_fd_sc_hd__clkinv_8_4/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__buf_2_6 vccd1 vssd1 BR128_3/C[109] BR128_1/C[109] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_509 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1508 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1519 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_11 vssd1 vccd1 out sky130_fd_sc_hd__o22ai_1_0/Y vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_0 sky130_fd_sc_hd__buf_12_0/A BR64_3/C[10] vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_306 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_317 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_328 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_339 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1305 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1316 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1327 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1338 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1349 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_840 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_851 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_862 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_873 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_884 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_895 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1850 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1861 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1872 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_103 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_114 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_125 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_136 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_147 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_158 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_169 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1102 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1113 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1124 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1135 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1146 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1157 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1168 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1179 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_670 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_681 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_692 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR128_1 BR128_1/RESET vccd1 BR64_3/C[0] BR64_3/C[1] BR64_3/C[2] BR64_3/C[3] BR64_3/C[4]
+ BR64_3/C[5] BR64_3/C[7] BR64_3/C[8] BR64_3/C[9] BR64_3/C[10] BR64_3/C[11] BR64_3/C[12]
+ BR64_3/C[13] BR64_3/C[14] BR32_2/C[15] BR32_2/C[16] BR64_1/C[17] BR64_1/C[18] BR64_1/C[19]
+ BR64_3/C[20] BR64_3/C[21] BR64_3/C[22] BR64_3/C[23] BR64_3/C[24] BR64_3/C[25] BR64_3/C[26]
+ BR64_3/C[27] BR64_3/C[28] BR64_3/C[29] BR64_3/C[30] BR64_3/C[6] BR64_3/C[31] BR64_3/C[32]
+ BR64_1/C[33] BR64_3/C[34] BR64_3/C[35] BR64_3/C[36] BR64_3/C[37] BR64_3/C[38] BR64_3/C[39]
+ BR64_3/C[40] BR64_3/C[41] BR64_3/C[42] BR64_3/C[43] BR64_3/C[44] BR64_3/C[45] BR64_3/C[46]
+ BR64_3/C[47] BR128_1/C[48] BR64_3/C[49] BR64_3/C[50] BR64_3/C[51] BR64_3/C[52] BR64_3/C[53]
+ BR64_3/C[54] BR64_3/C[55] BR64_3/C[56] BR64_3/C[57] BR64_1/C[58] BR64_1/C[59] BR64_3/C[60]
+ BR64_1/C[61] BR64_1/C[62] BR128_1/C[95] BR128_1/C[96] BR128_1/C[97] BR128_1/C[98]
+ BR128_1/C[99] BR128_1/C[100] BR128_1/C[101] BR128_1/C[102] BR128_1/C[103] BR128_1/C[104]
+ BR128_1/C[105] BR128_1/C[106] BR128_1/C[107] BR128_1/C[108] BR128_1/C[109] BR128_1/C[110]
+ BR128_3/C[111] BR128_3/C[112] BR128_3/C[113] BR128_3/C[114] BR128_2/C[115] BR128_2/C[116]
+ BR128_2/C[117] BR128_2/C[118] BR128_3/C[119] BR128_3/C[120] BR128_2/C[121] BR128_3/C[122]
+ BR128_3/C[123] BR128_3/C[124] BR128_2/C[125] BR128_2/C[126] BR128_1/C[127] BR64_1/C[63]
+ BR128_1/C[64] BR128_1/C[65] BR128_2/C[66] BR128_2/C[67] BR128_2/C[68] BR128_1/C[69]
+ BR128_3/C[70] BR128_3/C[71] BR128_3/C[72] BR128_3/C[73] BR128_3/C[74] BR128_3/C[75]
+ BR128_3/C[76] BR128_3/C[77] BR128_3/C[78] BR128_3/C[79] BR128_3/C[80] BR128_3/C[81]
+ BR128_3/C[82] BR128_3/C[83] BR128_3/C[84] BR128_3/C[85] BR128_3/C[86] BR128_3/C[87]
+ BR128_3/C[88] BR128_3/C[89] BR128_3/C[90] BR128_3/C[91] BR128_1/C[92] BR128_1/C[93]
+ BR128_1/C[94] BR128_1/OUT vssd1 BR128
Xsky130_fd_sc_hd__decap_12_1680 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1691 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_4 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__diode_2_1 BR128_2/C[66] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__dfrtp_2_19 BR128_1/C[108] rstn BR128_1/C[107] sky130_fd_sc_hd__clkinv_8_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__clkbuf_4_11 BR64_3/C[36] BR64_1/C[36] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_22 BR128_3/C[85] BR128_0/C[85] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_33 BR128_3/C[119] sky130_fd_sc_hd__dfrtp_2_8/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_44 BR64_3/C[48] BR128_1/C[48] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_55 BR64_3/C[21] BR64_1/C[21] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_66 BR128_3/C[80] BR128_0/C[80] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__dfrtp_2_109 sky130_fd_sc_hd__dfrtp_2_109/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR64_1/C[17] sky130_fd_sc_hd__clkinv_8_7/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__buf_2_7 vccd1 vssd1 BR128_3/C[108] BR128_1/C[108] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_1509 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_12 vssd1 vccd1 BR128_1/C[48] BR64_1/C[48] vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_1 sky130_fd_sc_hd__buf_12_1/A BR64_3/C[7] vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_307 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_318 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_329 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1306 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1317 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1328 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1339 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_830 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_841 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_852 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_863 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_874 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_885 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_896 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1840 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1851 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1862 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1873 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_0 BR128_1/C[127] sky130_fd_sc_hd__clkbuf_4_1/X BR128_2/C[126]
+ sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_104 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_115 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_126 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_137 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_148 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_159 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1103 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1114 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1125 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1136 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1147 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1158 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1169 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_660 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_671 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_682 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_693 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1670 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR128_2 BR128_2/RESET vccd1 BR64_3/C[0] BR64_3/C[1] BR64_3/C[2] BR64_3/C[3] BR64_3/C[4]
+ BR64_3/C[5] BR64_3/C[7] BR64_3/C[8] BR64_3/C[9] BR64_3/C[10] BR64_3/C[11] BR64_3/C[12]
+ BR64_3/C[13] BR64_3/C[14] BR64_3/C[15] BR64_3/C[16] BR64_3/C[17] BR64_3/C[18] BR64_3/C[19]
+ BR64_3/C[20] BR64_3/C[21] BR64_3/C[22] BR64_3/C[23] BR64_3/C[24] BR64_3/C[25] BR64_3/C[26]
+ BR64_3/C[27] BR64_3/C[28] BR64_3/C[29] BR64_3/C[30] BR64_3/C[6] BR64_3/C[31] BR64_3/C[32]
+ BR64_3/C[33] BR64_3/C[34] BR64_3/C[35] BR64_3/C[36] BR64_3/C[37] BR64_3/C[38] BR64_3/C[39]
+ BR64_3/C[40] BR64_3/C[41] BR64_3/C[42] BR64_3/C[43] BR64_3/C[44] BR64_3/C[45] BR64_3/C[46]
+ BR64_3/C[47] BR64_3/C[48] BR64_3/C[49] BR64_3/C[50] BR64_3/C[51] BR64_3/C[52] BR64_3/C[53]
+ BR64_3/C[54] BR64_3/C[55] BR64_3/C[56] BR64_3/C[57] BR64_3/C[58] BR64_3/C[59] BR64_3/C[60]
+ BR64_3/C[61] BR64_3/C[62] BR128_3/C[95] BR128_3/C[96] BR128_3/C[97] BR128_3/C[98]
+ BR128_3/C[99] BR128_3/C[100] BR128_3/C[101] BR128_3/C[102] BR128_3/C[103] BR128_3/C[104]
+ BR128_3/C[105] BR128_3/C[106] BR128_3/C[107] BR128_3/C[108] BR128_3/C[109] BR128_3/C[110]
+ BR128_3/C[111] BR128_3/C[112] BR128_3/C[113] BR128_3/C[114] BR128_2/C[115] BR128_2/C[116]
+ BR128_2/C[117] BR128_2/C[118] BR128_3/C[119] BR128_3/C[120] BR128_2/C[121] BR128_3/C[122]
+ BR128_3/C[123] BR128_3/C[124] BR128_2/C[125] BR128_2/C[126] so BR64_3/C[63] BR128_3/C[64]
+ BR128_3/C[65] BR128_2/C[66] BR128_2/C[67] BR128_2/C[68] BR128_2/C[69] BR128_3/C[70]
+ BR128_3/C[71] BR128_3/C[72] BR128_3/C[73] BR128_3/C[74] BR128_3/C[75] BR128_3/C[76]
+ BR128_3/C[77] BR128_3/C[78] BR128_3/C[79] BR128_3/C[80] BR128_3/C[81] BR128_3/C[82]
+ BR128_3/C[83] BR128_3/C[84] BR128_3/C[85] BR128_3/C[86] BR128_3/C[87] BR128_3/C[88]
+ BR128_3/C[89] BR128_3/C[90] BR128_3/C[91] BR128_3/C[92] BR128_3/C[93] BR128_3/C[94]
+ BR128_2/OUT vssd1 BR128
Xsky130_fd_sc_hd__decap_12_1681 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1692 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_5 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_490 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__diode_2_2 BR128_3/C[120] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkbuf_4_12 BR64_3/C[34] BR64_1/C[34] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_23 BR128_3/C[73] sky130_fd_sc_hd__dfrtp_2_54/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_34 BR128_3/C[112] sky130_fd_sc_hd__dfrtp_2_15/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_45 BR64_3/C[46] BR64_1/C[46] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_56 BR64_3/C[20] BR64_1/C[20] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_67 BR64_3/C[24] BR64_1/C[24] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__buf_2_8 vccd1 vssd1 BR128_3/C[107] BR128_1/C[107] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__clkbuf_1_13 vssd1 vccd1 BR128_2/C[69] BR128_1/C[69] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__buf_12_2 BR32_1/C[12] BR64_3/C[12] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__buf_12
Xsky130_fd_sc_hd__decap_12_308 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_319 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1307 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1318 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1329 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_820 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_831 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_842 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_853 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_864 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_875 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_886 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_897 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1830 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1841 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1852 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1863 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1874 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_1 BR128_2/C[126] sky130_fd_sc_hd__clkbuf_4_1/X BR128_2/C[125]
+ sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_105 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_116 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_127 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_138 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_149 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1104 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1115 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1126 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1137 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1148 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1159 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_650 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_661 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_672 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_683 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_694 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1660 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1671 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XBR128_3 BR128_3/RESET vccd1 BR64_3/C[0] BR64_3/C[1] BR64_3/C[2] BR64_3/C[3] BR64_3/C[4]
+ BR64_3/C[5] BR64_3/C[7] BR64_3/C[8] BR64_3/C[9] BR64_3/C[10] BR64_3/C[11] BR64_3/C[12]
+ BR64_3/C[13] BR64_3/C[14] BR64_3/C[15] BR64_3/C[16] BR64_3/C[17] BR64_3/C[18] BR64_3/C[19]
+ BR64_3/C[20] BR64_3/C[21] BR64_3/C[22] BR64_3/C[23] BR64_3/C[24] BR64_3/C[25] BR64_3/C[26]
+ BR64_3/C[27] BR64_3/C[28] BR64_3/C[29] BR64_3/C[30] BR64_3/C[6] BR64_3/C[31] BR64_3/C[32]
+ BR64_3/C[33] BR64_3/C[34] BR64_3/C[35] BR64_3/C[36] BR64_3/C[37] BR64_3/C[38] BR64_3/C[39]
+ BR64_3/C[40] BR64_3/C[41] BR64_3/C[42] BR64_3/C[43] BR64_3/C[44] BR64_3/C[45] BR64_3/C[46]
+ BR64_3/C[47] BR64_3/C[48] BR64_3/C[49] BR64_3/C[50] BR64_3/C[51] BR64_3/C[52] BR64_3/C[53]
+ BR64_3/C[54] BR64_3/C[55] BR64_3/C[56] BR64_3/C[57] BR64_3/C[58] BR64_3/C[59] BR64_3/C[60]
+ BR64_3/C[61] BR64_3/C[62] BR128_3/C[95] BR128_3/C[96] BR128_3/C[97] BR128_3/C[98]
+ BR128_3/C[99] BR128_3/C[100] BR128_3/C[101] BR128_3/C[102] BR128_3/C[103] BR128_3/C[104]
+ BR128_3/C[105] BR128_3/C[106] BR128_3/C[107] BR128_3/C[108] BR128_3/C[109] BR128_3/C[110]
+ BR128_3/C[111] BR128_3/C[112] BR128_3/C[113] BR128_3/C[114] BR128_3/C[115] BR128_3/C[116]
+ BR128_3/C[117] BR128_3/C[118] BR128_3/C[119] BR128_3/C[120] BR128_3/C[121] BR128_3/C[122]
+ BR128_3/C[123] BR128_3/C[124] BR128_3/C[125] BR128_3/C[126] so BR64_3/C[63] BR128_3/C[64]
+ BR128_3/C[65] BR128_3/C[66] BR128_3/C[67] BR128_3/C[68] BR128_3/C[69] BR128_3/C[70]
+ BR128_3/C[71] BR128_3/C[72] BR128_3/C[73] BR128_3/C[74] BR128_3/C[75] BR128_3/C[76]
+ BR128_3/C[77] BR128_3/C[78] BR128_3/C[79] BR128_3/C[80] BR128_3/C[81] BR128_3/C[82]
+ BR128_3/C[83] BR128_3/C[84] BR128_3/C[85] BR128_3/C[86] BR128_3/C[87] BR128_3/C[88]
+ BR128_3/C[89] BR128_3/C[90] BR128_3/C[91] BR128_3/C[92] BR128_3/C[93] BR128_3/C[94]
+ BR128_3/OUT vssd1 BR128
Xsky130_fd_sc_hd__decap_12_1682 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1693 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_6 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_480 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_491 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1490 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_30 vccd1 vssd1 BR64_3/C[58] BR64_1/C[58] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_3 BR64_3/C[6] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkbuf_4_13 BR64_3/C[30] BR64_1/C[30] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_24 BR128_3/C[90] sky130_fd_sc_hd__dfrtp_2_37/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_35 BR64_1/C[19] sky130_fd_sc_hd__dfrtp_2_108/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_46 BR64_3/C[45] BR64_1/C[45] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_57 BR64_3/C[19] BR64_1/C[19] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_68 BR128_3/C[79] BR128_0/C[79] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_6_0 vccd1 vssd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__buf_2_9 vccd1 vssd1 BR128_3/C[106] BR128_1/C[106] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_309 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1308 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1319 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_810 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_821 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_832 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_843 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_854 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_865 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_876 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_887 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_898 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1820 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1831 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1842 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1853 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1864 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1875 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_2 BR128_2/C[125] sky130_fd_sc_hd__clkbuf_4_1/X BR128_3/C[124]
+ sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_106 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_117 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_128 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_139 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1105 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1116 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1127 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1138 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1149 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_640 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_651 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_662 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_684 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_695 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1650 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1661 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1672 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1683 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1694 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_7 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_470 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_481 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_492 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1480 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1491 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_20 vccd1 vssd1 BR128_3/C[95] BR128_1/C[95] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_31 vccd1 vssd1 BR64_3/C[33] BR64_1/C[33] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_4 BR64_3/C[6] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkbuf_4_14 BR64_3/C[28] BR64_1/C[28] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_25 BR64_1/C[18] sky130_fd_sc_hd__dfrtp_2_109/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_36 BR128_3/C[122] sky130_fd_sc_hd__dfrtp_2_5/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_47 BR64_3/C[43] BR64_1/C[43] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_58 BR64_3/C[18] BR64_1/C[18] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_69 BR128_3/C[81] BR128_0/C[81] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_1309 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_800 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_811 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_822 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_833 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_844 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_855 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_866 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_877 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_888 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_899 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1810 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1821 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1832 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1843 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1854 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1865 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1876 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_3 sky130_fd_sc_hd__dfrtp_2_3/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_3/C[123] sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_107 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_118 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_129 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1106 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1117 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1128 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1139 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_630 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_652 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_663 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_674 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_696 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1640 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1651 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1662 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1684 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1695 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_8 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_460 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_471 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_482 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_493 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1470 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1481 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1492 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_10 vccd1 vssd1 BR128_3/C[105] BR128_1/C[105] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_21 vccd1 vssd1 BR128_3/C[94] BR128_1/C[94] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_5 BR64_3/C[6] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkbuf_4_15 BR64_3/C[27] BR64_1/C[27] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_26 BR128_3/C[91] sky130_fd_sc_hd__dfrtp_2_36/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_37 BR128_3/C[114] sky130_fd_sc_hd__dfrtp_2_13/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_48 BR64_3/C[42] BR64_1/C[42] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_59 BR64_3/C[17] BR64_1/C[17] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_290 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_801 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_812 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_823 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_834 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_845 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_856 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_867 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_878 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_889 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1800 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1811 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1822 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1833 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1844 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1855 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1866 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1877 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_4 sky130_fd_sc_hd__dfrtp_2_4/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_3/C[122] sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_108 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_119 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1107 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1118 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1129 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_620 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_631 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_642 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_653 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_664 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_675 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_686 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1630 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1652 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1663 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1674 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1696 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_450 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_461 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_472 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_483 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_494 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1460 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1471 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1482 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1493 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_11 vccd1 vssd1 BR128_3/C[104] BR128_1/C[104] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_22 vccd1 vssd1 BR128_3/C[93] BR128_1/C[93] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_6 BR64_3/C[6] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkbuf_4_16 BR64_3/C[25] BR64_1/C[25] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_27 BR128_3/C[71] sky130_fd_sc_hd__dfrtp_2_56/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_38 BR128_3/C[120] sky130_fd_sc_hd__dfrtp_2_7/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_49 BR64_3/C[39] BR64_1/C[39] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_280 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_291 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1290 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2b_1_0 BR128_0/RESET sky130_fd_sc_hd__nor2_1_2/B length1 vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__decap_12_802 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_813 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_824 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_835 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_846 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_857 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_868 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_879 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1801 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1812 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1823 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1834 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1845 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1856 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1867 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1878 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_5 sky130_fd_sc_hd__dfrtp_2_5/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_2/C[121] sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_109 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1108 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1119 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_610 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_621 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_632 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_643 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_654 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_665 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_676 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_687 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_698 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1620 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1631 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1642 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1653 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1664 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1675 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1686 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_440 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_451 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_462 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_473 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_484 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_495 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1450 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1461 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1472 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1483 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1494 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_12 vccd1 vssd1 BR128_3/C[103] BR128_1/C[103] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_23 vccd1 vssd1 BR128_3/C[92] BR128_1/C[92] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_7 BR64_3/C[6] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkbuf_4_17 BR64_3/C[22] BR64_1/C[22] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_28 BR128_3/C[72] sky130_fd_sc_hd__dfrtp_2_55/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_39 sky130_fd_sc_hd__nor2_1_5/A length1 vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_270 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_281 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_292 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1280 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1291 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2b_1_1 BR128_1/RESET sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__decap_12_803 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_814 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_825 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_836 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_847 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_858 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_869 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1802 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1813 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1824 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1835 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1846 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1857 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1868 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1879 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_6 BR128_2/C[121] sky130_fd_sc_hd__clkbuf_4_1/X BR128_3/C[120]
+ sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_1109 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_600 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_611 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_622 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_633 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_644 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_655 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_666 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_677 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_688 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_699 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1610 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1621 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1632 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1643 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1654 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1665 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1676 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1687 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1698 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_430 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_441 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_452 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_463 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_474 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_485 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_496 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1440 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1451 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1462 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1473 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1484 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1495 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_13 vccd1 vssd1 BR128_3/C[102] BR128_1/C[102] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_24 vccd1 vssd1 BR128_3/C[65] BR128_1/C[65] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__diode_2_8 BR64_3/C[6] vssd1 vccd1 vccd1 vssd1 sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__clkbuf_4_18 BR64_1/C[14] BR32_2/C[14] vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_29 BR128_3/C[70] sky130_fd_sc_hd__dfrtp_2_57/Q vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_260 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_271 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_282 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_293 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1270 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1281 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1292 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2b_1_2 BR128_2/RESET sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__nor2_1_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__decap_12_804 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_815 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_826 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_837 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_848 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_859 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1803 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1814 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1825 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1836 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1847 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1858 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1869 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_7 sky130_fd_sc_hd__dfrtp_2_7/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_3/C[119] sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_612 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_623 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_634 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_656 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_667 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_678 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_689 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1600 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1611 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1622 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1633 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1644 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1655 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1666 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1677 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1688 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_0 sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__nand2_1_2/B
+ sky130_fd_sc_hd__nor2_1_0/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_1699 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_420 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_431 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_442 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_453 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_464 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_475 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_486 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_497 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1430 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1441 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1452 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1463 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1474 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1485 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1496 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_14 vccd1 vssd1 BR128_3/C[101] BR128_1/C[101] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_25 vccd1 vssd1 BR128_3/C[64] BR128_1/C[64] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__clkbuf_4_19 BR128_3/C[82] BR128_0/C[82] vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__decap_12_250 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_261 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_272 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_283 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_294 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1260 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1271 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1282 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1293 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2b_1_3 BR128_3/RESET sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__nor2_1_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2b_1
Xsky130_fd_sc_hd__decap_12_1090 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_805 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_816 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_827 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_838 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_849 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1804 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1815 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1826 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1837 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1848 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1859 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_8 sky130_fd_sc_hd__dfrtp_2_8/Q sky130_fd_sc_hd__clkbuf_4_1/X
+ BR128_2/C[118] sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_602 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_624 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_635 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_646 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_668 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_679 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1612 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1623 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1634 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1656 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1667 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1678 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1689 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_1 sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__nor2_1_0/Y
+ puf_sel0 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_90 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_410 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_421 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_432 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_443 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_454 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_465 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_476 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_487 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_498 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1420 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1431 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1442 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1453 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1464 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1475 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1486 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1497 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_15 vccd1 vssd1 BR128_3/C[100] BR128_1/C[100] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_26 vccd1 vssd1 BR64_3/C[63] BR64_1/C[63] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__o21ai_2_0 sky130_fd_sc_hd__nand2_1_6/Y sky130_fd_sc_hd__o21ai_2_0/Y
+ sky130_fd_sc_hd__nor2_1_5/A sky130_fd_sc_hd__o22ai_1_4/Y vssd1 vccd1 vssd1 vccd1
+ sky130_fd_sc_hd__o21ai_2
Xsky130_fd_sc_hd__decap_12_240 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_251 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_262 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_273 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_284 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_295 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1250 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1261 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1272 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1283 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1294 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_0 vssd1 vccd1 BR128_3/C[67] BR128_2/C[67] vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_0 sky130_fd_sc_hd__nand2_1_2/B puf_sel0 vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1080 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1091 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_806 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_817 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_828 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_839 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1805 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1816 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1827 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1838 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1849 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_2_9 BR128_2/C[118] sky130_fd_sc_hd__clkbuf_4_1/X BR128_2/C[117]
+ sky130_fd_sc_hd__clkinv_8_8/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__dfrtp_2
Xsky130_fd_sc_hd__decap_12_603 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_614 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_625 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_636 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_647 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_658 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1602 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1624 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1635 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1646 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1668 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1679 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_2 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nand2_1_2/B
+ sky130_fd_sc_hd__nor2_1_1/Y vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_80 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_91 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_400 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_411 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_422 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_433 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_444 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_455 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_466 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_477 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_488 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_499 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1410 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1421 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1432 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1443 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1454 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1465 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1476 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1487 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1498 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_16 vccd1 vssd1 BR128_3/C[99] BR128_1/C[99] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_27 vccd1 vssd1 BR64_3/C[62] BR64_1/C[62] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_230 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_241 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_252 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_263 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_274 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_285 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_296 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1240 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1251 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1262 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1273 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1284 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1295 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_1 vssd1 vccd1 BR128_3/C[66] BR128_2/C[66] vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_1 sky130_fd_sc_hd__nor2_1_1/B puf_sel1 vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1070 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1081 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1092 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_807 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_818 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_829 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1806 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1817 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1828 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1839 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_604 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_615 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_626 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_637 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_648 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_659 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1603 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1614 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1625 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1636 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1647 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1658 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_3 sky130_fd_sc_hd__nand2_1_3/Y BR128_0/OUT length1 vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_70 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_81 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_92 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_401 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_412 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_423 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_434 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_445 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_456 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_467 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_478 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_489 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1400 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1411 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1422 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1433 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1444 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1455 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1466 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1477 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1488 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1499 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_17 vccd1 vssd1 BR128_3/C[98] BR128_1/C[98] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_28 vccd1 vssd1 BR64_3/C[61] BR64_1/C[61] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_990 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_220 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_231 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_242 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_253 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_264 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_275 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_286 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_297 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1230 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1241 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1252 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1263 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1274 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1285 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1296 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_2 vssd1 vccd1 BR128_3/C[115] BR128_2/C[115] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_2 sky130_fd_sc_hd__nand2_1_4/B length0 vssd1 vccd1 vssd1
+ vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1060 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1071 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1082 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1093 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_808 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_819 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1807 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1818 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1829 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_605 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_616 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_627 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_638 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_649 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1604 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1615 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1626 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1637 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1648 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1659 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_4 BR32_0/RESET sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nor2_1_2/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_60 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_71 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_82 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_93 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_402 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_413 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_424 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_435 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_446 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_457 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_468 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_479 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1401 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1412 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1423 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1434 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1445 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1456 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1467 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1478 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1489 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_18 vccd1 vssd1 BR128_3/C[97] BR128_1/C[97] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_29 vccd1 vssd1 BR64_3/C[59] BR64_1/C[59] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_980 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_991 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_210 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_232 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_243 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_254 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_265 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_276 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_287 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_298 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1220 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1231 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1242 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1253 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1264 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1275 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1286 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1297 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_3 vssd1 vccd1 BR32_3/C[14] BR32_2/C[14] vssd1 vccd1 sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__o21ai_0_0 vssd1 vccd1 sky130_fd_sc_hd__o21ai_0_0/Y sky130_fd_sc_hd__nand2_1_3/Y
+ length1 sky130_fd_sc_hd__o22ai_1_3/Y vssd1 vccd1 sky130_fd_sc_hd__o21ai_0
Xsky130_fd_sc_hd__clkinv_1_3 sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__nand2_1_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1050 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1061 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1072 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1083 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1094 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_809 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1808 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1819 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_606 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_628 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_639 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1605 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1616 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1627 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1638 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1649 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_5 BR64_0/RESET sky130_fd_sc_hd__nor2_1_2/Y length0 vssd1
+ vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_50 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_61 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_72 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_83 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_94 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_403 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_414 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_425 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_436 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_447 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_458 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_469 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1402 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1413 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1424 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1435 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1446 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1457 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1468 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1479 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_19 vccd1 vssd1 BR128_3/C[96] BR128_1/C[96] vssd1 vccd1 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_970 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_981 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_992 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_200 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_211 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_222 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_233 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_244 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_255 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_266 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_277 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_288 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_299 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1210 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1232 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1243 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1254 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1265 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1276 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1287 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1298 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_4 vssd1 vccd1 BR128_3/C[116] BR128_2/C[116] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_4 sky130_fd_sc_hd__o22ai_1_5/B1 sky130_fd_sc_hd__nand2_1_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1040 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1051 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1062 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1073 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1084 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1095 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1809 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_607 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_618 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1606 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1628 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1639 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_6 sky130_fd_sc_hd__nand2_1_6/Y BR128_1/OUT sky130_fd_sc_hd__nor2_1_5/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_40 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_51 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_62 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_73 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_84 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_95 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_404 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_415 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_426 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_437 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_448 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_459 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1403 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1414 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1425 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1436 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1447 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1458 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1469 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_960 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_971 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_982 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_993 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_201 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_212 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_223 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_234 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_245 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_256 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_267 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_278 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_289 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1200 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1211 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1222 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1233 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1244 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1255 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1266 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1277 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1288 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1299 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_790 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_5 vssd1 vccd1 BR128_3/C[118] BR128_2/C[118] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_5 sky130_fd_sc_hd__o22ai_1_6/B1 sky130_fd_sc_hd__nand2_1_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1030 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1041 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1052 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1063 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1074 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1085 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1096 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_608 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_619 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1607 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1618 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_7 BR32_1/RESET sky130_fd_sc_hd__nand2_1_7/B sky130_fd_sc_hd__nor2_1_3/Y
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_30 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_41 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_52 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_63 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_74 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_85 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_96 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_405 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_416 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_427 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_438 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_449 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1404 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1415 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1426 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1437 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1448 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1459 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_950 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_961 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_972 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_983 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_994 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_202 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_213 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_224 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_235 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_246 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_257 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_268 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_279 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1201 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1212 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1223 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1234 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1245 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1256 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1267 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1278 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1289 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_780 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_791 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1790 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_6 vssd1 vccd1 BR128_3/C[125] BR128_2/C[125] vssd1 vccd1
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkinv_1_6 sky130_fd_sc_hd__clkinv_4_0/A BR32_2/C[31] vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_12_1020 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1031 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1042 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1053 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1064 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1075 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1086 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1097 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_609 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1608 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1619 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_1_8 BR64_1/RESET sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__nand2_1_8/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_12_20 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_31 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_42 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_53 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_64 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_75 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_86 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_97 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_406 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_417 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_428 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_439 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1405 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1416 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1427 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1438 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1449 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_940 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_951 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_962 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_973 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_984 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_995 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_8_0 BR64_3/C[11] sky130_fd_sc_hd__clkbuf_8_0/A vssd1 vccd1
+ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_8
Xsky130_fd_sc_hd__decap_12_203 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_214 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_225 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_236 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_247 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_258 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_269 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1202 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1213 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1224 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1235 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1246 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1257 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1268 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_1279 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkinv_8_0 sky130_fd_sc_hd__clkinv_8_5/A sky130_fd_sc_hd__clkinv_8_0/A
+ vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_12_770 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_781 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_792 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
.ends

.subckt sky130_fd_pr__res_generic_m1_DBNWX4 m1_n500_n557# m1_n500_500#
R0 m1_n500_n557# m1_n500_500# sky130_fd_pr__res_generic_m1 w=5e+06u l=5e+06u
.ends

.subckt puf_top m1_44147_10052# puf_super_0/si puf_super_0/length0 puf_super_0/out
+ puf_super_0/clk puf_super_0/reset puf_super_0/puf_sel0 puf_super_0/length1 puf_super_0/puf_sel1
+ puf_super_0/vccd1 puf_super_0/so m1_40740_16650# VSUBS puf_super_0/rstn
Xpuf_super_0 puf_super_0/reset puf_super_0/clk puf_super_0/si puf_super_0/puf_sel1
+ puf_super_0/puf_sel0 puf_super_0/length1 puf_super_0/length0 puf_super_0/out puf_super_0/so
+ puf_super_0/vccd1 puf_super_0/rstn VSUBS puf_super
Xsky130_fd_pr__res_generic_m1_DBNWX4_0 puf_super_0/so m1_40740_16650# sky130_fd_pr__res_generic_m1_DBNWX4
Xsky130_fd_pr__res_generic_m1_DBNWX4_1 puf_super_0/out m1_44147_10052# sky130_fd_pr__res_generic_m1_DBNWX4
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xpuf_top_0 la_data_out[0] io_in[20] io_in[18] io_out[25] io_in[21] io_in[26] io_in[23]
+ io_in[17] io_in[22] vccd2 io_out[24] la_data_out[1] vssd2 io_in[19] puf_top
.ends

