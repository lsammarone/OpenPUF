magic
tech sky130A
magscale 1 2
timestamp 1654748177
<< error_p >>
rect 137227 243593 138743 243859
rect 33429 117817 33487 117819
rect 33551 117817 33609 117819
rect 33673 117817 33731 117819
rect 33795 117817 33853 117819
rect 36757 80121 36811 80125
rect 36851 80121 36905 80125
rect 36945 80121 36999 80125
rect 36811 80069 36813 80121
rect 36905 80069 36907 80121
rect 36999 80069 37001 80121
rect 6441 4799 6443 4861
rect 6529 4799 6531 4861
rect 6615 4799 6617 4861
rect 6719 4799 6721 4861
rect 6823 4799 6825 4861
rect 6911 4799 6913 4861
<< error_s >>
rect 157159 377037 158995 377135
rect 156931 376709 158995 377037
rect 157159 376579 158995 376709
rect 159373 376579 159929 377135
rect 48953 206341 49509 208177
<< metal2 >>
rect 3305 382079 3759 382237
rect 3305 381971 3427 382079
rect 3649 381971 3759 382079
rect 3305 379301 3759 381971
rect 3305 379165 3481 379301
rect 3597 379165 3759 379301
rect 3305 379121 3759 379165
rect 43661 344377 44243 344460
rect 43661 344307 43703 344377
rect 43767 344307 43841 344377
rect 43905 344307 43979 344377
rect 44043 344307 44117 344377
rect 44181 344307 44243 344377
rect 43661 336159 44243 344307
rect 43661 336041 43739 336159
rect 43871 336041 43991 336159
rect 44123 336041 44243 336159
rect 43661 335969 44243 336041
rect 43661 335851 43739 335969
rect 43871 335851 43991 335969
rect 44123 335851 44243 335969
rect 43661 335753 44243 335851
rect 43363 306697 43967 306767
rect 43363 306585 43393 306697
rect 43453 306585 43525 306697
rect 43585 306585 43657 306697
rect 43717 306585 43789 306697
rect 43849 306585 43967 306697
rect 43363 292947 43967 306585
rect 43363 292707 43447 292947
rect 43619 292707 43725 292947
rect 43897 292707 43967 292947
rect 43363 292543 43967 292707
rect 42575 268903 43475 269281
rect 42575 268749 42645 268903
rect 42711 268749 42811 268903
rect 42877 268749 42977 268903
rect 43043 268749 43143 268903
rect 43209 268749 43309 268903
rect 43375 268749 43475 268903
rect 42575 250345 43475 268749
rect 42575 249445 43691 250345
rect 26048 231191 26774 231576
rect 26048 231043 26105 231191
rect 26199 231043 26271 231191
rect 26365 231043 26437 231191
rect 26531 231043 26603 231191
rect 26697 231043 26774 231191
rect 26048 122707 26774 231043
rect 27939 193395 28791 193697
rect 27939 193181 28009 193395
rect 28117 193181 28213 193395
rect 28321 193181 28417 193395
rect 28525 193181 28621 193395
rect 28729 193181 28791 193395
rect 25805 122391 26907 122707
rect 25805 122085 25899 122391
rect 26121 122085 26405 122391
rect 26627 122085 26907 122391
rect 25805 121981 26907 122085
rect 27939 79147 28791 193181
rect 27939 78783 28021 79147
rect 28185 78783 28307 79147
rect 28471 78783 28593 79147
rect 28757 78783 28791 79147
rect 27939 78703 28791 78783
rect 30243 155645 31045 155996
rect 30243 155563 30311 155645
rect 30399 155563 30513 155645
rect 30601 155563 30715 155645
rect 30803 155563 30917 155645
rect 31005 155563 31045 155645
rect 6147 42407 6895 42465
rect 6147 42341 6279 42407
rect 6363 42341 6459 42407
rect 6543 42341 6639 42407
rect 6723 42341 6895 42407
rect 6147 42229 6895 42341
rect 6365 5125 6601 42229
rect 30243 35831 31045 155563
rect 30243 35593 30329 35831
rect 30469 35593 30585 35831
rect 30725 35593 30841 35831
rect 30981 35593 31045 35831
rect 30243 35273 31045 35593
rect 33371 117817 33899 118389
rect 33371 117763 33429 117817
rect 33487 117763 33551 117817
rect 33609 117763 33673 117817
rect 33731 117763 33795 117817
rect 33853 117763 33899 117817
rect 33371 13415 33899 117763
rect 32801 13189 33899 13415
rect 32801 13057 32959 13189
rect 33105 13057 33293 13189
rect 33439 13057 33627 13189
rect 33773 13057 33899 13189
rect 32801 12887 33899 13057
rect 36721 80121 37057 80259
rect 36721 80069 36757 80121
rect 36811 80069 36851 80121
rect 36905 80069 36945 80121
rect 36999 80069 37057 80121
rect 36721 8547 37057 80069
rect 36355 8445 37449 8547
rect 36355 8339 36469 8445
rect 36599 8339 36727 8445
rect 36857 8339 36985 8445
rect 37115 8339 37449 8445
rect 36355 8211 37449 8339
rect 6331 4861 6953 5125
rect 6331 4799 6387 4861
rect 6441 4799 6475 4861
rect 6529 4799 6561 4861
rect 6615 4799 6665 4861
rect 6719 4799 6769 4861
rect 6823 4799 6857 4861
rect 6911 4799 6953 4861
rect 6331 4683 6953 4799
<< via2 >>
rect 3427 381971 3649 382079
rect 3481 379165 3597 379301
rect 43703 344307 43767 344377
rect 43841 344307 43905 344377
rect 43979 344307 44043 344377
rect 44117 344307 44181 344377
rect 43739 336041 43871 336159
rect 43991 336041 44123 336159
rect 43739 335851 43871 335969
rect 43991 335851 44123 335969
rect 43393 306585 43453 306697
rect 43525 306585 43585 306697
rect 43657 306585 43717 306697
rect 43789 306585 43849 306697
rect 43447 292707 43619 292947
rect 43725 292707 43897 292947
rect 42645 268749 42711 268903
rect 42811 268749 42877 268903
rect 42977 268749 43043 268903
rect 43143 268749 43209 268903
rect 43309 268749 43375 268903
rect 26105 231043 26199 231191
rect 26271 231043 26365 231191
rect 26437 231043 26531 231191
rect 26603 231043 26697 231191
rect 28009 193181 28117 193395
rect 28213 193181 28321 193395
rect 28417 193181 28525 193395
rect 28621 193181 28729 193395
rect 25899 122085 26121 122391
rect 26405 122085 26627 122391
rect 28021 78783 28185 79147
rect 28307 78783 28471 79147
rect 28593 78783 28757 79147
rect 30311 155563 30399 155645
rect 30513 155563 30601 155645
rect 30715 155563 30803 155645
rect 30917 155563 31005 155645
rect 6279 42341 6363 42407
rect 6459 42341 6543 42407
rect 6639 42341 6723 42407
rect 30329 35593 30469 35831
rect 30585 35593 30725 35831
rect 30841 35593 30981 35831
rect 33429 117763 33487 117817
rect 33551 117763 33609 117817
rect 33673 117763 33731 117817
rect 33795 117763 33853 117817
rect 32959 13057 33105 13189
rect 33293 13057 33439 13189
rect 33627 13057 33773 13189
rect 36757 80069 36811 80121
rect 36851 80069 36905 80121
rect 36945 80069 36999 80121
rect 36469 8339 36599 8445
rect 36727 8339 36857 8445
rect 36985 8339 37115 8445
rect 6387 4799 6441 4861
rect 6475 4799 6529 4861
rect 6561 4799 6615 4861
rect 6665 4799 6719 4861
rect 6769 4799 6823 4861
rect 6857 4799 6911 4861
<< metal3 >>
rect 2485 649507 2785 649511
rect 2485 642919 9209 649507
rect 2485 636195 167671 642919
rect 2485 634711 9209 636195
rect 3059 382079 44891 382157
rect 3059 381971 3427 382079
rect 3649 382071 44891 382079
rect 3649 382011 58864 382071
rect 3649 381971 44891 382011
rect 3059 381893 44891 381971
rect 3289 379301 3795 379357
rect 3289 379299 3481 379301
rect 1147 379187 3481 379299
rect 3289 379165 3481 379187
rect 3597 379299 3795 379301
rect 3597 379187 3925 379299
rect 3597 379165 3795 379187
rect 3289 379089 3795 379165
rect 43667 344377 44241 344409
rect 43667 344373 43703 344377
rect 43637 344313 43703 344373
rect 43667 344307 43703 344313
rect 43767 344307 43841 344377
rect 43905 344307 43979 344377
rect 44043 344307 44117 344377
rect 44181 344373 44241 344377
rect 44181 344313 70640 344373
rect 44181 344307 44241 344313
rect 43667 344277 44241 344307
rect 1883 336159 44308 336253
rect 1883 336079 43739 336159
rect 1267 336041 43739 336079
rect 43871 336041 43991 336159
rect 44123 336041 44308 336159
rect 1267 335969 44308 336041
rect 1267 335967 43739 335969
rect 1883 335851 43739 335967
rect 43871 335851 43991 335969
rect 44123 335851 44308 335969
rect 1883 335799 44308 335851
rect 43365 306697 43967 306735
rect 43365 306675 43393 306697
rect 43287 306615 43393 306675
rect 43365 306585 43393 306615
rect 43453 306585 43525 306697
rect 43585 306585 43657 306697
rect 43717 306585 43789 306697
rect 43849 306675 43967 306697
rect 43849 306615 53344 306675
rect 43849 306585 43967 306615
rect 43365 306539 43967 306585
rect 2061 292947 44090 293027
rect 2061 292855 43447 292947
rect 1293 292743 43447 292855
rect 2061 292707 43447 292743
rect 43619 292707 43725 292947
rect 43897 292707 44090 292947
rect 2061 292641 44090 292707
rect 42545 268903 43585 268955
rect 42545 268749 42645 268903
rect 42711 268749 42811 268903
rect 42877 268749 42977 268903
rect 43043 268749 43143 268903
rect 43209 268749 43309 268903
rect 43375 268855 43585 268903
rect 43375 268795 50032 268855
rect 43375 268749 43585 268795
rect 42545 268691 43585 268749
rect 1745 249833 43911 249985
rect 1269 249721 43911 249833
rect 1745 249601 43911 249721
rect 25876 231191 45241 231223
rect 25876 231043 26105 231191
rect 26199 231043 26271 231191
rect 26365 231043 26437 231191
rect 26531 231043 26603 231191
rect 26697 231157 45241 231191
rect 26697 231097 60428 231157
rect 26697 231043 45241 231097
rect 25876 231013 45241 231043
rect 27720 193395 44835 193461
rect 27720 193181 28009 193395
rect 28117 193181 28213 193395
rect 28321 193181 28417 193395
rect 28525 193181 28621 193395
rect 28729 193337 44835 193395
rect 28729 193277 45340 193337
rect 28729 193181 44835 193277
rect 27720 193131 44835 193181
rect 2409 178001 3357 178557
rect 2409 177583 2553 178001
rect 2981 177583 3357 178001
rect 2409 177187 3357 177583
rect 2409 176769 2553 177187
rect 2981 176769 3357 177187
rect 2409 176373 3357 176769
rect 2409 175955 2553 176373
rect 2981 175955 3357 176373
rect 2409 175559 3357 175955
rect 2409 175141 2553 175559
rect 2981 175141 3357 175559
rect 2409 174745 3357 175141
rect 2409 174327 2553 174745
rect 2981 174327 3357 174745
rect 2409 168033 3357 174327
rect 2409 167615 2647 168033
rect 3075 167615 3357 168033
rect 2409 167219 3357 167615
rect 2409 166801 2647 167219
rect 3075 166801 3357 167219
rect 2409 166405 3357 166801
rect 2409 165987 2647 166405
rect 3075 165987 3357 166405
rect 2409 165591 3357 165987
rect 2409 165173 2647 165591
rect 3075 165173 3357 165591
rect 2409 164777 3357 165173
rect 2409 164359 2647 164777
rect 3075 164359 3357 164777
rect 2409 163757 3357 164359
rect 30058 155645 44623 155683
rect 30058 155563 30311 155645
rect 30399 155563 30513 155645
rect 30601 155563 30715 155645
rect 30803 155563 30917 155645
rect 31005 155639 44623 155645
rect 31005 155579 45340 155639
rect 31005 155563 44623 155579
rect 30058 155537 44623 155563
rect 25589 122391 27015 122505
rect 25589 122295 25899 122391
rect 1941 122211 25899 122295
rect 1233 122099 25899 122211
rect 1941 122085 25899 122099
rect 26121 122085 26405 122391
rect 26627 122295 27015 122391
rect 26627 122085 27413 122295
rect 1941 122035 27413 122085
rect 25589 121911 27015 122035
rect 33407 117819 33865 117845
rect 33313 117817 61716 117819
rect 33313 117763 33429 117817
rect 33487 117763 33551 117817
rect 33609 117763 33673 117817
rect 33731 117763 33795 117817
rect 33853 117763 61716 117817
rect 33313 117759 61716 117763
rect 33407 117741 33865 117759
rect 36729 80121 37045 80161
rect 36655 80069 36757 80121
rect 36811 80069 36851 80121
rect 36905 80069 36945 80121
rect 36999 80069 51320 80121
rect 36655 80061 51320 80069
rect 36729 80031 37045 80061
rect 27849 79147 28963 79339
rect 27849 79107 28021 79147
rect 1667 78989 28021 79107
rect 1239 78877 28021 78989
rect 1667 78813 28021 78877
rect 27849 78783 28021 78813
rect 28185 78783 28307 79147
rect 28471 78783 28593 79147
rect 28757 78783 28963 79147
rect 27849 78661 28963 78783
rect 6201 42423 6859 42483
rect 6109 42407 47916 42423
rect 6109 42363 6279 42407
rect 6201 42341 6279 42363
rect 6363 42341 6459 42407
rect 6543 42341 6639 42407
rect 6723 42363 47916 42407
rect 6723 42341 6859 42363
rect 6201 42275 6859 42341
rect 2177 35831 31469 35973
rect 2177 35767 30329 35831
rect 1255 35655 30329 35767
rect 2177 35593 30329 35655
rect 30469 35593 30585 35831
rect 30725 35593 30841 35831
rect 30981 35593 31469 35831
rect 2177 35469 31469 35593
rect 32869 13189 33823 13281
rect 32869 13163 32959 13189
rect 1257 13057 32959 13163
rect 33105 13057 33293 13189
rect 33439 13057 33627 13189
rect 33773 13163 33823 13189
rect 33773 13057 34231 13163
rect 1257 13051 34231 13057
rect 32869 12973 33823 13051
rect 36385 8445 37403 8507
rect 36385 8435 36469 8445
rect 1281 8339 36469 8435
rect 36599 8339 36727 8445
rect 36857 8339 36985 8445
rect 37115 8435 37403 8445
rect 37115 8339 38287 8435
rect 1281 8323 38287 8339
rect 36385 8277 37403 8323
rect 6635 4889 6981 4905
rect 1201 4861 6981 4889
rect 1201 4799 6387 4861
rect 6441 4799 6475 4861
rect 6529 4799 6561 4861
rect 6615 4799 6665 4861
rect 6719 4799 6769 4861
rect 6823 4799 6857 4861
rect 6911 4799 6981 4861
rect 1201 4777 6981 4799
rect 6635 4753 6981 4777
<< via3 >>
rect 2553 177583 2981 178001
rect 2553 176769 2981 177187
rect 2553 175955 2981 176373
rect 2553 175141 2981 175559
rect 2553 174327 2981 174745
rect 2647 167615 3075 168033
rect 2647 166801 3075 167219
rect 2647 165987 3075 166405
rect 2647 165173 3075 165591
rect 2647 164359 3075 164777
<< metal4 >>
rect 36623 207867 42195 210925
rect 36623 207179 37079 207867
rect 37965 207179 38705 207867
rect 39591 207179 40331 207867
rect 41217 207179 42195 207867
rect 36623 206541 42195 207179
rect 36623 205853 37079 206541
rect 37965 205853 38705 206541
rect 39591 205853 40331 206541
rect 41217 205853 42195 206541
rect 36623 205215 42195 205853
rect 36623 204527 37079 205215
rect 37965 204527 38705 205215
rect 39591 204527 40331 205215
rect 41217 204527 42195 205215
rect 2381 178001 3331 178263
rect 2381 177583 2553 178001
rect 2981 177723 3331 178001
rect 2381 177313 2703 177583
rect 3107 177313 3331 177723
rect 2381 177187 3331 177313
rect 2381 176769 2553 177187
rect 2981 177003 3331 177187
rect 2381 176593 2703 176769
rect 3107 176593 3331 177003
rect 2381 176373 3331 176593
rect 2381 175955 2553 176373
rect 2981 176283 3331 176373
rect 2381 175873 2703 175955
rect 3107 175873 3331 176283
rect 2381 175563 3331 175873
rect 2381 175559 2703 175563
rect 2381 175141 2553 175559
rect 3107 175153 3331 175563
rect 2981 175141 3331 175153
rect 2381 174843 3331 175141
rect 2381 174745 2703 174843
rect 2381 174327 2553 174745
rect 3107 174433 3331 174843
rect 2981 174327 3331 174433
rect 2381 174085 3331 174327
rect 36623 177819 42195 204527
rect 36623 177079 37179 177819
rect 37997 177079 38581 177819
rect 39399 177079 39983 177819
rect 40801 177079 42195 177819
rect 36623 176515 42195 177079
rect 36623 175775 37179 176515
rect 37997 175775 38581 176515
rect 39399 175775 39983 176515
rect 40801 175775 42195 176515
rect 36623 175211 42195 175775
rect 36623 174471 37179 175211
rect 37997 174471 38581 175211
rect 39399 174471 39983 175211
rect 40801 174471 42195 175211
rect 36623 173805 42195 174471
rect 48921 207699 49541 382259
rect 48921 207359 49047 207699
rect 49395 207359 49541 207699
rect 48921 206951 49541 207359
rect 48921 206611 49047 206951
rect 49395 206611 49541 206951
rect 48921 206203 49541 206611
rect 48921 205863 49047 206203
rect 49395 205863 49541 206203
rect 48921 205455 49541 205863
rect 48921 205115 49047 205455
rect 49395 205115 49541 205455
rect 48921 204707 49541 205115
rect 48921 204367 49047 204707
rect 49395 204367 49541 204707
rect 48921 177697 49541 204367
rect 48921 177343 49043 177697
rect 49419 177343 49541 177697
rect 48921 176953 49541 177343
rect 48921 176599 49043 176953
rect 49419 176599 49541 176953
rect 48921 176209 49541 176599
rect 48921 175855 49043 176209
rect 49419 175855 49541 176209
rect 48921 175465 49541 175855
rect 48921 175111 49043 175465
rect 49419 175111 49541 175465
rect 48921 174721 49541 175111
rect 48921 174367 49043 174721
rect 49419 174367 49541 174721
rect 2521 168033 3471 168383
rect 2521 167615 2647 168033
rect 3075 167771 3471 168033
rect 2521 167361 2803 167615
rect 3207 167361 3471 167771
rect 2521 167219 3471 167361
rect 2521 166801 2647 167219
rect 3075 167051 3471 167219
rect 2521 166641 2803 166801
rect 3207 166641 3471 167051
rect 2521 166405 3471 166641
rect 2521 165987 2647 166405
rect 3075 166331 3471 166405
rect 2521 165921 2803 165987
rect 3207 165921 3471 166331
rect 2521 165611 3471 165921
rect 2521 165591 2803 165611
rect 2521 165173 2647 165591
rect 3207 165201 3471 165611
rect 3075 165173 3471 165201
rect 2521 164891 3471 165173
rect 2521 164777 2803 164891
rect 2521 164359 2647 164777
rect 3207 164481 3471 164891
rect 3075 164359 3471 164481
rect 2521 164205 3471 164359
rect 48921 167855 49541 174367
rect 48921 167501 49073 167855
rect 49449 167501 49541 167855
rect 48921 167111 49541 167501
rect 48921 166757 49073 167111
rect 49449 166757 49541 167111
rect 48921 166367 49541 166757
rect 48921 166013 49073 166367
rect 49449 166013 49541 166367
rect 48921 165623 49541 166013
rect 48921 165269 49073 165623
rect 49449 165269 49541 165623
rect 48921 164879 49541 165269
rect 48921 164525 49073 164879
rect 49449 164525 49541 164879
rect 48921 42259 49541 164525
rect 50161 42259 50781 382259
rect 57627 376979 64351 644945
rect 57627 376651 57997 376979
rect 58325 376651 58781 376979
rect 59109 376651 59565 376979
rect 59893 376651 60349 376979
rect 60677 376651 61133 376979
rect 61461 376651 61917 376979
rect 62245 376651 62701 376979
rect 63029 376651 63485 376979
rect 63813 376651 64351 376979
rect 57627 376549 64351 376651
rect 76909 376989 83633 644945
rect 76909 376661 77541 376989
rect 77869 376661 78325 376989
rect 78653 376661 79109 376989
rect 79437 376661 79893 376989
rect 80221 376661 80677 376989
rect 81005 376661 81461 376989
rect 81789 376661 82245 376989
rect 82573 376661 83029 376989
rect 83357 376661 83633 376989
rect 76909 376549 83633 376661
rect 96191 377039 102915 644945
rect 96191 376711 96721 377039
rect 97049 376711 97505 377039
rect 97833 376711 98289 377039
rect 98617 376711 99073 377039
rect 99401 376711 99857 377039
rect 100185 376711 100641 377039
rect 100969 376711 101425 377039
rect 101753 376711 102209 377039
rect 102537 376711 102915 377039
rect 96191 376549 102915 376711
rect 115473 377011 122197 644945
rect 115473 376683 115889 377011
rect 116217 376683 116757 377011
rect 117085 376683 117625 377011
rect 117953 376683 118493 377011
rect 118821 376683 119361 377011
rect 119689 376683 120229 377011
rect 120557 376683 121097 377011
rect 121425 376683 122197 377011
rect 115473 376549 122197 376683
rect 134755 377027 141479 644945
rect 134755 376699 135141 377027
rect 135469 376699 136071 377027
rect 136399 376699 137001 377027
rect 137329 376699 137931 377027
rect 138259 376699 138861 377027
rect 139189 376699 139791 377027
rect 140119 376699 140721 377027
rect 141049 376699 141479 377027
rect 134755 376549 141479 376699
rect 154037 377037 160761 644945
rect 154037 376709 154453 377037
rect 154781 376709 155279 377037
rect 155607 376709 156105 377037
rect 156433 376709 156931 377037
rect 157259 376709 157757 377037
rect 158085 376709 158583 377037
rect 158911 376709 159409 377037
rect 159737 376709 160761 377037
rect 154037 376549 160761 376709
<< via4 >>
rect 37079 207179 37965 207867
rect 38705 207179 39591 207867
rect 40331 207179 41217 207867
rect 37079 205853 37965 206541
rect 38705 205853 39591 206541
rect 40331 205853 41217 206541
rect 37079 204527 37965 205215
rect 38705 204527 39591 205215
rect 40331 204527 41217 205215
rect 2703 177583 2981 177723
rect 2981 177583 3107 177723
rect 2703 177313 3107 177583
rect 2703 176769 2981 177003
rect 2981 176769 3107 177003
rect 2703 176593 3107 176769
rect 2703 175955 2981 176283
rect 2981 175955 3107 176283
rect 2703 175873 3107 175955
rect 2703 175559 3107 175563
rect 2703 175153 2981 175559
rect 2981 175153 3107 175559
rect 2703 174745 3107 174843
rect 2703 174433 2981 174745
rect 2981 174433 3107 174745
rect 37179 177079 37997 177819
rect 38581 177079 39399 177819
rect 39983 177079 40801 177819
rect 37179 175775 37997 176515
rect 38581 175775 39399 176515
rect 39983 175775 40801 176515
rect 37179 174471 37997 175211
rect 38581 174471 39399 175211
rect 39983 174471 40801 175211
rect 49047 207359 49395 207699
rect 49047 206611 49395 206951
rect 49047 205863 49395 206203
rect 49047 205115 49395 205455
rect 49047 204367 49395 204707
rect 49043 177343 49419 177697
rect 49043 176599 49419 176953
rect 49043 175855 49419 176209
rect 49043 175111 49419 175465
rect 49043 174367 49419 174721
rect 2803 167615 3075 167771
rect 3075 167615 3207 167771
rect 2803 167361 3207 167615
rect 2803 166801 3075 167051
rect 3075 166801 3207 167051
rect 2803 166641 3207 166801
rect 2803 165987 3075 166331
rect 3075 165987 3207 166331
rect 2803 165921 3207 165987
rect 2803 165591 3207 165611
rect 2803 165201 3075 165591
rect 3075 165201 3207 165591
rect 2803 164777 3207 164891
rect 2803 164481 3075 164777
rect 3075 164481 3207 164777
rect 49073 167501 49449 167855
rect 49073 166757 49449 167111
rect 49073 166013 49449 166367
rect 49073 165269 49449 165623
rect 49073 164525 49449 164879
rect 57997 376651 58325 376979
rect 58781 376651 59109 376979
rect 59565 376651 59893 376979
rect 60349 376651 60677 376979
rect 61133 376651 61461 376979
rect 61917 376651 62245 376979
rect 62701 376651 63029 376979
rect 63485 376651 63813 376979
rect 77541 376661 77869 376989
rect 78325 376661 78653 376989
rect 79109 376661 79437 376989
rect 79893 376661 80221 376989
rect 80677 376661 81005 376989
rect 81461 376661 81789 376989
rect 82245 376661 82573 376989
rect 83029 376661 83357 376989
rect 96721 376711 97049 377039
rect 97505 376711 97833 377039
rect 98289 376711 98617 377039
rect 99073 376711 99401 377039
rect 99857 376711 100185 377039
rect 100641 376711 100969 377039
rect 101425 376711 101753 377039
rect 102209 376711 102537 377039
rect 115889 376683 116217 377011
rect 116757 376683 117085 377011
rect 117625 376683 117953 377011
rect 118493 376683 118821 377011
rect 119361 376683 119689 377011
rect 120229 376683 120557 377011
rect 135141 376699 135469 377027
rect 136071 376699 136399 377027
rect 137001 376699 137329 377027
rect 137931 376699 138259 377027
rect 138861 376699 139189 377027
rect 139791 376699 140119 377027
rect 140721 376699 141049 377027
rect 154453 376709 154781 377037
rect 155279 376709 155607 377037
rect 156105 376709 156433 377037
rect 156931 376709 157259 377037
rect 157757 376709 158085 377037
rect 158583 376709 158911 377037
rect 159409 376709 159737 377037
<< metal5 >>
rect 45077 377787 165045 378407
rect 45077 377039 165045 377167
rect 45077 376989 96721 377039
rect 45077 376979 77541 376989
rect 45077 376651 57997 376979
rect 58325 376651 58781 376979
rect 59109 376651 59565 376979
rect 59893 376651 60349 376979
rect 60677 376651 61133 376979
rect 61461 376651 61917 376979
rect 62245 376651 62701 376979
rect 63029 376651 63485 376979
rect 63813 376661 77541 376979
rect 77869 376661 78325 376989
rect 78653 376661 79109 376989
rect 79437 376661 79893 376989
rect 80221 376661 80677 376989
rect 81005 376661 81461 376989
rect 81789 376661 82245 376989
rect 82573 376661 83029 376989
rect 83357 376711 96721 376989
rect 97049 376711 97505 377039
rect 97833 376711 98289 377039
rect 98617 376711 99073 377039
rect 99401 376711 99857 377039
rect 100185 376711 100641 377039
rect 100969 376711 101425 377039
rect 101753 376711 102209 377039
rect 102537 377037 165045 377039
rect 102537 377027 154453 377037
rect 102537 377011 135141 377027
rect 102537 376711 115889 377011
rect 83357 376683 115889 376711
rect 116217 376683 116757 377011
rect 117085 376683 117625 377011
rect 117953 376683 118493 377011
rect 118821 376683 119361 377011
rect 119689 376683 120229 377011
rect 120557 376699 135141 377011
rect 135469 376699 136071 377027
rect 136399 376699 137001 377027
rect 137329 376699 137931 377027
rect 138259 376699 138861 377027
rect 139189 376699 139791 377027
rect 140119 376699 140721 377027
rect 141049 376709 154453 377027
rect 154781 376709 155279 377037
rect 155607 376709 156105 377037
rect 156433 376709 156931 377037
rect 157259 376709 157757 377037
rect 158085 376709 158583 377037
rect 158911 376709 159409 377037
rect 159737 376709 165045 377037
rect 141049 376699 165045 376709
rect 120557 376683 165045 376699
rect 83357 376661 165045 376683
rect 63813 376651 165045 376661
rect 45077 376547 165045 376651
rect 36525 207867 49559 208537
rect 36525 207179 37079 207867
rect 37965 207179 38705 207867
rect 39591 207179 40331 207867
rect 41217 207699 49559 207867
rect 41217 207359 49047 207699
rect 49395 207359 49559 207699
rect 41217 207179 49559 207359
rect 36525 206951 49559 207179
rect 36525 206611 49047 206951
rect 49395 206611 49559 206951
rect 36525 206541 49559 206611
rect 36525 205853 37079 206541
rect 37965 205853 38705 206541
rect 39591 205853 40331 206541
rect 41217 206203 49559 206541
rect 41217 205863 49047 206203
rect 49395 205863 49559 206203
rect 41217 205853 49559 205863
rect 36525 205455 49559 205853
rect 36525 205215 49047 205455
rect 36525 204527 37079 205215
rect 37965 204527 38705 205215
rect 39591 204527 40331 205215
rect 41217 205115 49047 205215
rect 49395 205115 49559 205455
rect 41217 204707 49559 205115
rect 41217 204527 49047 204707
rect 36525 204367 49047 204527
rect 49395 204367 49559 204707
rect 36525 204165 49559 204367
rect 2523 177819 49694 178147
rect 2523 177723 37179 177819
rect 2523 177313 2703 177723
rect 3107 177313 37179 177723
rect 2523 177079 37179 177313
rect 37997 177079 38581 177819
rect 39399 177079 39983 177819
rect 40801 177697 49694 177819
rect 40801 177343 49043 177697
rect 49419 177343 49694 177697
rect 40801 177079 49694 177343
rect 2523 177003 49694 177079
rect 2523 176593 2703 177003
rect 3107 176953 49694 177003
rect 3107 176599 49043 176953
rect 49419 176599 49694 176953
rect 3107 176593 49694 176599
rect 2523 176515 49694 176593
rect 2523 176283 37179 176515
rect 2523 175873 2703 176283
rect 3107 175873 37179 176283
rect 2523 175775 37179 175873
rect 37997 175775 38581 176515
rect 39399 175775 39983 176515
rect 40801 176209 49694 176515
rect 40801 175855 49043 176209
rect 49419 175855 49694 176209
rect 40801 175775 49694 175855
rect 2523 175563 49694 175775
rect 2523 175153 2703 175563
rect 3107 175465 49694 175563
rect 3107 175211 49043 175465
rect 3107 175153 37179 175211
rect 2523 174843 37179 175153
rect 2523 174433 2703 174843
rect 3107 174471 37179 174843
rect 37997 174471 38581 175211
rect 39399 174471 39983 175211
rect 40801 175111 49043 175211
rect 49419 175111 49694 175465
rect 40801 174721 49694 175111
rect 40801 174471 49043 174721
rect 3107 174433 49043 174471
rect 2523 174367 49043 174433
rect 49419 174367 49694 174721
rect 2523 174217 49694 174367
rect 2613 167855 49836 168229
rect 2613 167771 49073 167855
rect 2613 167361 2803 167771
rect 3207 167501 49073 167771
rect 49449 167501 49836 167855
rect 3207 167361 49836 167501
rect 2613 167111 49836 167361
rect 2613 167051 49073 167111
rect 2613 166641 2803 167051
rect 3207 166757 49073 167051
rect 49449 166757 49836 167111
rect 3207 166641 49836 166757
rect 2613 166367 49836 166641
rect 2613 166331 49073 166367
rect 2613 165921 2803 166331
rect 3207 166013 49073 166331
rect 49449 166013 49836 166367
rect 3207 165921 49836 166013
rect 2613 165623 49836 165921
rect 2613 165611 49073 165623
rect 2613 165201 2803 165611
rect 3207 165269 49073 165611
rect 49449 165269 49836 165623
rect 3207 165201 49836 165269
rect 2613 164891 49836 165201
rect 2613 164481 2803 164891
rect 3207 164879 49836 164891
rect 3207 164525 49073 164879
rect 49449 164525 49836 164879
rect 3207 164481 49836 164525
rect 2613 164299 49836 164481
use puf_super  puf_super_0
timestamp 1654736712
transform 1 0 45077 0 1 42259
box 0 0 119968 340000
<< end >>
