magic
tech sky130A
magscale 1 2
timestamp 1656729169
<< metal3 >>
rect -1139 152 1138 180
rect -1139 -152 -1112 152
rect 1112 -152 1138 152
rect -1139 -180 1138 -152
<< via3 >>
rect -1112 -152 1112 152
<< metal4 >>
rect -1139 152 1138 180
rect -1139 -152 -1112 152
rect 1112 -152 1138 152
rect -1139 -180 1138 -152
<< properties >>
string GDS_END 9347970
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/merge/design_merged.gds
string GDS_START 9340670
<< end >>
