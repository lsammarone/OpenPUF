magic
tech sky130A
magscale 1 2
timestamp 1656715967
<< error_p >>
rect -23 17 23 29
rect -23 -17 17 17
rect -23 -29 23 -17
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -23 17 23 29
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -29 23 -17
<< properties >>
string GDS_END 9298302
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/design_merged.gds
string GDS_START 9298106
<< end >>
