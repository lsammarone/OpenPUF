magic
tech sky130A
magscale 1 2
timestamp 1656729169
<< nwell >>
rect -406 636 388 882
rect -574 -766 -356 -198
rect -62 -278 382 -258
rect -62 -444 416 -278
rect 690 -416 1048 -200
rect -62 -452 434 -444
rect 202 -594 434 -452
<< locali >>
rect 92 452 142 456
rect 460 452 526 484
rect 92 443 526 452
rect 92 409 100 443
rect 134 436 526 443
rect 134 409 580 436
rect 92 402 580 409
rect 92 400 142 402
rect -342 319 -304 322
rect -342 285 -340 319
rect -306 285 -304 319
rect -342 282 -304 285
rect -164 317 -124 318
rect -164 283 -161 317
rect -127 283 -124 317
rect -164 282 -124 283
rect -252 219 -208 224
rect -252 185 -247 219
rect -213 185 -208 219
rect -252 180 -208 185
rect -248 -63 -204 -58
rect -248 -97 -243 -63
rect -209 -97 -204 -63
rect -248 -102 -204 -97
rect -342 -161 -304 -158
rect -342 -195 -340 -161
rect -306 -195 -304 -161
rect -342 -198 -304 -195
rect -164 -161 -126 -158
rect -164 -195 -162 -161
rect -128 -195 -126 -161
rect -164 -198 -126 -195
rect 1044 -165 1082 -162
rect 1044 -199 1046 -165
rect 1080 -199 1082 -165
rect 1044 -202 1082 -199
rect 1218 -357 1256 -354
rect 1218 -391 1220 -357
rect 1254 -391 1256 -357
rect 1218 -394 1256 -391
rect 276 -599 334 -590
rect 276 -633 284 -599
rect 318 -602 334 -599
rect 464 -602 530 -522
rect 318 -633 588 -602
rect 276 -636 588 -633
rect 276 -642 334 -636
rect -384 -769 -288 -764
rect -384 -803 -372 -769
rect -338 -803 -288 -769
rect -384 -810 -288 -803
rect -176 -771 10 -764
rect -176 -805 -62 -771
rect -28 -805 10 -771
rect -176 -810 10 -805
rect 1040 -781 1078 -778
rect 1040 -815 1042 -781
rect 1076 -815 1078 -781
rect 1040 -818 1078 -815
rect 80 -849 118 -846
rect 80 -883 82 -849
rect 116 -883 118 -849
rect 80 -886 118 -883
<< viali >>
rect 100 409 134 443
rect -340 285 -306 319
rect -161 283 -127 317
rect -247 185 -213 219
rect -243 -97 -209 -63
rect -340 -195 -306 -161
rect -162 -195 -128 -161
rect 1046 -199 1080 -165
rect 1220 -391 1254 -357
rect 284 -633 318 -599
rect -372 -803 -338 -769
rect -62 -805 -28 -771
rect 1042 -815 1076 -781
rect 82 -883 116 -849
<< metal1 >>
rect -574 1120 1322 1192
rect -574 1004 961 1120
rect 1269 1004 1322 1120
rect -574 938 1322 1004
rect -366 634 -300 938
rect 92 456 146 458
rect -16 454 146 456
rect -16 402 -6 454
rect 46 443 146 454
rect 46 409 100 443
rect 134 409 146 443
rect 46 402 146 409
rect -16 400 146 402
rect 92 394 146 400
rect -428 328 -296 338
rect -428 276 -422 328
rect -370 319 -296 328
rect -370 285 -340 319
rect -306 285 -296 319
rect -370 276 -296 285
rect -178 336 -102 344
rect -178 284 -168 336
rect -116 332 -102 336
rect 258 342 406 350
rect -116 284 -60 332
rect -178 283 -161 284
rect -127 283 -60 284
rect -178 276 -60 283
rect 258 290 270 342
rect 322 290 406 342
rect 258 280 406 290
rect -428 266 -296 276
rect -266 230 94 234
rect -266 219 20 230
rect -266 185 -247 219
rect -213 185 20 219
rect -266 178 20 185
rect 72 178 94 230
rect -266 168 94 178
rect -118 34 432 110
rect -262 -52 98 -48
rect -262 -63 24 -52
rect -262 -97 -243 -63
rect -209 -97 24 -63
rect -262 -104 24 -97
rect 76 -104 98 -52
rect 850 -64 920 938
rect -262 -114 98 -104
rect 206 -140 920 -64
rect -428 -152 -296 -142
rect -428 -204 -422 -152
rect -370 -161 -296 -152
rect -370 -195 -340 -161
rect -306 -195 -296 -161
rect -370 -204 -296 -195
rect -428 -214 -296 -204
rect -178 -161 -96 -152
rect -178 -166 -162 -161
rect -128 -166 -96 -161
rect -178 -218 -166 -166
rect -114 -218 -96 -166
rect -178 -230 -96 -218
rect 206 -176 282 -140
rect 258 -228 282 -176
rect 800 -228 810 -176
rect 206 -434 282 -228
rect 792 -236 810 -228
rect 628 -285 686 -282
rect 392 -294 462 -286
rect 392 -346 401 -294
rect 453 -346 462 -294
rect 628 -337 631 -285
rect 683 -337 686 -285
rect 628 -340 686 -337
rect 392 -354 462 -346
rect 186 -458 282 -434
rect 186 -510 208 -458
rect 260 -510 282 -458
rect 186 -530 282 -510
rect 844 -454 920 -140
rect 986 -150 1096 -134
rect 986 -202 998 -150
rect 1050 -165 1096 -150
rect 1080 -199 1096 -165
rect 1050 -202 1096 -199
rect 986 -210 1096 -202
rect 1202 -357 1298 -326
rect 1202 -391 1220 -357
rect 1254 -391 1298 -357
rect 1202 -404 1298 -391
rect 844 -530 1052 -454
rect 268 -599 334 -590
rect 268 -600 284 -599
rect -50 -632 284 -600
rect -50 -730 -18 -632
rect 268 -633 284 -632
rect 318 -633 334 -599
rect 268 -642 334 -633
rect -534 -766 -320 -754
rect -56 -760 -12 -730
rect -534 -818 -526 -766
rect -474 -769 -320 -766
rect -474 -803 -372 -769
rect -338 -803 -320 -769
rect -474 -818 -320 -803
rect -80 -762 -12 -760
rect -80 -814 -70 -762
rect -18 -814 -12 -762
rect 972 -772 1096 -756
rect -534 -826 -320 -818
rect 972 -824 982 -772
rect 1034 -781 1096 -772
rect 1034 -815 1042 -781
rect 1076 -815 1096 -781
rect 1034 -824 1096 -815
rect 972 -830 1096 -824
rect 68 -849 134 -834
rect 68 -883 82 -849
rect 116 -850 134 -849
rect 116 -883 500 -850
rect 68 -894 500 -883
rect -566 -970 1224 -930
rect -566 -1022 -264 -970
rect -212 -1022 -186 -970
rect -134 -1004 1224 -970
rect 1284 -1004 1322 -930
rect -134 -1022 961 -1004
rect -566 -1120 961 -1022
rect 1269 -1120 1322 -1004
rect -566 -1184 1322 -1120
<< via1 >>
rect 961 1004 1269 1120
rect -6 402 46 454
rect -422 276 -370 328
rect -168 317 -116 336
rect -168 284 -161 317
rect -161 284 -127 317
rect -127 284 -116 317
rect 270 290 322 342
rect 642 252 694 304
rect 20 178 72 230
rect 746 156 798 208
rect -266 38 -214 90
rect 24 -104 76 -52
rect 1112 28 1164 80
rect -422 -204 -370 -152
rect -166 -195 -162 -166
rect -162 -195 -128 -166
rect -128 -195 -114 -166
rect -166 -218 -114 -195
rect 206 -228 258 -176
rect 748 -228 800 -176
rect 401 -346 453 -294
rect 631 -337 683 -285
rect 208 -510 260 -458
rect 998 -165 1050 -150
rect 998 -199 1046 -165
rect 1046 -199 1050 -165
rect 998 -202 1050 -199
rect -526 -818 -474 -766
rect -70 -771 -18 -762
rect -70 -805 -62 -771
rect -62 -805 -28 -771
rect -28 -805 -18 -771
rect -70 -814 -18 -805
rect 982 -824 1034 -772
rect -264 -1022 -212 -970
rect -186 -1022 -134 -970
rect 961 -1120 1269 -1004
<< metal2 >>
rect 940 1120 1290 1134
rect 940 1004 961 1120
rect 1269 1004 1290 1120
rect 940 990 1290 1004
rect -566 816 1050 844
rect -436 332 -364 346
rect -124 344 -96 816
rect 528 512 600 520
rect -574 328 -364 332
rect -574 276 -422 328
rect -370 276 -364 328
rect -178 336 -96 344
rect -178 284 -168 336
rect -116 284 -96 336
rect -178 276 -96 284
rect -574 270 -364 276
rect -436 260 -364 270
rect -266 90 -214 110
rect -436 -144 -396 -134
rect -436 -148 -364 -144
rect -574 -152 -364 -148
rect -574 -204 -422 -152
rect -370 -204 -364 -152
rect -574 -210 -364 -204
rect -436 -220 -364 -210
rect -554 -754 -510 -398
rect -554 -766 -462 -754
rect -554 -818 -526 -766
rect -474 -818 -462 -766
rect -554 -826 -462 -818
rect -554 -1014 -510 -826
rect -266 -962 -214 38
rect -124 -152 -96 276
rect -178 -166 -96 -152
rect -178 -218 -166 -166
rect -114 -218 -96 -166
rect -178 -230 -96 -218
rect -36 454 46 464
rect -36 402 -6 454
rect 528 456 532 512
rect 588 456 600 512
rect 528 450 600 456
rect 1002 512 1082 528
rect 1002 456 1014 512
rect 1070 456 1082 512
rect 1002 450 1082 456
rect 1196 512 1272 522
rect 1196 456 1208 512
rect 1264 456 1272 512
rect -36 396 46 402
rect -36 -748 -8 396
rect 258 342 344 350
rect 258 290 270 342
rect 322 290 344 342
rect 20 231 122 236
rect 20 230 35 231
rect 20 175 35 178
rect 91 175 122 231
rect 20 170 122 175
rect 24 -51 126 -46
rect 24 -52 39 -51
rect 24 -107 39 -104
rect 95 -107 126 -51
rect 316 -52 344 290
rect 622 304 710 306
rect 622 252 642 304
rect 694 252 710 304
rect 622 238 710 252
rect 384 232 470 236
rect 384 176 396 232
rect 452 176 470 232
rect 24 -112 126 -107
rect 258 -108 272 -52
rect 328 -108 344 -52
rect 258 -112 344 -108
rect 206 -176 258 -166
rect 206 -448 258 -228
rect 442 -286 470 176
rect 622 182 640 238
rect 696 182 710 238
rect 622 172 710 182
rect 742 208 808 214
rect 742 156 746 208
rect 798 156 808 208
rect 742 144 808 156
rect 384 -294 470 -286
rect 384 -346 401 -294
rect 453 -346 470 -294
rect 622 -48 696 -33
rect 622 -104 631 -48
rect 687 -104 696 -48
rect 622 -285 696 -104
rect 742 -170 796 144
rect 1022 -134 1050 450
rect 1196 448 1272 456
rect 1244 332 1272 448
rect 1244 270 1322 332
rect 1112 80 1164 116
rect 986 -150 1058 -134
rect 742 -176 808 -170
rect 742 -228 748 -176
rect 800 -228 808 -176
rect 986 -202 998 -150
rect 1050 -202 1058 -150
rect 986 -210 1058 -202
rect 742 -236 808 -228
rect 622 -337 631 -285
rect 683 -337 696 -285
rect 622 -344 696 -337
rect 384 -360 470 -346
rect 578 -440 614 -420
rect 188 -458 282 -448
rect 188 -510 208 -458
rect 260 -510 282 -458
rect 536 -496 538 -440
rect 594 -496 614 -440
rect 578 -506 614 -496
rect 996 -440 1076 -424
rect 996 -496 1008 -440
rect 1064 -496 1076 -440
rect 996 -502 1076 -496
rect 188 -530 282 -510
rect -80 -762 -8 -748
rect 1016 -754 1044 -502
rect -80 -814 -70 -762
rect -18 -814 -8 -762
rect 970 -772 1046 -754
rect 970 -824 982 -772
rect 1034 -824 1046 -772
rect 970 -832 1046 -824
rect -276 -970 -124 -962
rect -276 -1022 -264 -970
rect -212 -1022 -186 -970
rect -134 -1022 -124 -970
rect 1112 -990 1164 28
rect 1218 -210 1322 -148
rect 1218 -430 1246 -210
rect 1206 -440 1276 -430
rect 1206 -496 1208 -440
rect 1264 -496 1276 -440
rect 1206 -506 1276 -496
rect -276 -1028 -124 -1022
rect 940 -1004 1290 -990
rect 940 -1120 961 -1004
rect 1269 -1120 1290 -1004
rect 940 -1134 1290 -1120
<< via2 >>
rect 967 1034 1023 1090
rect 1047 1034 1103 1090
rect 1127 1034 1183 1090
rect 1207 1034 1263 1090
rect 532 456 588 512
rect 1014 456 1070 512
rect 1208 456 1264 512
rect 35 230 91 231
rect 35 178 72 230
rect 72 178 91 230
rect 35 175 91 178
rect 39 -52 95 -51
rect 39 -104 76 -52
rect 76 -104 95 -52
rect 39 -107 95 -104
rect 396 176 452 232
rect 272 -108 328 -52
rect 640 182 696 238
rect 631 -104 687 -48
rect 538 -496 594 -440
rect 1008 -496 1064 -440
rect 1208 -496 1264 -440
rect 967 -1090 1023 -1034
rect 1047 -1090 1103 -1034
rect 1127 -1090 1183 -1034
rect 1207 -1090 1263 -1034
<< metal3 >>
rect -574 1090 1322 1192
rect -574 1034 967 1090
rect 1023 1034 1047 1090
rect 1103 1034 1127 1090
rect 1183 1034 1207 1090
rect 1263 1034 1322 1090
rect -574 938 1322 1034
rect 514 512 1278 520
rect 514 456 532 512
rect 588 456 1014 512
rect 1070 456 1208 512
rect 1264 456 1278 512
rect 514 450 1278 456
rect 10 237 162 250
rect 626 238 706 244
rect 626 237 640 238
rect 10 232 640 237
rect 10 231 396 232
rect 10 175 35 231
rect 91 176 396 231
rect 452 182 640 232
rect 696 237 706 238
rect 696 182 717 237
rect 452 176 717 182
rect 91 175 717 176
rect 10 171 717 175
rect 10 158 162 171
rect 14 -45 166 -32
rect 622 -45 696 -32
rect 14 -48 721 -45
rect 14 -51 631 -48
rect 14 -107 39 -51
rect 95 -52 631 -51
rect 95 -107 272 -52
rect 14 -108 272 -107
rect 328 -104 631 -52
rect 687 -104 721 -48
rect 328 -108 721 -104
rect 14 -111 721 -108
rect 14 -124 166 -111
rect 258 -118 344 -111
rect 526 -440 1276 -420
rect 526 -496 538 -440
rect 594 -496 1008 -440
rect 1064 -496 1208 -440
rect 1264 -496 1276 -440
rect 526 -506 1276 -496
rect -566 -1034 1322 -930
rect -566 -1090 967 -1034
rect 1023 -1090 1047 -1034
rect 1103 -1090 1127 -1034
rect 1183 -1090 1207 -1034
rect 1263 -1090 1322 -1034
rect -566 -1185 1322 -1090
use mux  mux_0
timestamp 1656729169
transform 1 0 432 0 1 146
box -54 -122 366 878
use mux  mux_1
timestamp 1656729169
transform 1 0 436 0 1 -892
box -54 -122 366 878
use mux  mux_2
timestamp 1656729169
transform 1 0 432 0 1 146
box -54 -122 366 878
use mux  mux_3
timestamp 1656729169
transform 1 0 436 0 1 -892
box -54 -122 366 878
use mux  mux_4
timestamp 1656729169
transform 1 0 432 0 1 146
box -54 -122 366 878
use mux  mux_5
timestamp 1656729169
transform 1 0 436 0 1 -892
box -54 -122 366 878
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_0
timestamp 1656729169
transform 1 0 1008 0 1 -1027
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_1
timestamp 1656729169
transform 1 0 1008 0 -1 61
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_2
timestamp 1656729169
transform 1 0 1008 0 1 -1027
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_3
timestamp 1656729169
transform 1 0 1008 0 -1 61
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_4
timestamp 1656729169
transform 1 0 1008 0 1 -1027
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_5
timestamp 1656729169
transform 1 0 1008 0 -1 61
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1#0  sky130_fd_sc_hd__inv_1#0_0
timestamp 1656729169
transform 1 0 -90 0 1 -1026
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1#0  sky130_fd_sc_hd__inv_1#0_1
timestamp 1656729169
transform 1 0 -366 0 1 -1026
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1#0  sky130_fd_sc_hd__inv_1#0_2
timestamp 1656729169
transform 1 0 -90 0 1 -1026
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1#0  sky130_fd_sc_hd__inv_1#0_3
timestamp 1656729169
transform 1 0 -366 0 1 -1026
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1#0  sky130_fd_sc_hd__inv_1_0
timestamp 1656729169
transform 1 0 -90 0 1 -1026
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1#0  sky130_fd_sc_hd__inv_1_1
timestamp 1656729169
transform 1 0 -366 0 1 -1026
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_0
timestamp 1656729169
transform 1 0 -366 0 1 62
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_1
timestamp 1656729169
transform 1 0 -366 0 -1 62
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_2
timestamp 1656729169
transform 1 0 -366 0 1 62
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_3
timestamp 1656729169
transform 1 0 -366 0 -1 62
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_4
timestamp 1656729169
transform 1 0 -366 0 1 62
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_5
timestamp 1656729169
transform 1 0 -366 0 -1 62
box -38 -48 314 592
<< properties >>
string GDS_END 10039168
string GDS_FILE /scratch/users/lsammaro/OpenPUF/mag/merge/design_merged.gds
string GDS_START 9995172
<< end >>
