magic
tech sky130A
timestamp 1483428465
<< checkpaint >>
rect -716 -654 716 654
<< metal3 >>
rect -86 16 86 24
rect -86 -16 -76 16
rect -44 -16 -36 16
rect -4 -16 4 16
rect 36 -16 44 16
rect 76 -16 86 16
rect -86 -24 86 -16
<< via3 >>
rect -76 -16 -44 16
rect -36 -16 -4 16
rect 4 -16 36 16
rect 44 -16 76 16
<< metal4 >>
rect -86 16 86 24
rect -86 -16 -76 16
rect -44 -16 -36 16
rect -4 -16 4 16
rect 36 -16 44 16
rect 76 -16 86 16
rect -86 -24 86 -16
<< end >>
