magic
tech sky130A
timestamp 1483428465
<< checkpaint >>
rect -1130 -1130 1130 1130
<< metal4 >>
rect -500 459 500 500
rect -500 -459 -459 459
rect 459 -459 500 459
rect -500 -500 500 -459
<< via4 >>
rect -459 -459 459 459
<< metal5 >>
rect -500 459 500 500
rect -500 -459 -459 459
rect 459 -459 500 459
rect -500 -500 500 -459
<< end >>
