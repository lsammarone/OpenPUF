magic
tech sky130A
timestamp 1483428465
<< checkpaint >>
rect -1130 -994 1130 994
<< metal4 >>
rect -500 299 500 364
rect -500 -299 -459 299
rect 459 -299 500 299
rect -500 -364 500 -299
<< via4 >>
rect -459 -299 459 299
<< metal5 >>
rect -500 299 500 364
rect -500 -299 -459 299
rect 459 -299 500 299
rect -500 -364 500 -299
<< end >>
