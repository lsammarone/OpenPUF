magic
tech sky130A
magscale 1 2
timestamp 1483428465
<< checkpaint >>
rect -1652 -2223 1652 2223
<< metal4 >>
rect -392 918 392 963
rect -392 -918 -278 918
rect 278 -918 392 918
rect -392 -963 392 -918
<< via4 >>
rect -278 -918 278 918
<< metal5 >>
rect -392 918 392 963
rect -392 -918 -278 918
rect 278 -918 392 918
rect -392 -963 392 -918
<< end >>
