magic
tech sky130A
timestamp 1483428465
<< checkpaint >>
rect -902 -720 902 720
<< metal3 >>
rect -272 76 272 90
rect -272 -76 -256 76
rect 256 -76 272 76
rect -272 -90 272 -76
<< via3 >>
rect -256 -76 256 76
<< metal4 >>
rect -272 76 272 90
rect -272 -76 -256 76
rect 256 -76 272 76
rect -272 -90 272 -76
<< end >>
